// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Dec 6 2024 13:45:26

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    CMA,
    DRA,
    A,
    TSn,
    CLMBEn,
    AWEn,
    RESETn,
    CASn,
    BANK0,
    VBENn,
    CUMBEn,
    CLKRAM,
    C3,
    ASn,
    LDSn,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CASLn,
    RAMSPACEn,
    WEn,
    REGENn,
    DBRn,
    CLK40C,
    CLK40_IN,
    REGSPACEn,
    RAMENn,
    RASn,
    TACKn,
    CLKEN,
    C1);

    input [1:0] SIZ;
    output [10:0] CMA;
    input [9:0] DRA;
    input [20:0] A;
    input TSn;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CASn;
    output BANK0;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    input C3;
    output ASn;
    output LDSn;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    input CASLn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    input DBRn;
    output CLK40C;
    input CLK40_IN;
    input REGSPACEn;
    output RAMENn;
    output RASn;
    output TACKn;
    output CLKEN;
    input C1;

    wire N__10065;
    wire N__10064;
    wire N__10063;
    wire N__10056;
    wire N__10055;
    wire N__10054;
    wire N__10047;
    wire N__10046;
    wire N__10045;
    wire N__10038;
    wire N__10037;
    wire N__10036;
    wire N__10029;
    wire N__10028;
    wire N__10027;
    wire N__10020;
    wire N__10019;
    wire N__10018;
    wire N__10011;
    wire N__10010;
    wire N__10009;
    wire N__10002;
    wire N__10001;
    wire N__10000;
    wire N__9993;
    wire N__9992;
    wire N__9991;
    wire N__9984;
    wire N__9983;
    wire N__9982;
    wire N__9975;
    wire N__9974;
    wire N__9973;
    wire N__9966;
    wire N__9965;
    wire N__9964;
    wire N__9957;
    wire N__9956;
    wire N__9955;
    wire N__9948;
    wire N__9947;
    wire N__9946;
    wire N__9939;
    wire N__9938;
    wire N__9937;
    wire N__9930;
    wire N__9929;
    wire N__9928;
    wire N__9921;
    wire N__9920;
    wire N__9919;
    wire N__9912;
    wire N__9911;
    wire N__9910;
    wire N__9903;
    wire N__9902;
    wire N__9901;
    wire N__9894;
    wire N__9893;
    wire N__9892;
    wire N__9885;
    wire N__9884;
    wire N__9883;
    wire N__9876;
    wire N__9875;
    wire N__9874;
    wire N__9867;
    wire N__9866;
    wire N__9865;
    wire N__9858;
    wire N__9857;
    wire N__9856;
    wire N__9849;
    wire N__9848;
    wire N__9847;
    wire N__9840;
    wire N__9839;
    wire N__9838;
    wire N__9831;
    wire N__9830;
    wire N__9829;
    wire N__9822;
    wire N__9821;
    wire N__9820;
    wire N__9813;
    wire N__9812;
    wire N__9811;
    wire N__9804;
    wire N__9803;
    wire N__9802;
    wire N__9795;
    wire N__9794;
    wire N__9793;
    wire N__9786;
    wire N__9785;
    wire N__9784;
    wire N__9777;
    wire N__9776;
    wire N__9775;
    wire N__9768;
    wire N__9767;
    wire N__9766;
    wire N__9759;
    wire N__9758;
    wire N__9757;
    wire N__9750;
    wire N__9749;
    wire N__9748;
    wire N__9741;
    wire N__9740;
    wire N__9739;
    wire N__9732;
    wire N__9731;
    wire N__9730;
    wire N__9723;
    wire N__9722;
    wire N__9721;
    wire N__9714;
    wire N__9713;
    wire N__9712;
    wire N__9705;
    wire N__9704;
    wire N__9703;
    wire N__9696;
    wire N__9695;
    wire N__9694;
    wire N__9687;
    wire N__9686;
    wire N__9685;
    wire N__9678;
    wire N__9677;
    wire N__9676;
    wire N__9669;
    wire N__9668;
    wire N__9667;
    wire N__9660;
    wire N__9659;
    wire N__9658;
    wire N__9651;
    wire N__9650;
    wire N__9649;
    wire N__9642;
    wire N__9641;
    wire N__9640;
    wire N__9633;
    wire N__9632;
    wire N__9631;
    wire N__9624;
    wire N__9623;
    wire N__9622;
    wire N__9615;
    wire N__9614;
    wire N__9613;
    wire N__9606;
    wire N__9605;
    wire N__9604;
    wire N__9597;
    wire N__9596;
    wire N__9595;
    wire N__9588;
    wire N__9587;
    wire N__9586;
    wire N__9579;
    wire N__9578;
    wire N__9577;
    wire N__9570;
    wire N__9569;
    wire N__9568;
    wire N__9561;
    wire N__9560;
    wire N__9559;
    wire N__9552;
    wire N__9551;
    wire N__9550;
    wire N__9543;
    wire N__9542;
    wire N__9541;
    wire N__9534;
    wire N__9533;
    wire N__9532;
    wire N__9525;
    wire N__9524;
    wire N__9523;
    wire N__9516;
    wire N__9515;
    wire N__9514;
    wire N__9507;
    wire N__9506;
    wire N__9505;
    wire N__9498;
    wire N__9497;
    wire N__9496;
    wire N__9489;
    wire N__9488;
    wire N__9487;
    wire N__9480;
    wire N__9479;
    wire N__9478;
    wire N__9471;
    wire N__9470;
    wire N__9469;
    wire N__9462;
    wire N__9461;
    wire N__9460;
    wire N__9453;
    wire N__9452;
    wire N__9451;
    wire N__9444;
    wire N__9443;
    wire N__9442;
    wire N__9435;
    wire N__9434;
    wire N__9433;
    wire N__9426;
    wire N__9425;
    wire N__9424;
    wire N__9417;
    wire N__9416;
    wire N__9415;
    wire N__9408;
    wire N__9407;
    wire N__9406;
    wire N__9399;
    wire N__9398;
    wire N__9397;
    wire N__9390;
    wire N__9389;
    wire N__9388;
    wire N__9381;
    wire N__9380;
    wire N__9379;
    wire N__9372;
    wire N__9371;
    wire N__9370;
    wire N__9363;
    wire N__9362;
    wire N__9361;
    wire N__9354;
    wire N__9353;
    wire N__9352;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9328;
    wire N__9325;
    wire N__9322;
    wire N__9317;
    wire N__9314;
    wire N__9311;
    wire N__9308;
    wire N__9305;
    wire N__9302;
    wire N__9299;
    wire N__9298;
    wire N__9295;
    wire N__9292;
    wire N__9287;
    wire N__9284;
    wire N__9283;
    wire N__9282;
    wire N__9281;
    wire N__9280;
    wire N__9279;
    wire N__9278;
    wire N__9277;
    wire N__9276;
    wire N__9275;
    wire N__9274;
    wire N__9273;
    wire N__9272;
    wire N__9271;
    wire N__9270;
    wire N__9269;
    wire N__9268;
    wire N__9267;
    wire N__9266;
    wire N__9265;
    wire N__9264;
    wire N__9263;
    wire N__9262;
    wire N__9261;
    wire N__9260;
    wire N__9259;
    wire N__9258;
    wire N__9257;
    wire N__9256;
    wire N__9255;
    wire N__9254;
    wire N__9253;
    wire N__9252;
    wire N__9251;
    wire N__9250;
    wire N__9249;
    wire N__9248;
    wire N__9247;
    wire N__9246;
    wire N__9245;
    wire N__9242;
    wire N__9241;
    wire N__9240;
    wire N__9239;
    wire N__9238;
    wire N__9237;
    wire N__9236;
    wire N__9235;
    wire N__9234;
    wire N__9233;
    wire N__9232;
    wire N__9231;
    wire N__9230;
    wire N__9125;
    wire N__9122;
    wire N__9121;
    wire N__9120;
    wire N__9119;
    wire N__9118;
    wire N__9117;
    wire N__9116;
    wire N__9113;
    wire N__9112;
    wire N__9111;
    wire N__9110;
    wire N__9107;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9085;
    wire N__9082;
    wire N__9081;
    wire N__9080;
    wire N__9079;
    wire N__9078;
    wire N__9077;
    wire N__9076;
    wire N__9073;
    wire N__9072;
    wire N__9071;
    wire N__9070;
    wire N__9069;
    wire N__9068;
    wire N__9067;
    wire N__9066;
    wire N__9065;
    wire N__9064;
    wire N__9063;
    wire N__9062;
    wire N__9061;
    wire N__9060;
    wire N__9059;
    wire N__9058;
    wire N__9057;
    wire N__9056;
    wire N__9055;
    wire N__9054;
    wire N__9053;
    wire N__9052;
    wire N__9051;
    wire N__9048;
    wire N__9045;
    wire N__9044;
    wire N__9043;
    wire N__9042;
    wire N__9041;
    wire N__9038;
    wire N__9037;
    wire N__9036;
    wire N__9035;
    wire N__9034;
    wire N__9033;
    wire N__9030;
    wire N__9027;
    wire N__9026;
    wire N__9025;
    wire N__9024;
    wire N__9023;
    wire N__9022;
    wire N__9019;
    wire N__9018;
    wire N__9015;
    wire N__9014;
    wire N__9013;
    wire N__9012;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8894;
    wire N__8891;
    wire N__8888;
    wire N__8885;
    wire N__8882;
    wire N__8879;
    wire N__8876;
    wire N__8873;
    wire N__8870;
    wire N__8867;
    wire N__8864;
    wire N__8863;
    wire N__8862;
    wire N__8861;
    wire N__8858;
    wire N__8857;
    wire N__8856;
    wire N__8853;
    wire N__8852;
    wire N__8851;
    wire N__8850;
    wire N__8849;
    wire N__8848;
    wire N__8845;
    wire N__8844;
    wire N__8843;
    wire N__8842;
    wire N__8841;
    wire N__8840;
    wire N__8839;
    wire N__8838;
    wire N__8835;
    wire N__8832;
    wire N__8827;
    wire N__8826;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8802;
    wire N__8797;
    wire N__8796;
    wire N__8795;
    wire N__8794;
    wire N__8791;
    wire N__8788;
    wire N__8787;
    wire N__8784;
    wire N__8777;
    wire N__8774;
    wire N__8769;
    wire N__8768;
    wire N__8767;
    wire N__8766;
    wire N__8765;
    wire N__8764;
    wire N__8761;
    wire N__8758;
    wire N__8755;
    wire N__8750;
    wire N__8745;
    wire N__8742;
    wire N__8737;
    wire N__8734;
    wire N__8727;
    wire N__8724;
    wire N__8721;
    wire N__8718;
    wire N__8711;
    wire N__8704;
    wire N__8699;
    wire N__8690;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8653;
    wire N__8650;
    wire N__8647;
    wire N__8646;
    wire N__8645;
    wire N__8640;
    wire N__8637;
    wire N__8634;
    wire N__8633;
    wire N__8628;
    wire N__8625;
    wire N__8622;
    wire N__8621;
    wire N__8618;
    wire N__8617;
    wire N__8616;
    wire N__8613;
    wire N__8610;
    wire N__8607;
    wire N__8604;
    wire N__8601;
    wire N__8598;
    wire N__8585;
    wire N__8584;
    wire N__8583;
    wire N__8582;
    wire N__8581;
    wire N__8578;
    wire N__8577;
    wire N__8576;
    wire N__8575;
    wire N__8574;
    wire N__8569;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8557;
    wire N__8556;
    wire N__8553;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8538;
    wire N__8535;
    wire N__8532;
    wire N__8529;
    wire N__8526;
    wire N__8523;
    wire N__8518;
    wire N__8511;
    wire N__8510;
    wire N__8509;
    wire N__8506;
    wire N__8503;
    wire N__8500;
    wire N__8495;
    wire N__8492;
    wire N__8487;
    wire N__8474;
    wire N__8473;
    wire N__8472;
    wire N__8471;
    wire N__8470;
    wire N__8467;
    wire N__8464;
    wire N__8463;
    wire N__8462;
    wire N__8461;
    wire N__8458;
    wire N__8455;
    wire N__8454;
    wire N__8451;
    wire N__8446;
    wire N__8443;
    wire N__8442;
    wire N__8437;
    wire N__8434;
    wire N__8433;
    wire N__8430;
    wire N__8427;
    wire N__8424;
    wire N__8421;
    wire N__8418;
    wire N__8417;
    wire N__8416;
    wire N__8413;
    wire N__8410;
    wire N__8407;
    wire N__8404;
    wire N__8401;
    wire N__8398;
    wire N__8395;
    wire N__8390;
    wire N__8389;
    wire N__8386;
    wire N__8383;
    wire N__8380;
    wire N__8375;
    wire N__8370;
    wire N__8365;
    wire N__8362;
    wire N__8357;
    wire N__8342;
    wire N__8341;
    wire N__8338;
    wire N__8335;
    wire N__8330;
    wire N__8327;
    wire N__8324;
    wire N__8323;
    wire N__8320;
    wire N__8317;
    wire N__8314;
    wire N__8311;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8299;
    wire N__8294;
    wire N__8291;
    wire N__8288;
    wire N__8285;
    wire N__8282;
    wire N__8281;
    wire N__8280;
    wire N__8279;
    wire N__8276;
    wire N__8273;
    wire N__8270;
    wire N__8267;
    wire N__8266;
    wire N__8263;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8251;
    wire N__8250;
    wire N__8247;
    wire N__8244;
    wire N__8241;
    wire N__8238;
    wire N__8235;
    wire N__8232;
    wire N__8219;
    wire N__8216;
    wire N__8215;
    wire N__8212;
    wire N__8209;
    wire N__8206;
    wire N__8203;
    wire N__8200;
    wire N__8197;
    wire N__8194;
    wire N__8191;
    wire N__8188;
    wire N__8185;
    wire N__8180;
    wire N__8177;
    wire N__8176;
    wire N__8173;
    wire N__8170;
    wire N__8167;
    wire N__8164;
    wire N__8161;
    wire N__8158;
    wire N__8155;
    wire N__8152;
    wire N__8147;
    wire N__8144;
    wire N__8141;
    wire N__8138;
    wire N__8135;
    wire N__8134;
    wire N__8133;
    wire N__8130;
    wire N__8129;
    wire N__8126;
    wire N__8125;
    wire N__8124;
    wire N__8123;
    wire N__8120;
    wire N__8119;
    wire N__8118;
    wire N__8117;
    wire N__8116;
    wire N__8115;
    wire N__8114;
    wire N__8111;
    wire N__8108;
    wire N__8105;
    wire N__8102;
    wire N__8099;
    wire N__8096;
    wire N__8093;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8067;
    wire N__8062;
    wire N__8061;
    wire N__8060;
    wire N__8057;
    wire N__8054;
    wire N__8051;
    wire N__8048;
    wire N__8045;
    wire N__8042;
    wire N__8039;
    wire N__8036;
    wire N__8029;
    wire N__8026;
    wire N__8025;
    wire N__8022;
    wire N__8017;
    wire N__8012;
    wire N__8005;
    wire N__8002;
    wire N__7999;
    wire N__7994;
    wire N__7979;
    wire N__7976;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7957;
    wire N__7956;
    wire N__7953;
    wire N__7950;
    wire N__7947;
    wire N__7942;
    wire N__7941;
    wire N__7938;
    wire N__7935;
    wire N__7932;
    wire N__7931;
    wire N__7928;
    wire N__7925;
    wire N__7922;
    wire N__7919;
    wire N__7910;
    wire N__7907;
    wire N__7904;
    wire N__7901;
    wire N__7900;
    wire N__7897;
    wire N__7894;
    wire N__7889;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7877;
    wire N__7874;
    wire N__7871;
    wire N__7868;
    wire N__7865;
    wire N__7864;
    wire N__7861;
    wire N__7858;
    wire N__7853;
    wire N__7850;
    wire N__7847;
    wire N__7844;
    wire N__7841;
    wire N__7838;
    wire N__7835;
    wire N__7832;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7816;
    wire N__7813;
    wire N__7810;
    wire N__7805;
    wire N__7802;
    wire N__7799;
    wire N__7796;
    wire N__7793;
    wire N__7790;
    wire N__7789;
    wire N__7786;
    wire N__7783;
    wire N__7780;
    wire N__7777;
    wire N__7774;
    wire N__7771;
    wire N__7768;
    wire N__7765;
    wire N__7762;
    wire N__7757;
    wire N__7754;
    wire N__7751;
    wire N__7750;
    wire N__7749;
    wire N__7746;
    wire N__7743;
    wire N__7740;
    wire N__7733;
    wire N__7732;
    wire N__7729;
    wire N__7726;
    wire N__7721;
    wire N__7718;
    wire N__7717;
    wire N__7714;
    wire N__7711;
    wire N__7706;
    wire N__7703;
    wire N__7700;
    wire N__7697;
    wire N__7694;
    wire N__7691;
    wire N__7688;
    wire N__7685;
    wire N__7682;
    wire N__7679;
    wire N__7676;
    wire N__7673;
    wire N__7670;
    wire N__7667;
    wire N__7664;
    wire N__7661;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7637;
    wire N__7634;
    wire N__7631;
    wire N__7628;
    wire N__7627;
    wire N__7626;
    wire N__7623;
    wire N__7618;
    wire N__7613;
    wire N__7610;
    wire N__7607;
    wire N__7604;
    wire N__7601;
    wire N__7598;
    wire N__7597;
    wire N__7596;
    wire N__7593;
    wire N__7592;
    wire N__7589;
    wire N__7586;
    wire N__7583;
    wire N__7580;
    wire N__7575;
    wire N__7572;
    wire N__7567;
    wire N__7566;
    wire N__7565;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7544;
    wire N__7541;
    wire N__7538;
    wire N__7535;
    wire N__7532;
    wire N__7529;
    wire N__7526;
    wire N__7523;
    wire N__7520;
    wire N__7517;
    wire N__7514;
    wire N__7511;
    wire N__7508;
    wire N__7507;
    wire N__7504;
    wire N__7501;
    wire N__7500;
    wire N__7497;
    wire N__7494;
    wire N__7491;
    wire N__7490;
    wire N__7487;
    wire N__7482;
    wire N__7479;
    wire N__7472;
    wire N__7471;
    wire N__7470;
    wire N__7469;
    wire N__7466;
    wire N__7465;
    wire N__7462;
    wire N__7461;
    wire N__7460;
    wire N__7457;
    wire N__7454;
    wire N__7451;
    wire N__7444;
    wire N__7441;
    wire N__7440;
    wire N__7439;
    wire N__7434;
    wire N__7429;
    wire N__7426;
    wire N__7423;
    wire N__7420;
    wire N__7417;
    wire N__7406;
    wire N__7403;
    wire N__7400;
    wire N__7397;
    wire N__7394;
    wire N__7391;
    wire N__7388;
    wire N__7385;
    wire N__7384;
    wire N__7381;
    wire N__7378;
    wire N__7375;
    wire N__7372;
    wire N__7369;
    wire N__7366;
    wire N__7363;
    wire N__7358;
    wire N__7355;
    wire N__7352;
    wire N__7349;
    wire N__7346;
    wire N__7343;
    wire N__7340;
    wire N__7337;
    wire N__7334;
    wire N__7331;
    wire N__7328;
    wire N__7325;
    wire N__7322;
    wire N__7319;
    wire N__7316;
    wire N__7313;
    wire N__7310;
    wire N__7307;
    wire N__7304;
    wire N__7301;
    wire N__7298;
    wire N__7295;
    wire N__7292;
    wire N__7289;
    wire N__7286;
    wire N__7283;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7271;
    wire N__7268;
    wire N__7265;
    wire N__7262;
    wire N__7259;
    wire N__7256;
    wire N__7253;
    wire N__7250;
    wire N__7247;
    wire N__7244;
    wire N__7241;
    wire N__7238;
    wire N__7235;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7223;
    wire N__7220;
    wire N__7217;
    wire N__7214;
    wire N__7211;
    wire N__7208;
    wire N__7205;
    wire N__7202;
    wire N__7199;
    wire N__7196;
    wire N__7193;
    wire N__7190;
    wire N__7187;
    wire N__7184;
    wire N__7181;
    wire N__7178;
    wire N__7175;
    wire N__7172;
    wire N__7169;
    wire N__7166;
    wire N__7163;
    wire N__7160;
    wire N__7157;
    wire N__7154;
    wire N__7151;
    wire N__7148;
    wire N__7145;
    wire N__7142;
    wire N__7139;
    wire N__7136;
    wire N__7135;
    wire N__7134;
    wire N__7133;
    wire N__7132;
    wire N__7129;
    wire N__7126;
    wire N__7123;
    wire N__7120;
    wire N__7117;
    wire N__7112;
    wire N__7109;
    wire N__7106;
    wire N__7103;
    wire N__7100;
    wire N__7095;
    wire N__7088;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7078;
    wire N__7075;
    wire N__7074;
    wire N__7071;
    wire N__7068;
    wire N__7065;
    wire N__7062;
    wire N__7057;
    wire N__7054;
    wire N__7051;
    wire N__7048;
    wire N__7045;
    wire N__7040;
    wire N__7037;
    wire N__7034;
    wire N__7031;
    wire N__7028;
    wire N__7025;
    wire N__7022;
    wire N__7019;
    wire N__7016;
    wire N__7015;
    wire N__7014;
    wire N__7011;
    wire N__7008;
    wire N__7005;
    wire N__7000;
    wire N__6999;
    wire N__6996;
    wire N__6993;
    wire N__6990;
    wire N__6983;
    wire N__6982;
    wire N__6981;
    wire N__6978;
    wire N__6977;
    wire N__6976;
    wire N__6973;
    wire N__6972;
    wire N__6971;
    wire N__6970;
    wire N__6967;
    wire N__6964;
    wire N__6961;
    wire N__6958;
    wire N__6955;
    wire N__6952;
    wire N__6947;
    wire N__6932;
    wire N__6929;
    wire N__6926;
    wire N__6923;
    wire N__6920;
    wire N__6917;
    wire N__6914;
    wire N__6911;
    wire N__6908;
    wire N__6905;
    wire N__6902;
    wire N__6899;
    wire N__6896;
    wire N__6893;
    wire N__6890;
    wire N__6887;
    wire N__6884;
    wire N__6881;
    wire N__6878;
    wire N__6875;
    wire N__6872;
    wire N__6869;
    wire N__6866;
    wire N__6863;
    wire N__6860;
    wire N__6857;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6845;
    wire N__6842;
    wire N__6839;
    wire N__6836;
    wire N__6833;
    wire N__6830;
    wire N__6827;
    wire N__6824;
    wire N__6821;
    wire N__6818;
    wire N__6815;
    wire N__6812;
    wire N__6809;
    wire N__6806;
    wire N__6803;
    wire N__6800;
    wire N__6797;
    wire N__6794;
    wire N__6791;
    wire N__6788;
    wire N__6785;
    wire N__6782;
    wire N__6779;
    wire N__6776;
    wire N__6773;
    wire N__6770;
    wire N__6767;
    wire N__6764;
    wire N__6761;
    wire N__6758;
    wire N__6757;
    wire N__6756;
    wire N__6753;
    wire N__6750;
    wire N__6747;
    wire N__6746;
    wire N__6745;
    wire N__6740;
    wire N__6737;
    wire N__6736;
    wire N__6731;
    wire N__6728;
    wire N__6725;
    wire N__6722;
    wire N__6719;
    wire N__6712;
    wire N__6709;
    wire N__6706;
    wire N__6703;
    wire N__6700;
    wire N__6695;
    wire N__6692;
    wire N__6689;
    wire N__6686;
    wire N__6683;
    wire N__6682;
    wire N__6679;
    wire N__6678;
    wire N__6675;
    wire N__6672;
    wire N__6669;
    wire N__6666;
    wire N__6659;
    wire N__6656;
    wire N__6653;
    wire N__6650;
    wire N__6647;
    wire N__6644;
    wire N__6641;
    wire N__6638;
    wire N__6635;
    wire N__6632;
    wire N__6631;
    wire N__6630;
    wire N__6629;
    wire N__6628;
    wire N__6627;
    wire N__6626;
    wire N__6625;
    wire N__6624;
    wire N__6621;
    wire N__6618;
    wire N__6609;
    wire N__6606;
    wire N__6603;
    wire N__6600;
    wire N__6591;
    wire N__6588;
    wire N__6587;
    wire N__6584;
    wire N__6581;
    wire N__6578;
    wire N__6575;
    wire N__6570;
    wire N__6565;
    wire N__6562;
    wire N__6559;
    wire N__6554;
    wire N__6551;
    wire N__6548;
    wire N__6545;
    wire N__6542;
    wire N__6539;
    wire N__6536;
    wire N__6533;
    wire N__6530;
    wire N__6527;
    wire N__6524;
    wire N__6521;
    wire N__6520;
    wire N__6517;
    wire N__6514;
    wire N__6511;
    wire N__6508;
    wire N__6507;
    wire N__6502;
    wire N__6501;
    wire N__6500;
    wire N__6497;
    wire N__6494;
    wire N__6489;
    wire N__6482;
    wire N__6479;
    wire N__6476;
    wire N__6473;
    wire N__6470;
    wire N__6467;
    wire N__6464;
    wire N__6461;
    wire N__6458;
    wire N__6455;
    wire N__6452;
    wire N__6449;
    wire N__6446;
    wire N__6443;
    wire N__6440;
    wire N__6437;
    wire N__6436;
    wire N__6433;
    wire N__6430;
    wire N__6427;
    wire N__6424;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6412;
    wire N__6409;
    wire N__6406;
    wire N__6401;
    wire N__6398;
    wire N__6395;
    wire N__6392;
    wire N__6389;
    wire N__6386;
    wire N__6383;
    wire N__6382;
    wire N__6379;
    wire N__6376;
    wire N__6371;
    wire N__6368;
    wire N__6365;
    wire N__6362;
    wire N__6361;
    wire N__6358;
    wire N__6355;
    wire N__6350;
    wire N__6347;
    wire N__6344;
    wire N__6343;
    wire N__6340;
    wire N__6337;
    wire N__6334;
    wire N__6331;
    wire N__6328;
    wire N__6325;
    wire N__6320;
    wire N__6317;
    wire N__6314;
    wire N__6311;
    wire N__6308;
    wire N__6305;
    wire N__6302;
    wire N__6301;
    wire N__6298;
    wire N__6295;
    wire N__6292;
    wire N__6287;
    wire N__6284;
    wire N__6283;
    wire N__6282;
    wire N__6279;
    wire N__6276;
    wire N__6275;
    wire N__6274;
    wire N__6273;
    wire N__6272;
    wire N__6271;
    wire N__6270;
    wire N__6269;
    wire N__6268;
    wire N__6265;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6249;
    wire N__6246;
    wire N__6243;
    wire N__6238;
    wire N__6221;
    wire N__6220;
    wire N__6217;
    wire N__6214;
    wire N__6211;
    wire N__6208;
    wire N__6205;
    wire N__6204;
    wire N__6203;
    wire N__6202;
    wire N__6201;
    wire N__6200;
    wire N__6199;
    wire N__6198;
    wire N__6197;
    wire N__6194;
    wire N__6191;
    wire N__6188;
    wire N__6185;
    wire N__6182;
    wire N__6179;
    wire N__6176;
    wire N__6173;
    wire N__6168;
    wire N__6149;
    wire N__6148;
    wire N__6147;
    wire N__6144;
    wire N__6143;
    wire N__6140;
    wire N__6137;
    wire N__6134;
    wire N__6133;
    wire N__6132;
    wire N__6131;
    wire N__6128;
    wire N__6125;
    wire N__6122;
    wire N__6119;
    wire N__6114;
    wire N__6111;
    wire N__6098;
    wire N__6097;
    wire N__6094;
    wire N__6093;
    wire N__6090;
    wire N__6087;
    wire N__6086;
    wire N__6085;
    wire N__6082;
    wire N__6079;
    wire N__6076;
    wire N__6071;
    wire N__6062;
    wire N__6061;
    wire N__6060;
    wire N__6059;
    wire N__6058;
    wire N__6057;
    wire N__6056;
    wire N__6053;
    wire N__6052;
    wire N__6051;
    wire N__6046;
    wire N__6045;
    wire N__6044;
    wire N__6043;
    wire N__6042;
    wire N__6041;
    wire N__6040;
    wire N__6039;
    wire N__6038;
    wire N__6035;
    wire N__6030;
    wire N__6027;
    wire N__6024;
    wire N__6019;
    wire N__6016;
    wire N__6011;
    wire N__6006;
    wire N__6003;
    wire N__5996;
    wire N__5991;
    wire N__5972;
    wire N__5971;
    wire N__5970;
    wire N__5969;
    wire N__5968;
    wire N__5967;
    wire N__5966;
    wire N__5965;
    wire N__5964;
    wire N__5963;
    wire N__5962;
    wire N__5959;
    wire N__5958;
    wire N__5953;
    wire N__5952;
    wire N__5951;
    wire N__5946;
    wire N__5945;
    wire N__5944;
    wire N__5943;
    wire N__5940;
    wire N__5933;
    wire N__5932;
    wire N__5929;
    wire N__5924;
    wire N__5921;
    wire N__5918;
    wire N__5913;
    wire N__5910;
    wire N__5907;
    wire N__5902;
    wire N__5897;
    wire N__5894;
    wire N__5873;
    wire N__5870;
    wire N__5867;
    wire N__5866;
    wire N__5863;
    wire N__5862;
    wire N__5861;
    wire N__5860;
    wire N__5859;
    wire N__5856;
    wire N__5853;
    wire N__5850;
    wire N__5843;
    wire N__5834;
    wire N__5831;
    wire N__5828;
    wire N__5827;
    wire N__5824;
    wire N__5821;
    wire N__5816;
    wire N__5813;
    wire N__5810;
    wire N__5807;
    wire N__5804;
    wire N__5801;
    wire N__5798;
    wire N__5795;
    wire N__5792;
    wire N__5789;
    wire N__5786;
    wire N__5783;
    wire N__5780;
    wire N__5777;
    wire N__5774;
    wire N__5771;
    wire N__5768;
    wire N__5765;
    wire N__5764;
    wire N__5763;
    wire N__5762;
    wire N__5759;
    wire N__5758;
    wire N__5757;
    wire N__5756;
    wire N__5755;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5732;
    wire N__5717;
    wire N__5714;
    wire N__5713;
    wire N__5710;
    wire N__5707;
    wire N__5704;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5681;
    wire N__5680;
    wire N__5677;
    wire N__5674;
    wire N__5671;
    wire N__5666;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5654;
    wire N__5651;
    wire N__5648;
    wire N__5645;
    wire N__5644;
    wire N__5641;
    wire N__5638;
    wire N__5635;
    wire N__5630;
    wire N__5629;
    wire N__5626;
    wire N__5623;
    wire N__5618;
    wire N__5617;
    wire N__5616;
    wire N__5613;
    wire N__5608;
    wire N__5603;
    wire N__5602;
    wire N__5599;
    wire N__5596;
    wire N__5591;
    wire N__5588;
    wire N__5585;
    wire N__5584;
    wire N__5583;
    wire N__5580;
    wire N__5575;
    wire N__5570;
    wire N__5569;
    wire N__5566;
    wire N__5563;
    wire N__5560;
    wire N__5555;
    wire N__5552;
    wire N__5551;
    wire N__5548;
    wire N__5545;
    wire N__5540;
    wire N__5537;
    wire N__5534;
    wire N__5531;
    wire N__5528;
    wire N__5525;
    wire N__5522;
    wire N__5519;
    wire N__5516;
    wire N__5513;
    wire N__5510;
    wire N__5507;
    wire N__5504;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5489;
    wire N__5486;
    wire N__5483;
    wire N__5480;
    wire N__5477;
    wire N__5474;
    wire N__5471;
    wire N__5468;
    wire N__5467;
    wire N__5466;
    wire N__5463;
    wire N__5460;
    wire N__5457;
    wire N__5450;
    wire N__5449;
    wire N__5446;
    wire N__5443;
    wire N__5438;
    wire N__5435;
    wire N__5432;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5422;
    wire N__5421;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5409;
    wire N__5402;
    wire N__5399;
    wire N__5398;
    wire N__5397;
    wire N__5394;
    wire N__5389;
    wire N__5384;
    wire N__5381;
    wire N__5380;
    wire N__5379;
    wire N__5378;
    wire N__5375;
    wire N__5368;
    wire N__5363;
    wire N__5360;
    wire N__5359;
    wire N__5358;
    wire N__5357;
    wire N__5350;
    wire N__5347;
    wire N__5342;
    wire N__5339;
    wire N__5336;
    wire N__5335;
    wire N__5332;
    wire N__5329;
    wire N__5324;
    wire N__5321;
    wire N__5318;
    wire N__5315;
    wire N__5312;
    wire N__5309;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5288;
    wire N__5285;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5243;
    wire N__5240;
    wire N__5237;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5222;
    wire N__5219;
    wire N__5216;
    wire N__5213;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5203;
    wire N__5200;
    wire N__5197;
    wire N__5192;
    wire N__5189;
    wire N__5186;
    wire N__5183;
    wire N__5182;
    wire N__5181;
    wire N__5180;
    wire N__5173;
    wire N__5170;
    wire N__5165;
    wire N__5164;
    wire N__5161;
    wire N__5158;
    wire N__5155;
    wire N__5152;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5137;
    wire N__5136;
    wire N__5135;
    wire N__5132;
    wire N__5125;
    wire N__5120;
    wire N__5117;
    wire N__5114;
    wire N__5113;
    wire N__5110;
    wire N__5109;
    wire N__5106;
    wire N__5105;
    wire N__5102;
    wire N__5095;
    wire N__5090;
    wire N__5087;
    wire N__5084;
    wire N__5081;
    wire N__5078;
    wire N__5075;
    wire N__5072;
    wire N__5069;
    wire N__5066;
    wire N__5063;
    wire N__5060;
    wire N__5057;
    wire N__5054;
    wire N__5051;
    wire N__5048;
    wire N__5045;
    wire N__5042;
    wire N__5039;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5027;
    wire N__5024;
    wire N__5023;
    wire N__5020;
    wire N__5017;
    wire N__5012;
    wire N__5011;
    wire N__5008;
    wire N__5005;
    wire N__5000;
    wire N__4999;
    wire N__4996;
    wire N__4993;
    wire N__4990;
    wire N__4985;
    wire N__4984;
    wire N__4981;
    wire N__4978;
    wire N__4973;
    wire N__4972;
    wire N__4969;
    wire N__4966;
    wire N__4961;
    wire N__4960;
    wire N__4957;
    wire N__4954;
    wire N__4949;
    wire N__4946;
    wire N__4943;
    wire N__4942;
    wire N__4939;
    wire N__4936;
    wire N__4933;
    wire N__4930;
    wire N__4927;
    wire N__4924;
    wire N__4919;
    wire N__4916;
    wire N__4913;
    wire N__4912;
    wire N__4909;
    wire N__4906;
    wire N__4905;
    wire N__4900;
    wire N__4897;
    wire N__4894;
    wire N__4891;
    wire N__4888;
    wire N__4885;
    wire N__4882;
    wire N__4879;
    wire N__4876;
    wire N__4871;
    wire N__4870;
    wire N__4867;
    wire N__4866;
    wire N__4863;
    wire N__4860;
    wire N__4857;
    wire N__4850;
    wire N__4849;
    wire N__4846;
    wire N__4845;
    wire N__4840;
    wire N__4839;
    wire N__4836;
    wire N__4833;
    wire N__4830;
    wire N__4827;
    wire N__4820;
    wire N__4819;
    wire N__4814;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4793;
    wire N__4790;
    wire N__4787;
    wire N__4784;
    wire N__4781;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4753;
    wire N__4752;
    wire N__4749;
    wire N__4746;
    wire N__4743;
    wire N__4736;
    wire N__4735;
    wire N__4734;
    wire N__4731;
    wire N__4728;
    wire N__4723;
    wire N__4720;
    wire N__4715;
    wire N__4712;
    wire N__4709;
    wire N__4706;
    wire N__4703;
    wire N__4700;
    wire N__4697;
    wire N__4694;
    wire N__4693;
    wire N__4690;
    wire N__4689;
    wire N__4686;
    wire N__4683;
    wire N__4680;
    wire N__4677;
    wire N__4670;
    wire N__4669;
    wire N__4666;
    wire N__4663;
    wire N__4658;
    wire N__4655;
    wire N__4652;
    wire N__4649;
    wire N__4648;
    wire N__4645;
    wire N__4644;
    wire N__4641;
    wire N__4638;
    wire N__4635;
    wire N__4632;
    wire N__4629;
    wire N__4624;
    wire N__4621;
    wire N__4618;
    wire N__4615;
    wire N__4612;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4586;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4562;
    wire N__4559;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4541;
    wire N__4540;
    wire N__4537;
    wire N__4534;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4522;
    wire N__4519;
    wire N__4516;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire N__4498;
    wire N__4495;
    wire N__4492;
    wire N__4487;
    wire N__4484;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4474;
    wire N__4471;
    wire N__4468;
    wire N__4467;
    wire N__4464;
    wire N__4461;
    wire N__4458;
    wire N__4451;
    wire N__4450;
    wire N__4449;
    wire N__4446;
    wire N__4443;
    wire N__4440;
    wire N__4437;
    wire N__4434;
    wire N__4431;
    wire N__4424;
    wire N__4423;
    wire N__4420;
    wire N__4417;
    wire N__4412;
    wire N__4411;
    wire N__4410;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4395;
    wire N__4392;
    wire N__4389;
    wire N__4386;
    wire N__4383;
    wire N__4378;
    wire N__4375;
    wire N__4372;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4360;
    wire N__4355;
    wire N__4354;
    wire N__4353;
    wire N__4350;
    wire N__4345;
    wire N__4340;
    wire N__4337;
    wire N__4336;
    wire N__4333;
    wire N__4330;
    wire N__4325;
    wire N__4322;
    wire N__4319;
    wire N__4316;
    wire N__4315;
    wire N__4312;
    wire N__4309;
    wire N__4304;
    wire N__4301;
    wire N__4298;
    wire N__4295;
    wire N__4292;
    wire N__4289;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4277;
    wire N__4276;
    wire N__4273;
    wire N__4270;
    wire N__4265;
    wire N__4264;
    wire N__4261;
    wire N__4258;
    wire N__4257;
    wire N__4252;
    wire N__4249;
    wire N__4244;
    wire N__4241;
    wire N__4238;
    wire N__4235;
    wire N__4232;
    wire N__4229;
    wire N__4226;
    wire N__4223;
    wire N__4220;
    wire N__4217;
    wire N__4214;
    wire N__4211;
    wire N__4208;
    wire N__4205;
    wire N__4202;
    wire N__4199;
    wire N__4196;
    wire N__4193;
    wire N__4190;
    wire N__4187;
    wire N__4184;
    wire N__4181;
    wire N__4180;
    wire N__4179;
    wire N__4178;
    wire N__4175;
    wire N__4172;
    wire N__4169;
    wire N__4166;
    wire N__4163;
    wire N__4160;
    wire N__4151;
    wire N__4150;
    wire N__4147;
    wire N__4144;
    wire N__4141;
    wire N__4140;
    wire N__4139;
    wire N__4138;
    wire N__4135;
    wire N__4134;
    wire N__4133;
    wire N__4132;
    wire N__4129;
    wire N__4126;
    wire N__4121;
    wire N__4118;
    wire N__4111;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4090;
    wire N__4089;
    wire N__4088;
    wire N__4085;
    wire N__4080;
    wire N__4077;
    wire N__4070;
    wire N__4069;
    wire N__4068;
    wire N__4063;
    wire N__4060;
    wire N__4055;
    wire N__4052;
    wire N__4049;
    wire N__4048;
    wire N__4045;
    wire N__4042;
    wire N__4037;
    wire N__4036;
    wire N__4035;
    wire N__4034;
    wire N__4033;
    wire N__4032;
    wire N__4029;
    wire N__4024;
    wire N__4021;
    wire N__4020;
    wire N__4017;
    wire N__4014;
    wire N__4009;
    wire N__4006;
    wire N__4003;
    wire N__4000;
    wire N__3989;
    wire N__3988;
    wire N__3987;
    wire N__3986;
    wire N__3985;
    wire N__3982;
    wire N__3979;
    wire N__3976;
    wire N__3973;
    wire N__3968;
    wire N__3959;
    wire N__3956;
    wire N__3953;
    wire N__3952;
    wire N__3951;
    wire N__3950;
    wire N__3949;
    wire N__3948;
    wire N__3945;
    wire N__3942;
    wire N__3939;
    wire N__3932;
    wire N__3923;
    wire N__3920;
    wire N__3917;
    wire N__3916;
    wire N__3915;
    wire N__3912;
    wire N__3909;
    wire N__3906;
    wire N__3901;
    wire N__3896;
    wire N__3893;
    wire N__3892;
    wire N__3891;
    wire N__3890;
    wire N__3887;
    wire N__3880;
    wire N__3875;
    wire N__3874;
    wire N__3871;
    wire N__3868;
    wire N__3865;
    wire N__3864;
    wire N__3861;
    wire N__3858;
    wire N__3855;
    wire N__3848;
    wire N__3845;
    wire N__3842;
    wire N__3839;
    wire N__3836;
    wire N__3833;
    wire N__3830;
    wire N__3827;
    wire N__3826;
    wire N__3823;
    wire N__3820;
    wire N__3815;
    wire N__3814;
    wire N__3811;
    wire N__3810;
    wire N__3807;
    wire N__3806;
    wire N__3803;
    wire N__3800;
    wire N__3797;
    wire N__3794;
    wire N__3785;
    wire N__3782;
    wire N__3779;
    wire N__3776;
    wire N__3773;
    wire N__3770;
    wire N__3769;
    wire N__3766;
    wire N__3763;
    wire N__3758;
    wire N__3755;
    wire N__3752;
    wire N__3749;
    wire N__3746;
    wire N__3745;
    wire N__3742;
    wire N__3741;
    wire N__3738;
    wire N__3735;
    wire N__3732;
    wire N__3725;
    wire N__3722;
    wire N__3721;
    wire N__3720;
    wire N__3713;
    wire N__3710;
    wire N__3709;
    wire N__3704;
    wire N__3701;
    wire N__3700;
    wire N__3699;
    wire N__3696;
    wire N__3693;
    wire N__3690;
    wire N__3683;
    wire N__3680;
    wire N__3677;
    wire N__3676;
    wire N__3673;
    wire N__3670;
    wire N__3667;
    wire N__3664;
    wire N__3661;
    wire N__3658;
    wire N__3653;
    wire N__3650;
    wire N__3647;
    wire N__3644;
    wire N__3641;
    wire N__3640;
    wire N__3639;
    wire N__3636;
    wire N__3631;
    wire N__3626;
    wire N__3623;
    wire N__3620;
    wire N__3617;
    wire N__3614;
    wire N__3611;
    wire N__3608;
    wire N__3607;
    wire N__3604;
    wire N__3601;
    wire N__3596;
    wire N__3593;
    wire N__3590;
    wire N__3587;
    wire N__3584;
    wire N__3581;
    wire N__3578;
    wire N__3575;
    wire N__3572;
    wire N__3569;
    wire N__3566;
    wire N__3563;
    wire N__3562;
    wire N__3559;
    wire N__3556;
    wire N__3553;
    wire N__3550;
    wire N__3547;
    wire N__3544;
    wire N__3541;
    wire N__3538;
    wire N__3535;
    wire N__3532;
    wire N__3531;
    wire N__3526;
    wire N__3523;
    wire N__3518;
    wire N__3515;
    wire N__3512;
    wire N__3509;
    wire N__3506;
    wire N__3503;
    wire N__3500;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire CLK40_OUT_i_i;
    wire CLK80_OUT_i_i;
    wire ASn_c;
    wire \U712_REG_SM.REG_TACK_7_0_cascade_ ;
    wire \U712_REG_SM.un1_STATE_COUNT_5_0_1 ;
    wire \U712_REG_SM.N_183_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_6 ;
    wire \U712_REG_SM.DS_EN_0_sqmuxa_1_0_a3_0_cascade_ ;
    wire C1_c;
    wire \U712_REG_SM.N_162_0_cascade_ ;
    wire \U712_REG_SM.N_166_0 ;
    wire C3_c;
    wire VBENn_c;
    wire \U712_REG_SM.N_162_0 ;
    wire \U712_REG_SM.N_171_0_cascade_ ;
    wire \U712_REG_SM.RnW_m ;
    wire \U712_REG_SM.un1_LDS_OUT_0_sqmuxa_1_0_cascade_ ;
    wire \U712_REG_SM.N_165_0 ;
    wire \U712_REG_SM.N_167_0_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_2 ;
    wire \U712_REG_SM.N_167_0 ;
    wire \U712_REG_SM.N_176_0_cascade_ ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_2 ;
    wire \U712_REG_SM.N_157_0 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_2 ;
    wire \U712_REG_SM.N_157_0_cascade_ ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire \U712_REG_SM.N_176_0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_5 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_REG_SM.N_192 ;
    wire TACK_OUTn;
    wire \U712_REG_SM.N_171_0 ;
    wire \U712_REG_SM.UDS_OUT_2_0_0 ;
    wire \U712_REG_SM.LDS_OUTZ0 ;
    wire U712_REG_SM_un1_LDSn_i;
    wire \U712_REG_SM.UDS_OUTZ0 ;
    wire \U712_REG_SM.DS_ENZ0 ;
    wire U712_REG_SM_un1_UDSn_i;
    wire A_c_13;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_4_cascade_ ;
    wire A_c_6;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \U712_REG_SM.N_163_0 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_REG_SM.N_186 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_1 ;
    wire \U712_REG_SM.N_188 ;
    wire REG_TACK;
    wire \U712_CYCLE_TERM.TACK_EN6_0_cascade_ ;
    wire \U712_CYCLE_TERM.N_45_0_0_en_cascade_ ;
    wire REGSPACEn_c;
    wire \U712_REG_SM.DS_EN_0_sqmuxa_1 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_0 ;
    wire CPU_TACKm;
    wire CLK40_OUT_i;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire DBRn_c;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_CYCLE_TERM.N_45_0_0_en_0 ;
    wire \U712_REG_SM.LDS_OUT_2_0_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_2 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0 ;
    wire SIZ_c_0;
    wire TACK_EN_i_ess;
    wire N_614_i;
    wire \U712_CHIP_RAM.N_36 ;
    wire CMA_c_4;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire bfn_10_7_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire C1_c_g;
    wire \U712_CHIP_RAM.N_49_cascade_ ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_a2_0_0_cascade_ ;
    wire RAMENn_c;
    wire TSn_c;
    wire U712_REG_SM_DBR_SYNC_1;
    wire U712_REG_SM_DBR_SYNC_0;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_57_cascade_ ;
    wire \U712_CHIP_RAM.N_58_cascade_ ;
    wire \U712_CHIP_RAM.N_40_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_0 ;
    wire \U712_CHIP_RAM.N_99_cascade_ ;
    wire \U712_CHIP_RAM.N_85 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_a2_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_a2_0_0 ;
    wire \U712_CHIP_RAM.N_65_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_ ;
    wire \U712_CHIP_RAM.N_58 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_a2_0_cascade_ ;
    wire SIZ_c_1;
    wire A_c_0;
    wire \U712_BYTE_ENABLE.LLBE_0_0_tz ;
    wire \U712_BYTE_ENABLE.LW_TRANS_0 ;
    wire \U712_BYTE_ENABLE.LLBE_0_0_tz_cascade_ ;
    wire A_c_1;
    wire CMA_c_2;
    wire A_c_4;
    wire A_c_11;
    wire \U712_CHIP_RAM.N_34 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_2 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_CHIP_RAM.N_74_cascade_ ;
    wire \U712_CHIP_RAM.N_50_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_75 ;
    wire \U712_CHIP_RAM.N_60 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_1 ;
    wire \U712_CHIP_RAM.N_77 ;
    wire \U712_CHIP_RAM.N_40 ;
    wire \U712_CHIP_RAM.N_62_cascade_ ;
    wire \U712_CHIP_RAM.N_13_cascade_ ;
    wire \U712_CHIP_RAM.N_44_cascade_ ;
    wire \U712_CHIP_RAM.N_93 ;
    wire \U712_CHIP_RAM.N_13 ;
    wire \U712_CHIP_RAM.N_65 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_i_1_0_cascade_ ;
    wire \U712_CHIP_RAM.N_62 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.N_57 ;
    wire \U712_BYTE_ENABLE.un2_CLLBEnZ0 ;
    wire CLLBEn_c;
    wire \U712_CHIP_RAM.DMA_CYCLE_7 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_0 ;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.un1_CMA31_0_i ;
    wire A_c_15;
    wire A_c_8;
    wire \U712_CHIP_RAM.N_38 ;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_6 ;
    wire \U712_CHIP_RAM.N_44 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0 ;
    wire \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.REFRESH_CYCLEZ0 ;
    wire \U712_CHIP_RAM.N_47 ;
    wire \U712_CHIP_RAM.N_47_cascade_ ;
    wire \U712_CHIP_RAM.N_89 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_a2_6_0 ;
    wire \U712_CHIP_RAM.N_100 ;
    wire \U712_CHIP_RAM.N_100_cascade_ ;
    wire \U712_CHIP_RAM.N_101 ;
    wire AWEn_c;
    wire \U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_0_a2_1 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_0_cascade_ ;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.N_56 ;
    wire \U712_CHIP_RAM.N_42 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.N_42_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.N_98 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0 ;
    wire RnW_c;
    wire DBDIR_c;
    wire DRDDIR_0_i;
    wire RESETn_c;
    wire RESETn_c_i;
    wire CRCSn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CMA_c_10;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0 ;
    wire \U712_CHIP_RAM.N_45 ;
    wire A_c_16;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_7_cascade_ ;
    wire A_c_18;
    wire CMA_c_0;
    wire CMA_c_3;
    wire A_c_5;
    wire A_c_12;
    wire \U712_CHIP_RAM.N_35 ;
    wire A_c_7;
    wire A_c_14;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_5 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_3 ;
    wire A_c_3;
    wire A_c_10;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_ ;
    wire \U712_CHIP_RAM.N_33 ;
    wire A_c_9;
    wire A_c_2;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_ ;
    wire \U712_CHIP_RAM.N_32 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_BYTE_ENABLE.un2_CUMBEnZ0 ;
    wire CASLn_c;
    wire CUMBEn_c;
    wire \U712_BYTE_ENABLE.un2_CLMBEnZ0 ;
    wire CLMBEn_c;
    wire CASUn_c;
    wire DBENn_c;
    wire \U712_BYTE_ENABLE.un2_CUUBEnZ0 ;
    wire CUUBEn_c;
    wire REG_CYCLEm;
    wire DMA_CYCLEm;
    wire N_52_i;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.N_37 ;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.N_39 ;
    wire CMA_c_7;
    wire A_c_19;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ;
    wire DRA_c_6;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire DRA_c_1;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire RASn_c;
    wire WEn_c;
    wire A_c_17;
    wire CPU_CYCLEm;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.un1_CMA31_0_i_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire \U712_CHIP_RAM.CMA_5_0_8 ;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ;
    wire CONSTANT_ONE_NET;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire CASn_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_1 ;
    wire RAS0n_c;
    wire RAS1n_c;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_0 ;
    wire _gnd_net_;
    wire CLK80_OUT;
    wire RESETn_c_i_g;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_OUT_i),
            .REFERENCECLK(N__3518),
            .RESETB(N__8215),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_OUT),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__10065),
            .DIN(N__10064),
            .DOUT(N__10063),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__10065),
            .PADOUT(N__10064),
            .PADIN(N__10063),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7598),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__10056),
            .DIN(N__10055),
            .DOUT(N__10054),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__10056),
            .PADOUT(N__10055),
            .PADIN(N__10054),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__10047),
            .DIN(N__10046),
            .DOUT(N__10045),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__10047),
            .PADOUT(N__10046),
            .PADIN(N__10045),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7979),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__10038),
            .DIN(N__10037),
            .DOUT(N__10036),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__10038),
            .PADOUT(N__10037),
            .PADIN(N__10036),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6659),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__10029),
            .DIN(N__10028),
            .DOUT(N__10027),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__10029),
            .PADOUT(N__10028),
            .PADIN(N__10027),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKEN_obuf_iopad (
            .OE(N__10020),
            .DIN(N__10019),
            .DOUT(N__10018),
            .PACKAGEPIN(CLKEN));
    defparam CLKEN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKEN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKEN_obuf_preio (
            .PADOEN(N__10020),
            .PADOUT(N__10019),
            .PADIN(N__10018),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8219),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__10011),
            .DIN(N__10010),
            .DOUT(N__10009),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__10011),
            .PADOUT(N__10010),
            .PADIN(N__10009),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__10002),
            .DIN(N__10001),
            .DOUT(N__10000),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__10002),
            .PADOUT(N__10001),
            .PADIN(N__10000),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__9993),
            .DIN(N__9992),
            .DOUT(N__9991),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__9993),
            .PADOUT(N__9992),
            .PADIN(N__9991),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS1n_ibuf_iopad (
            .OE(N__9984),
            .DIN(N__9983),
            .DOUT(N__9982),
            .PACKAGEPIN(RAS1n));
    defparam RAS1n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS1n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS1n_ibuf_preio (
            .PADOEN(N__9984),
            .PADOUT(N__9983),
            .PADIN(N__9982),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS1n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__9975),
            .DIN(N__9974),
            .DOUT(N__9973),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__9975),
            .PADOUT(N__9974),
            .PADIN(N__9973),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__9966),
            .DIN(N__9965),
            .DOUT(N__9964),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__9966),
            .PADOUT(N__9965),
            .PADIN(N__9964),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7313),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuf_iopad (
            .OE(N__9957),
            .DIN(N__9956),
            .DOUT(N__9955),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMENn_obuf_preio (
            .PADOEN(N__9957),
            .PADOUT(N__9956),
            .PADIN(N__9955),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4942),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__9948),
            .DIN(N__9947),
            .DOUT(N__9946),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__9948),
            .PADOUT(N__9947),
            .PADIN(N__9946),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__9939),
            .DIN(N__9938),
            .DOUT(N__9937),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__9939),
            .PADOUT(N__9938),
            .PADIN(N__9937),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__9930),
            .DIN(N__9929),
            .DOUT(N__9928),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__9930),
            .PADOUT(N__9929),
            .PADIN(N__9928),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3785),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__9921),
            .DIN(N__9920),
            .DOUT(N__9919),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__9921),
            .PADOUT(N__9920),
            .PADIN(N__9919),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__9912),
            .DIN(N__9911),
            .DOUT(N__9910),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__9912),
            .PADOUT(N__9911),
            .PADIN(N__9910),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__9903),
            .DIN(N__9902),
            .DOUT(N__9901),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__9903),
            .PADOUT(N__9902),
            .PADIN(N__9901),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6899),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__9894),
            .DIN(N__9893),
            .DOUT(N__9892),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__9894),
            .PADOUT(N__9893),
            .PADIN(N__9892),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__9885),
            .DIN(N__9884),
            .DOUT(N__9883),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__9885),
            .PADOUT(N__9884),
            .PADIN(N__9883),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6542),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__9876),
            .DIN(N__9875),
            .DOUT(N__9874),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__9876),
            .PADOUT(N__9875),
            .PADIN(N__9874),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__9867),
            .DIN(N__9866),
            .DOUT(N__9865),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__9867),
            .PADOUT(N__9866),
            .PADIN(N__9865),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__9858),
            .DIN(N__9857),
            .DOUT(N__9856),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__9858),
            .PADOUT(N__9857),
            .PADIN(N__9856),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__9849),
            .DIN(N__9848),
            .DOUT(N__9847),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__9849),
            .PADOUT(N__9848),
            .PADIN(N__9847),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__9840),
            .DIN(N__9839),
            .DOUT(N__9838),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__9840),
            .PADOUT(N__9839),
            .PADIN(N__9838),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__9831),
            .DIN(N__9830),
            .DOUT(N__9829),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__9831),
            .PADOUT(N__9830),
            .PADIN(N__9829),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__9822),
            .DIN(N__9821),
            .DOUT(N__9820),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__9822),
            .PADOUT(N__9821),
            .PADIN(N__9820),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__9813),
            .DIN(N__9812),
            .DOUT(N__9811),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__9813),
            .PADOUT(N__9812),
            .PADIN(N__9811),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__9804),
            .DIN(N__9803),
            .DOUT(N__9802),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__9804),
            .PADOUT(N__9803),
            .PADIN(N__9802),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__9795),
            .DIN(N__9794),
            .DOUT(N__9793),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__9795),
            .PADOUT(N__9794),
            .PADIN(N__9793),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__9786),
            .DIN(N__9785),
            .DOUT(N__9784),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__9786),
            .PADOUT(N__9785),
            .PADIN(N__9784),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5501),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__9777),
            .DIN(N__9776),
            .DOUT(N__9775),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__9777),
            .PADOUT(N__9776),
            .PADIN(N__9775),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__9768),
            .DIN(N__9767),
            .DOUT(N__9766),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__9768),
            .PADOUT(N__9767),
            .PADIN(N__9766),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__9759),
            .DIN(N__9758),
            .DOUT(N__9757),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__9759),
            .PADOUT(N__9758),
            .PADIN(N__9757),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__9750),
            .DIN(N__9749),
            .DOUT(N__9748),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__9750),
            .PADOUT(N__9749),
            .PADIN(N__9748),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_obuf_iopad (
            .OE(N__9741),
            .DIN(N__9740),
            .DOUT(N__9739),
            .PACKAGEPIN(CLK40C));
    defparam CLK40C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_obuf_preio (
            .PADOEN(N__9741),
            .PADOUT(N__9740),
            .PADIN(N__9739),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3593),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__9732),
            .DIN(N__9731),
            .DOUT(N__9730),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__9732),
            .PADOUT(N__9731),
            .PADIN(N__9730),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4304),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__9723),
            .DIN(N__9722),
            .DOUT(N__9721),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__9723),
            .PADOUT(N__9722),
            .PADIN(N__9721),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__9714),
            .DIN(N__9713),
            .DOUT(N__9712),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__9714),
            .PADOUT(N__9713),
            .PADIN(N__9712),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7679),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__9705),
            .DIN(N__9704),
            .DOUT(N__9703),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__9705),
            .PADOUT(N__9704),
            .PADIN(N__9703),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__9696),
            .DIN(N__9695),
            .DOUT(N__9694),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__9696),
            .PADOUT(N__9695),
            .PADIN(N__9694),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__9687),
            .DIN(N__9686),
            .DOUT(N__9685),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__9687),
            .PADOUT(N__9686),
            .PADIN(N__9685),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3584),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__9678),
            .DIN(N__9677),
            .DOUT(N__9676),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__9678),
            .PADOUT(N__9677),
            .PADIN(N__9676),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__9669),
            .DIN(N__9668),
            .DOUT(N__9667),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__9669),
            .PADOUT(N__9668),
            .PADIN(N__9667),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3566),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__9660),
            .DIN(N__9659),
            .DOUT(N__9658),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__9660),
            .PADOUT(N__9659),
            .PADIN(N__9658),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6881),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__9651),
            .DIN(N__9650),
            .DOUT(N__9649),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__9651),
            .PADOUT(N__9650),
            .PADIN(N__9649),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__9642),
            .DIN(N__9641),
            .DOUT(N__9640),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__9642),
            .PADOUT(N__9641),
            .PADIN(N__9640),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_0_iopad (
            .OE(N__9633),
            .DIN(N__9632),
            .DOUT(N__9631),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__9633),
            .PADOUT(N__9632),
            .PADIN(N__9631),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__9624),
            .DIN(N__9623),
            .DOUT(N__9622),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__9624),
            .PADOUT(N__9623),
            .PADIN(N__9622),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6482),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__9615),
            .DIN(N__9614),
            .DOUT(N__9613),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__9615),
            .PADOUT(N__9614),
            .PADIN(N__9613),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__9606),
            .DIN(N__9605),
            .DOUT(N__9604),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__9606),
            .PADOUT(N__9605),
            .PADIN(N__9604),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4571),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__9597),
            .DIN(N__9596),
            .DOUT(N__9595),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__9597),
            .PADOUT(N__9596),
            .PADIN(N__9595),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7406),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__9588),
            .DIN(N__9587),
            .DOUT(N__9586),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__9588),
            .PADOUT(N__9587),
            .PADIN(N__9586),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5534),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__9579),
            .DIN(N__9578),
            .DOUT(N__9577),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__9579),
            .PADOUT(N__9578),
            .PADIN(N__9577),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7271),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__9570),
            .DIN(N__9569),
            .DOUT(N__9568),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__9570),
            .PADOUT(N__9569),
            .PADIN(N__9568),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3562),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__9561),
            .DIN(N__9560),
            .DOUT(N__9559),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__9561),
            .PADOUT(N__9560),
            .PADIN(N__9559),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__9552),
            .DIN(N__9551),
            .DOUT(N__9550),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__9552),
            .PADOUT(N__9551),
            .PADIN(N__9550),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__9543),
            .DIN(N__9542),
            .DOUT(N__9541),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__9543),
            .PADOUT(N__9542),
            .PADIN(N__9541),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7649),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__9534),
            .DIN(N__9533),
            .DOUT(N__9532),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__9534),
            .PADOUT(N__9533),
            .PADIN(N__9532),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8897),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__9525),
            .DIN(N__9524),
            .DOUT(N__9523),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__9525),
            .PADOUT(N__9524),
            .PADIN(N__9523),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6695),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__9516),
            .DIN(N__9515),
            .DOUT(N__9514),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__9516),
            .PADOUT(N__9515),
            .PADIN(N__9514),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7037),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__9507),
            .DIN(N__9506),
            .DOUT(N__9505),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__9507),
            .PADOUT(N__9506),
            .PADIN(N__9505),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__9498),
            .DIN(N__9497),
            .DOUT(N__9496),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__9498),
            .PADOUT(N__9497),
            .PADIN(N__9496),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__9489),
            .DIN(N__9488),
            .DOUT(N__9487),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__9489),
            .PADOUT(N__9488),
            .PADIN(N__9487),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__9480),
            .DIN(N__9479),
            .DOUT(N__9478),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__9480),
            .PADOUT(N__9479),
            .PADIN(N__9478),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__9471),
            .DIN(N__9470),
            .DOUT(N__9469),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__9471),
            .PADOUT(N__9470),
            .PADIN(N__9469),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6464),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__9462),
            .DIN(N__9461),
            .DOUT(N__9460),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__9462),
            .PADOUT(N__9461),
            .PADIN(N__9460),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__9453),
            .DIN(N__9452),
            .DOUT(N__9451),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__9453),
            .PADOUT(N__9452),
            .PADIN(N__9451),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7532),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__9444),
            .DIN(N__9443),
            .DOUT(N__9442),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__9444),
            .PADOUT(N__9443),
            .PADIN(N__9442),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4598),
            .DIN0(),
            .DOUT0(N__3842),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__9435),
            .DIN(N__9434),
            .DOUT(N__9433),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__9435),
            .PADOUT(N__9434),
            .PADIN(N__9433),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5075),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__9426),
            .DIN(N__9425),
            .DOUT(N__9424),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__9426),
            .PADOUT(N__9425),
            .PADIN(N__9424),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__9417),
            .DIN(N__9416),
            .DOUT(N__9415),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__9417),
            .PADOUT(N__9416),
            .PADIN(N__9415),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__9408),
            .DIN(N__9407),
            .DOUT(N__9406),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__9408),
            .PADOUT(N__9407),
            .PADIN(N__9406),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8675),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__9399),
            .DIN(N__9398),
            .DOUT(N__9397),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__9399),
            .PADOUT(N__9398),
            .PADIN(N__9397),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__9390),
            .DIN(N__9389),
            .DOUT(N__9388),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__9390),
            .PADOUT(N__9389),
            .PADIN(N__9388),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__9381),
            .DIN(N__9380),
            .DOUT(N__9379),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__9381),
            .PADOUT(N__9380),
            .PADIN(N__9379),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__9372),
            .DIN(N__9371),
            .DOUT(N__9370),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__9372),
            .PADOUT(N__9371),
            .PADIN(N__9370),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__9363),
            .DIN(N__9362),
            .DOUT(N__9361),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__9363),
            .PADOUT(N__9362),
            .PADIN(N__9361),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7340),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__9354),
            .DIN(N__9353),
            .DOUT(N__9352),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__9354),
            .PADOUT(N__9353),
            .PADIN(N__9352),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4244),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__2241 (
            .O(N__9335),
            .I(N__9332));
    InMux I__2240 (
            .O(N__9332),
            .I(N__9329));
    LocalMux I__2239 (
            .O(N__9329),
            .I(N__9325));
    InMux I__2238 (
            .O(N__9328),
            .I(N__9322));
    Span4Mux_h I__2237 (
            .O(N__9325),
            .I(N__9317));
    LocalMux I__2236 (
            .O(N__9322),
            .I(N__9317));
    Span4Mux_v I__2235 (
            .O(N__9317),
            .I(N__9314));
    Sp12to4 I__2234 (
            .O(N__9314),
            .I(N__9311));
    Odrv12 I__2233 (
            .O(N__9311),
            .I(RAS0n_c));
    InMux I__2232 (
            .O(N__9308),
            .I(N__9305));
    LocalMux I__2231 (
            .O(N__9305),
            .I(N__9302));
    Odrv12 I__2230 (
            .O(N__9302),
            .I(RAS1n_c));
    InMux I__2229 (
            .O(N__9299),
            .I(N__9295));
    InMux I__2228 (
            .O(N__9298),
            .I(N__9292));
    LocalMux I__2227 (
            .O(N__9295),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    LocalMux I__2226 (
            .O(N__9292),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    InMux I__2225 (
            .O(N__9287),
            .I(N__9284));
    LocalMux I__2224 (
            .O(N__9284),
            .I(N__9242));
    ClkMux I__2223 (
            .O(N__9283),
            .I(N__9125));
    ClkMux I__2222 (
            .O(N__9282),
            .I(N__9125));
    ClkMux I__2221 (
            .O(N__9281),
            .I(N__9125));
    ClkMux I__2220 (
            .O(N__9280),
            .I(N__9125));
    ClkMux I__2219 (
            .O(N__9279),
            .I(N__9125));
    ClkMux I__2218 (
            .O(N__9278),
            .I(N__9125));
    ClkMux I__2217 (
            .O(N__9277),
            .I(N__9125));
    ClkMux I__2216 (
            .O(N__9276),
            .I(N__9125));
    ClkMux I__2215 (
            .O(N__9275),
            .I(N__9125));
    ClkMux I__2214 (
            .O(N__9274),
            .I(N__9125));
    ClkMux I__2213 (
            .O(N__9273),
            .I(N__9125));
    ClkMux I__2212 (
            .O(N__9272),
            .I(N__9125));
    ClkMux I__2211 (
            .O(N__9271),
            .I(N__9125));
    ClkMux I__2210 (
            .O(N__9270),
            .I(N__9125));
    ClkMux I__2209 (
            .O(N__9269),
            .I(N__9125));
    ClkMux I__2208 (
            .O(N__9268),
            .I(N__9125));
    ClkMux I__2207 (
            .O(N__9267),
            .I(N__9125));
    ClkMux I__2206 (
            .O(N__9266),
            .I(N__9125));
    ClkMux I__2205 (
            .O(N__9265),
            .I(N__9125));
    ClkMux I__2204 (
            .O(N__9264),
            .I(N__9125));
    ClkMux I__2203 (
            .O(N__9263),
            .I(N__9125));
    ClkMux I__2202 (
            .O(N__9262),
            .I(N__9125));
    ClkMux I__2201 (
            .O(N__9261),
            .I(N__9125));
    ClkMux I__2200 (
            .O(N__9260),
            .I(N__9125));
    ClkMux I__2199 (
            .O(N__9259),
            .I(N__9125));
    ClkMux I__2198 (
            .O(N__9258),
            .I(N__9125));
    ClkMux I__2197 (
            .O(N__9257),
            .I(N__9125));
    ClkMux I__2196 (
            .O(N__9256),
            .I(N__9125));
    ClkMux I__2195 (
            .O(N__9255),
            .I(N__9125));
    ClkMux I__2194 (
            .O(N__9254),
            .I(N__9125));
    ClkMux I__2193 (
            .O(N__9253),
            .I(N__9125));
    ClkMux I__2192 (
            .O(N__9252),
            .I(N__9125));
    ClkMux I__2191 (
            .O(N__9251),
            .I(N__9125));
    ClkMux I__2190 (
            .O(N__9250),
            .I(N__9125));
    ClkMux I__2189 (
            .O(N__9249),
            .I(N__9125));
    ClkMux I__2188 (
            .O(N__9248),
            .I(N__9125));
    ClkMux I__2187 (
            .O(N__9247),
            .I(N__9125));
    ClkMux I__2186 (
            .O(N__9246),
            .I(N__9125));
    ClkMux I__2185 (
            .O(N__9245),
            .I(N__9125));
    Glb2LocalMux I__2184 (
            .O(N__9242),
            .I(N__9125));
    ClkMux I__2183 (
            .O(N__9241),
            .I(N__9125));
    ClkMux I__2182 (
            .O(N__9240),
            .I(N__9125));
    ClkMux I__2181 (
            .O(N__9239),
            .I(N__9125));
    ClkMux I__2180 (
            .O(N__9238),
            .I(N__9125));
    ClkMux I__2179 (
            .O(N__9237),
            .I(N__9125));
    ClkMux I__2178 (
            .O(N__9236),
            .I(N__9125));
    ClkMux I__2177 (
            .O(N__9235),
            .I(N__9125));
    ClkMux I__2176 (
            .O(N__9234),
            .I(N__9125));
    ClkMux I__2175 (
            .O(N__9233),
            .I(N__9125));
    ClkMux I__2174 (
            .O(N__9232),
            .I(N__9125));
    ClkMux I__2173 (
            .O(N__9231),
            .I(N__9125));
    ClkMux I__2172 (
            .O(N__9230),
            .I(N__9125));
    GlobalMux I__2171 (
            .O(N__9125),
            .I(CLK80_OUT));
    CascadeMux I__2170 (
            .O(N__9122),
            .I(N__9113));
    InMux I__2169 (
            .O(N__9121),
            .I(N__9107));
    InMux I__2168 (
            .O(N__9120),
            .I(N__9104));
    InMux I__2167 (
            .O(N__9119),
            .I(N__9101));
    InMux I__2166 (
            .O(N__9118),
            .I(N__9098));
    InMux I__2165 (
            .O(N__9117),
            .I(N__9095));
    InMux I__2164 (
            .O(N__9116),
            .I(N__9092));
    InMux I__2163 (
            .O(N__9113),
            .I(N__9085));
    InMux I__2162 (
            .O(N__9112),
            .I(N__9085));
    InMux I__2161 (
            .O(N__9111),
            .I(N__9085));
    InMux I__2160 (
            .O(N__9110),
            .I(N__9082));
    LocalMux I__2159 (
            .O(N__9107),
            .I(N__9073));
    LocalMux I__2158 (
            .O(N__9104),
            .I(N__9048));
    LocalMux I__2157 (
            .O(N__9101),
            .I(N__9045));
    LocalMux I__2156 (
            .O(N__9098),
            .I(N__9038));
    LocalMux I__2155 (
            .O(N__9095),
            .I(N__9030));
    LocalMux I__2154 (
            .O(N__9092),
            .I(N__9027));
    LocalMux I__2153 (
            .O(N__9085),
            .I(N__9019));
    LocalMux I__2152 (
            .O(N__9082),
            .I(N__9015));
    SRMux I__2151 (
            .O(N__9081),
            .I(N__8903));
    SRMux I__2150 (
            .O(N__9080),
            .I(N__8903));
    SRMux I__2149 (
            .O(N__9079),
            .I(N__8903));
    SRMux I__2148 (
            .O(N__9078),
            .I(N__8903));
    SRMux I__2147 (
            .O(N__9077),
            .I(N__8903));
    SRMux I__2146 (
            .O(N__9076),
            .I(N__8903));
    Glb2LocalMux I__2145 (
            .O(N__9073),
            .I(N__8903));
    SRMux I__2144 (
            .O(N__9072),
            .I(N__8903));
    SRMux I__2143 (
            .O(N__9071),
            .I(N__8903));
    SRMux I__2142 (
            .O(N__9070),
            .I(N__8903));
    SRMux I__2141 (
            .O(N__9069),
            .I(N__8903));
    SRMux I__2140 (
            .O(N__9068),
            .I(N__8903));
    SRMux I__2139 (
            .O(N__9067),
            .I(N__8903));
    SRMux I__2138 (
            .O(N__9066),
            .I(N__8903));
    SRMux I__2137 (
            .O(N__9065),
            .I(N__8903));
    SRMux I__2136 (
            .O(N__9064),
            .I(N__8903));
    SRMux I__2135 (
            .O(N__9063),
            .I(N__8903));
    SRMux I__2134 (
            .O(N__9062),
            .I(N__8903));
    SRMux I__2133 (
            .O(N__9061),
            .I(N__8903));
    SRMux I__2132 (
            .O(N__9060),
            .I(N__8903));
    SRMux I__2131 (
            .O(N__9059),
            .I(N__8903));
    SRMux I__2130 (
            .O(N__9058),
            .I(N__8903));
    SRMux I__2129 (
            .O(N__9057),
            .I(N__8903));
    SRMux I__2128 (
            .O(N__9056),
            .I(N__8903));
    SRMux I__2127 (
            .O(N__9055),
            .I(N__8903));
    SRMux I__2126 (
            .O(N__9054),
            .I(N__8903));
    SRMux I__2125 (
            .O(N__9053),
            .I(N__8903));
    SRMux I__2124 (
            .O(N__9052),
            .I(N__8903));
    SRMux I__2123 (
            .O(N__9051),
            .I(N__8903));
    Glb2LocalMux I__2122 (
            .O(N__9048),
            .I(N__8903));
    Glb2LocalMux I__2121 (
            .O(N__9045),
            .I(N__8903));
    SRMux I__2120 (
            .O(N__9044),
            .I(N__8903));
    SRMux I__2119 (
            .O(N__9043),
            .I(N__8903));
    SRMux I__2118 (
            .O(N__9042),
            .I(N__8903));
    SRMux I__2117 (
            .O(N__9041),
            .I(N__8903));
    Glb2LocalMux I__2116 (
            .O(N__9038),
            .I(N__8903));
    SRMux I__2115 (
            .O(N__9037),
            .I(N__8903));
    SRMux I__2114 (
            .O(N__9036),
            .I(N__8903));
    SRMux I__2113 (
            .O(N__9035),
            .I(N__8903));
    SRMux I__2112 (
            .O(N__9034),
            .I(N__8903));
    SRMux I__2111 (
            .O(N__9033),
            .I(N__8903));
    Glb2LocalMux I__2110 (
            .O(N__9030),
            .I(N__8903));
    Glb2LocalMux I__2109 (
            .O(N__9027),
            .I(N__8903));
    SRMux I__2108 (
            .O(N__9026),
            .I(N__8903));
    SRMux I__2107 (
            .O(N__9025),
            .I(N__8903));
    SRMux I__2106 (
            .O(N__9024),
            .I(N__8903));
    SRMux I__2105 (
            .O(N__9023),
            .I(N__8903));
    SRMux I__2104 (
            .O(N__9022),
            .I(N__8903));
    Glb2LocalMux I__2103 (
            .O(N__9019),
            .I(N__8903));
    SRMux I__2102 (
            .O(N__9018),
            .I(N__8903));
    Glb2LocalMux I__2101 (
            .O(N__9015),
            .I(N__8903));
    SRMux I__2100 (
            .O(N__9014),
            .I(N__8903));
    SRMux I__2099 (
            .O(N__9013),
            .I(N__8903));
    SRMux I__2098 (
            .O(N__9012),
            .I(N__8903));
    GlobalMux I__2097 (
            .O(N__8903),
            .I(N__8900));
    gio2CtrlBuf I__2096 (
            .O(N__8900),
            .I(RESETn_c_i_g));
    IoInMux I__2095 (
            .O(N__8897),
            .I(N__8894));
    LocalMux I__2094 (
            .O(N__8894),
            .I(N__8891));
    Span4Mux_s2_h I__2093 (
            .O(N__8891),
            .I(N__8888));
    Sp12to4 I__2092 (
            .O(N__8888),
            .I(N__8885));
    Span12Mux_s8_v I__2091 (
            .O(N__8885),
            .I(N__8882));
    Odrv12 I__2090 (
            .O(N__8882),
            .I(WEn_c));
    InMux I__2089 (
            .O(N__8879),
            .I(N__8876));
    LocalMux I__2088 (
            .O(N__8876),
            .I(N__8873));
    Span12Mux_v I__2087 (
            .O(N__8873),
            .I(N__8870));
    Span12Mux_h I__2086 (
            .O(N__8870),
            .I(N__8867));
    Odrv12 I__2085 (
            .O(N__8867),
            .I(A_c_17));
    InMux I__2084 (
            .O(N__8864),
            .I(N__8858));
    CascadeMux I__2083 (
            .O(N__8863),
            .I(N__8853));
    InMux I__2082 (
            .O(N__8862),
            .I(N__8845));
    InMux I__2081 (
            .O(N__8861),
            .I(N__8835));
    LocalMux I__2080 (
            .O(N__8858),
            .I(N__8832));
    InMux I__2079 (
            .O(N__8857),
            .I(N__8827));
    InMux I__2078 (
            .O(N__8856),
            .I(N__8827));
    InMux I__2077 (
            .O(N__8853),
            .I(N__8819));
    InMux I__2076 (
            .O(N__8852),
            .I(N__8819));
    InMux I__2075 (
            .O(N__8851),
            .I(N__8819));
    InMux I__2074 (
            .O(N__8850),
            .I(N__8816));
    InMux I__2073 (
            .O(N__8849),
            .I(N__8813));
    InMux I__2072 (
            .O(N__8848),
            .I(N__8810));
    LocalMux I__2071 (
            .O(N__8845),
            .I(N__8807));
    InMux I__2070 (
            .O(N__8844),
            .I(N__8802));
    InMux I__2069 (
            .O(N__8843),
            .I(N__8802));
    InMux I__2068 (
            .O(N__8842),
            .I(N__8797));
    InMux I__2067 (
            .O(N__8841),
            .I(N__8797));
    InMux I__2066 (
            .O(N__8840),
            .I(N__8791));
    InMux I__2065 (
            .O(N__8839),
            .I(N__8788));
    InMux I__2064 (
            .O(N__8838),
            .I(N__8784));
    LocalMux I__2063 (
            .O(N__8835),
            .I(N__8777));
    Span4Mux_v I__2062 (
            .O(N__8832),
            .I(N__8777));
    LocalMux I__2061 (
            .O(N__8827),
            .I(N__8777));
    InMux I__2060 (
            .O(N__8826),
            .I(N__8774));
    LocalMux I__2059 (
            .O(N__8819),
            .I(N__8769));
    LocalMux I__2058 (
            .O(N__8816),
            .I(N__8769));
    LocalMux I__2057 (
            .O(N__8813),
            .I(N__8761));
    LocalMux I__2056 (
            .O(N__8810),
            .I(N__8758));
    Span4Mux_v I__2055 (
            .O(N__8807),
            .I(N__8755));
    LocalMux I__2054 (
            .O(N__8802),
            .I(N__8750));
    LocalMux I__2053 (
            .O(N__8797),
            .I(N__8750));
    InMux I__2052 (
            .O(N__8796),
            .I(N__8745));
    InMux I__2051 (
            .O(N__8795),
            .I(N__8745));
    InMux I__2050 (
            .O(N__8794),
            .I(N__8742));
    LocalMux I__2049 (
            .O(N__8791),
            .I(N__8737));
    LocalMux I__2048 (
            .O(N__8788),
            .I(N__8737));
    InMux I__2047 (
            .O(N__8787),
            .I(N__8734));
    LocalMux I__2046 (
            .O(N__8784),
            .I(N__8727));
    Span4Mux_v I__2045 (
            .O(N__8777),
            .I(N__8727));
    LocalMux I__2044 (
            .O(N__8774),
            .I(N__8727));
    Span4Mux_v I__2043 (
            .O(N__8769),
            .I(N__8724));
    InMux I__2042 (
            .O(N__8768),
            .I(N__8721));
    InMux I__2041 (
            .O(N__8767),
            .I(N__8718));
    InMux I__2040 (
            .O(N__8766),
            .I(N__8711));
    InMux I__2039 (
            .O(N__8765),
            .I(N__8711));
    InMux I__2038 (
            .O(N__8764),
            .I(N__8711));
    Span4Mux_v I__2037 (
            .O(N__8761),
            .I(N__8704));
    Span4Mux_h I__2036 (
            .O(N__8758),
            .I(N__8704));
    Span4Mux_v I__2035 (
            .O(N__8755),
            .I(N__8704));
    Span4Mux_v I__2034 (
            .O(N__8750),
            .I(N__8699));
    LocalMux I__2033 (
            .O(N__8745),
            .I(N__8699));
    LocalMux I__2032 (
            .O(N__8742),
            .I(N__8690));
    Span4Mux_h I__2031 (
            .O(N__8737),
            .I(N__8690));
    LocalMux I__2030 (
            .O(N__8734),
            .I(N__8690));
    Span4Mux_h I__2029 (
            .O(N__8727),
            .I(N__8690));
    Odrv4 I__2028 (
            .O(N__8724),
            .I(CPU_CYCLEm));
    LocalMux I__2027 (
            .O(N__8721),
            .I(CPU_CYCLEm));
    LocalMux I__2026 (
            .O(N__8718),
            .I(CPU_CYCLEm));
    LocalMux I__2025 (
            .O(N__8711),
            .I(CPU_CYCLEm));
    Odrv4 I__2024 (
            .O(N__8704),
            .I(CPU_CYCLEm));
    Odrv4 I__2023 (
            .O(N__8699),
            .I(CPU_CYCLEm));
    Odrv4 I__2022 (
            .O(N__8690),
            .I(CPU_CYCLEm));
    IoInMux I__2021 (
            .O(N__8675),
            .I(N__8672));
    LocalMux I__2020 (
            .O(N__8672),
            .I(N__8669));
    IoSpan4Mux I__2019 (
            .O(N__8669),
            .I(N__8666));
    Span4Mux_s3_h I__2018 (
            .O(N__8666),
            .I(N__8663));
    Span4Mux_h I__2017 (
            .O(N__8663),
            .I(N__8660));
    Span4Mux_h I__2016 (
            .O(N__8660),
            .I(N__8657));
    Odrv4 I__2015 (
            .O(N__8657),
            .I(CMA_c_8));
    CEMux I__2014 (
            .O(N__8654),
            .I(N__8650));
    CEMux I__2013 (
            .O(N__8653),
            .I(N__8647));
    LocalMux I__2012 (
            .O(N__8650),
            .I(N__8640));
    LocalMux I__2011 (
            .O(N__8647),
            .I(N__8640));
    CEMux I__2010 (
            .O(N__8646),
            .I(N__8637));
    CEMux I__2009 (
            .O(N__8645),
            .I(N__8634));
    Span4Mux_h I__2008 (
            .O(N__8640),
            .I(N__8628));
    LocalMux I__2007 (
            .O(N__8637),
            .I(N__8628));
    LocalMux I__2006 (
            .O(N__8634),
            .I(N__8625));
    CEMux I__2005 (
            .O(N__8633),
            .I(N__8622));
    Span4Mux_h I__2004 (
            .O(N__8628),
            .I(N__8618));
    Span4Mux_v I__2003 (
            .O(N__8625),
            .I(N__8613));
    LocalMux I__2002 (
            .O(N__8622),
            .I(N__8610));
    CEMux I__2001 (
            .O(N__8621),
            .I(N__8607));
    Span4Mux_h I__2000 (
            .O(N__8618),
            .I(N__8604));
    CEMux I__1999 (
            .O(N__8617),
            .I(N__8601));
    CEMux I__1998 (
            .O(N__8616),
            .I(N__8598));
    Odrv4 I__1997 (
            .O(N__8613),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    Odrv12 I__1996 (
            .O(N__8610),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    LocalMux I__1995 (
            .O(N__8607),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    Odrv4 I__1994 (
            .O(N__8604),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    LocalMux I__1993 (
            .O(N__8601),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    LocalMux I__1992 (
            .O(N__8598),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    InMux I__1991 (
            .O(N__8585),
            .I(N__8578));
    InMux I__1990 (
            .O(N__8584),
            .I(N__8569));
    InMux I__1989 (
            .O(N__8583),
            .I(N__8569));
    InMux I__1988 (
            .O(N__8582),
            .I(N__8564));
    InMux I__1987 (
            .O(N__8581),
            .I(N__8564));
    LocalMux I__1986 (
            .O(N__8578),
            .I(N__8561));
    InMux I__1985 (
            .O(N__8577),
            .I(N__8558));
    InMux I__1984 (
            .O(N__8576),
            .I(N__8553));
    InMux I__1983 (
            .O(N__8575),
            .I(N__8549));
    InMux I__1982 (
            .O(N__8574),
            .I(N__8546));
    LocalMux I__1981 (
            .O(N__8569),
            .I(N__8543));
    LocalMux I__1980 (
            .O(N__8564),
            .I(N__8538));
    Span4Mux_h I__1979 (
            .O(N__8561),
            .I(N__8538));
    LocalMux I__1978 (
            .O(N__8558),
            .I(N__8535));
    CascadeMux I__1977 (
            .O(N__8557),
            .I(N__8532));
    InMux I__1976 (
            .O(N__8556),
            .I(N__8529));
    LocalMux I__1975 (
            .O(N__8553),
            .I(N__8526));
    InMux I__1974 (
            .O(N__8552),
            .I(N__8523));
    LocalMux I__1973 (
            .O(N__8549),
            .I(N__8518));
    LocalMux I__1972 (
            .O(N__8546),
            .I(N__8518));
    Span4Mux_v I__1971 (
            .O(N__8543),
            .I(N__8511));
    Span4Mux_v I__1970 (
            .O(N__8538),
            .I(N__8511));
    Span4Mux_h I__1969 (
            .O(N__8535),
            .I(N__8511));
    InMux I__1968 (
            .O(N__8532),
            .I(N__8506));
    LocalMux I__1967 (
            .O(N__8529),
            .I(N__8503));
    Span4Mux_v I__1966 (
            .O(N__8526),
            .I(N__8500));
    LocalMux I__1965 (
            .O(N__8523),
            .I(N__8495));
    Span4Mux_h I__1964 (
            .O(N__8518),
            .I(N__8495));
    Span4Mux_h I__1963 (
            .O(N__8511),
            .I(N__8492));
    InMux I__1962 (
            .O(N__8510),
            .I(N__8487));
    InMux I__1961 (
            .O(N__8509),
            .I(N__8487));
    LocalMux I__1960 (
            .O(N__8506),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    Odrv12 I__1959 (
            .O(N__8503),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    Odrv4 I__1958 (
            .O(N__8500),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    Odrv4 I__1957 (
            .O(N__8495),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    Odrv4 I__1956 (
            .O(N__8492),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    LocalMux I__1955 (
            .O(N__8487),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    CascadeMux I__1954 (
            .O(N__8474),
            .I(N__8467));
    CascadeMux I__1953 (
            .O(N__8473),
            .I(N__8464));
    CascadeMux I__1952 (
            .O(N__8472),
            .I(N__8458));
    CascadeMux I__1951 (
            .O(N__8471),
            .I(N__8455));
    InMux I__1950 (
            .O(N__8470),
            .I(N__8451));
    InMux I__1949 (
            .O(N__8467),
            .I(N__8446));
    InMux I__1948 (
            .O(N__8464),
            .I(N__8446));
    InMux I__1947 (
            .O(N__8463),
            .I(N__8443));
    InMux I__1946 (
            .O(N__8462),
            .I(N__8437));
    InMux I__1945 (
            .O(N__8461),
            .I(N__8437));
    InMux I__1944 (
            .O(N__8458),
            .I(N__8434));
    InMux I__1943 (
            .O(N__8455),
            .I(N__8430));
    InMux I__1942 (
            .O(N__8454),
            .I(N__8427));
    LocalMux I__1941 (
            .O(N__8451),
            .I(N__8424));
    LocalMux I__1940 (
            .O(N__8446),
            .I(N__8421));
    LocalMux I__1939 (
            .O(N__8443),
            .I(N__8418));
    InMux I__1938 (
            .O(N__8442),
            .I(N__8413));
    LocalMux I__1937 (
            .O(N__8437),
            .I(N__8410));
    LocalMux I__1936 (
            .O(N__8434),
            .I(N__8407));
    InMux I__1935 (
            .O(N__8433),
            .I(N__8404));
    LocalMux I__1934 (
            .O(N__8430),
            .I(N__8401));
    LocalMux I__1933 (
            .O(N__8427),
            .I(N__8398));
    Span4Mux_v I__1932 (
            .O(N__8424),
            .I(N__8395));
    Span4Mux_v I__1931 (
            .O(N__8421),
            .I(N__8390));
    Span4Mux_h I__1930 (
            .O(N__8418),
            .I(N__8390));
    CascadeMux I__1929 (
            .O(N__8417),
            .I(N__8386));
    InMux I__1928 (
            .O(N__8416),
            .I(N__8383));
    LocalMux I__1927 (
            .O(N__8413),
            .I(N__8380));
    Span4Mux_h I__1926 (
            .O(N__8410),
            .I(N__8375));
    Span4Mux_h I__1925 (
            .O(N__8407),
            .I(N__8375));
    LocalMux I__1924 (
            .O(N__8404),
            .I(N__8370));
    Span4Mux_h I__1923 (
            .O(N__8401),
            .I(N__8370));
    Span4Mux_v I__1922 (
            .O(N__8398),
            .I(N__8365));
    Span4Mux_h I__1921 (
            .O(N__8395),
            .I(N__8365));
    Span4Mux_h I__1920 (
            .O(N__8390),
            .I(N__8362));
    InMux I__1919 (
            .O(N__8389),
            .I(N__8357));
    InMux I__1918 (
            .O(N__8386),
            .I(N__8357));
    LocalMux I__1917 (
            .O(N__8383),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv12 I__1916 (
            .O(N__8380),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1915 (
            .O(N__8375),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1914 (
            .O(N__8370),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1913 (
            .O(N__8365),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1912 (
            .O(N__8362),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1911 (
            .O(N__8357),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    InMux I__1910 (
            .O(N__8342),
            .I(N__8338));
    InMux I__1909 (
            .O(N__8341),
            .I(N__8335));
    LocalMux I__1908 (
            .O(N__8338),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    LocalMux I__1907 (
            .O(N__8335),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    InMux I__1906 (
            .O(N__8330),
            .I(N__8327));
    LocalMux I__1905 (
            .O(N__8327),
            .I(N__8324));
    Span4Mux_v I__1904 (
            .O(N__8324),
            .I(N__8320));
    InMux I__1903 (
            .O(N__8323),
            .I(N__8317));
    Sp12to4 I__1902 (
            .O(N__8320),
            .I(N__8314));
    LocalMux I__1901 (
            .O(N__8317),
            .I(N__8311));
    Span12Mux_h I__1900 (
            .O(N__8314),
            .I(N__8308));
    Span12Mux_v I__1899 (
            .O(N__8311),
            .I(N__8305));
    Span12Mux_v I__1898 (
            .O(N__8308),
            .I(N__8302));
    Span12Mux_h I__1897 (
            .O(N__8305),
            .I(N__8299));
    Odrv12 I__1896 (
            .O(N__8302),
            .I(DRA_c_4));
    Odrv12 I__1895 (
            .O(N__8299),
            .I(DRA_c_4));
    InMux I__1894 (
            .O(N__8294),
            .I(N__8291));
    LocalMux I__1893 (
            .O(N__8291),
            .I(N__8288));
    Odrv4 I__1892 (
            .O(N__8288),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    CEMux I__1891 (
            .O(N__8285),
            .I(N__8282));
    LocalMux I__1890 (
            .O(N__8282),
            .I(N__8276));
    CEMux I__1889 (
            .O(N__8281),
            .I(N__8273));
    CEMux I__1888 (
            .O(N__8280),
            .I(N__8270));
    CEMux I__1887 (
            .O(N__8279),
            .I(N__8267));
    Span4Mux_h I__1886 (
            .O(N__8276),
            .I(N__8263));
    LocalMux I__1885 (
            .O(N__8273),
            .I(N__8258));
    LocalMux I__1884 (
            .O(N__8270),
            .I(N__8258));
    LocalMux I__1883 (
            .O(N__8267),
            .I(N__8255));
    CEMux I__1882 (
            .O(N__8266),
            .I(N__8252));
    Span4Mux_h I__1881 (
            .O(N__8263),
            .I(N__8247));
    Span4Mux_h I__1880 (
            .O(N__8258),
            .I(N__8244));
    Span4Mux_v I__1879 (
            .O(N__8255),
            .I(N__8241));
    LocalMux I__1878 (
            .O(N__8252),
            .I(N__8238));
    CEMux I__1877 (
            .O(N__8251),
            .I(N__8235));
    CEMux I__1876 (
            .O(N__8250),
            .I(N__8232));
    Odrv4 I__1875 (
            .O(N__8247),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    Odrv4 I__1874 (
            .O(N__8244),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    Odrv4 I__1873 (
            .O(N__8241),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    Odrv12 I__1872 (
            .O(N__8238),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    LocalMux I__1871 (
            .O(N__8235),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    LocalMux I__1870 (
            .O(N__8232),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    IoInMux I__1869 (
            .O(N__8219),
            .I(N__8216));
    LocalMux I__1868 (
            .O(N__8216),
            .I(N__8212));
    IoInMux I__1867 (
            .O(N__8215),
            .I(N__8209));
    IoSpan4Mux I__1866 (
            .O(N__8212),
            .I(N__8206));
    LocalMux I__1865 (
            .O(N__8209),
            .I(N__8203));
    IoSpan4Mux I__1864 (
            .O(N__8206),
            .I(N__8200));
    Span4Mux_s2_v I__1863 (
            .O(N__8203),
            .I(N__8197));
    Span4Mux_s3_h I__1862 (
            .O(N__8200),
            .I(N__8194));
    Span4Mux_v I__1861 (
            .O(N__8197),
            .I(N__8191));
    Span4Mux_h I__1860 (
            .O(N__8194),
            .I(N__8188));
    Span4Mux_v I__1859 (
            .O(N__8191),
            .I(N__8185));
    Odrv4 I__1858 (
            .O(N__8188),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1857 (
            .O(N__8185),
            .I(CONSTANT_ONE_NET));
    InMux I__1856 (
            .O(N__8180),
            .I(N__8177));
    LocalMux I__1855 (
            .O(N__8177),
            .I(N__8173));
    InMux I__1854 (
            .O(N__8176),
            .I(N__8170));
    Span4Mux_v I__1853 (
            .O(N__8173),
            .I(N__8167));
    LocalMux I__1852 (
            .O(N__8170),
            .I(N__8164));
    Sp12to4 I__1851 (
            .O(N__8167),
            .I(N__8161));
    Span4Mux_v I__1850 (
            .O(N__8164),
            .I(N__8158));
    Span12Mux_h I__1849 (
            .O(N__8161),
            .I(N__8155));
    Sp12to4 I__1848 (
            .O(N__8158),
            .I(N__8152));
    Odrv12 I__1847 (
            .O(N__8155),
            .I(DRA_c_8));
    Odrv12 I__1846 (
            .O(N__8152),
            .I(DRA_c_8));
    CascadeMux I__1845 (
            .O(N__8147),
            .I(N__8144));
    InMux I__1844 (
            .O(N__8144),
            .I(N__8141));
    LocalMux I__1843 (
            .O(N__8141),
            .I(N__8138));
    Odrv4 I__1842 (
            .O(N__8138),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__1841 (
            .O(N__8135),
            .I(N__8130));
    CascadeMux I__1840 (
            .O(N__8134),
            .I(N__8126));
    CascadeMux I__1839 (
            .O(N__8133),
            .I(N__8120));
    LocalMux I__1838 (
            .O(N__8130),
            .I(N__8111));
    InMux I__1837 (
            .O(N__8129),
            .I(N__8108));
    InMux I__1836 (
            .O(N__8126),
            .I(N__8105));
    CascadeMux I__1835 (
            .O(N__8125),
            .I(N__8102));
    CascadeMux I__1834 (
            .O(N__8124),
            .I(N__8099));
    InMux I__1833 (
            .O(N__8123),
            .I(N__8096));
    InMux I__1832 (
            .O(N__8120),
            .I(N__8093));
    InMux I__1831 (
            .O(N__8119),
            .I(N__8090));
    CascadeMux I__1830 (
            .O(N__8118),
            .I(N__8087));
    InMux I__1829 (
            .O(N__8117),
            .I(N__8084));
    CascadeMux I__1828 (
            .O(N__8116),
            .I(N__8081));
    CascadeMux I__1827 (
            .O(N__8115),
            .I(N__8078));
    CascadeMux I__1826 (
            .O(N__8114),
            .I(N__8075));
    Span4Mux_v I__1825 (
            .O(N__8111),
            .I(N__8072));
    LocalMux I__1824 (
            .O(N__8108),
            .I(N__8067));
    LocalMux I__1823 (
            .O(N__8105),
            .I(N__8067));
    InMux I__1822 (
            .O(N__8102),
            .I(N__8062));
    InMux I__1821 (
            .O(N__8099),
            .I(N__8062));
    LocalMux I__1820 (
            .O(N__8096),
            .I(N__8057));
    LocalMux I__1819 (
            .O(N__8093),
            .I(N__8054));
    LocalMux I__1818 (
            .O(N__8090),
            .I(N__8051));
    InMux I__1817 (
            .O(N__8087),
            .I(N__8048));
    LocalMux I__1816 (
            .O(N__8084),
            .I(N__8045));
    InMux I__1815 (
            .O(N__8081),
            .I(N__8042));
    InMux I__1814 (
            .O(N__8078),
            .I(N__8039));
    InMux I__1813 (
            .O(N__8075),
            .I(N__8036));
    Span4Mux_h I__1812 (
            .O(N__8072),
            .I(N__8029));
    Span4Mux_v I__1811 (
            .O(N__8067),
            .I(N__8029));
    LocalMux I__1810 (
            .O(N__8062),
            .I(N__8029));
    CascadeMux I__1809 (
            .O(N__8061),
            .I(N__8026));
    InMux I__1808 (
            .O(N__8060),
            .I(N__8022));
    Span4Mux_v I__1807 (
            .O(N__8057),
            .I(N__8017));
    Span4Mux_v I__1806 (
            .O(N__8054),
            .I(N__8017));
    Span4Mux_h I__1805 (
            .O(N__8051),
            .I(N__8012));
    LocalMux I__1804 (
            .O(N__8048),
            .I(N__8012));
    Span12Mux_v I__1803 (
            .O(N__8045),
            .I(N__8005));
    LocalMux I__1802 (
            .O(N__8042),
            .I(N__8005));
    LocalMux I__1801 (
            .O(N__8039),
            .I(N__8005));
    LocalMux I__1800 (
            .O(N__8036),
            .I(N__8002));
    Span4Mux_h I__1799 (
            .O(N__8029),
            .I(N__7999));
    InMux I__1798 (
            .O(N__8026),
            .I(N__7994));
    InMux I__1797 (
            .O(N__8025),
            .I(N__7994));
    LocalMux I__1796 (
            .O(N__8022),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1795 (
            .O(N__8017),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1794 (
            .O(N__8012),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv12 I__1793 (
            .O(N__8005),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1792 (
            .O(N__8002),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1791 (
            .O(N__7999),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1790 (
            .O(N__7994),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    IoInMux I__1789 (
            .O(N__7979),
            .I(N__7976));
    LocalMux I__1788 (
            .O(N__7976),
            .I(N__7973));
    IoSpan4Mux I__1787 (
            .O(N__7973),
            .I(N__7970));
    Sp12to4 I__1786 (
            .O(N__7970),
            .I(N__7967));
    Span12Mux_s9_v I__1785 (
            .O(N__7967),
            .I(N__7964));
    Odrv12 I__1784 (
            .O(N__7964),
            .I(CASn_c));
    CEMux I__1783 (
            .O(N__7961),
            .I(N__7958));
    LocalMux I__1782 (
            .O(N__7958),
            .I(N__7953));
    CEMux I__1781 (
            .O(N__7957),
            .I(N__7950));
    CEMux I__1780 (
            .O(N__7956),
            .I(N__7947));
    Span4Mux_v I__1779 (
            .O(N__7953),
            .I(N__7942));
    LocalMux I__1778 (
            .O(N__7950),
            .I(N__7942));
    LocalMux I__1777 (
            .O(N__7947),
            .I(N__7938));
    Span4Mux_h I__1776 (
            .O(N__7942),
            .I(N__7935));
    CEMux I__1775 (
            .O(N__7941),
            .I(N__7932));
    Span4Mux_h I__1774 (
            .O(N__7938),
            .I(N__7928));
    Span4Mux_h I__1773 (
            .O(N__7935),
            .I(N__7925));
    LocalMux I__1772 (
            .O(N__7932),
            .I(N__7922));
    CEMux I__1771 (
            .O(N__7931),
            .I(N__7919));
    Odrv4 I__1770 (
            .O(N__7928),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    Odrv4 I__1769 (
            .O(N__7925),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    Odrv4 I__1768 (
            .O(N__7922),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    LocalMux I__1767 (
            .O(N__7919),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    InMux I__1766 (
            .O(N__7910),
            .I(N__7907));
    LocalMux I__1765 (
            .O(N__7907),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ));
    InMux I__1764 (
            .O(N__7904),
            .I(N__7901));
    LocalMux I__1763 (
            .O(N__7901),
            .I(N__7897));
    InMux I__1762 (
            .O(N__7900),
            .I(N__7894));
    Span4Mux_h I__1761 (
            .O(N__7897),
            .I(N__7889));
    LocalMux I__1760 (
            .O(N__7894),
            .I(N__7889));
    Span4Mux_h I__1759 (
            .O(N__7889),
            .I(N__7886));
    Sp12to4 I__1758 (
            .O(N__7886),
            .I(N__7883));
    Span12Mux_v I__1757 (
            .O(N__7883),
            .I(N__7880));
    Odrv12 I__1756 (
            .O(N__7880),
            .I(DRA_c_6));
    InMux I__1755 (
            .O(N__7877),
            .I(N__7874));
    LocalMux I__1754 (
            .O(N__7874),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__1753 (
            .O(N__7871),
            .I(N__7868));
    LocalMux I__1752 (
            .O(N__7868),
            .I(N__7865));
    Span4Mux_v I__1751 (
            .O(N__7865),
            .I(N__7861));
    InMux I__1750 (
            .O(N__7864),
            .I(N__7858));
    Span4Mux_h I__1749 (
            .O(N__7861),
            .I(N__7853));
    LocalMux I__1748 (
            .O(N__7858),
            .I(N__7853));
    Span4Mux_h I__1747 (
            .O(N__7853),
            .I(N__7850));
    Sp12to4 I__1746 (
            .O(N__7850),
            .I(N__7847));
    Span12Mux_v I__1745 (
            .O(N__7847),
            .I(N__7844));
    Odrv12 I__1744 (
            .O(N__7844),
            .I(DRA_c_5));
    InMux I__1743 (
            .O(N__7841),
            .I(N__7838));
    LocalMux I__1742 (
            .O(N__7838),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__1741 (
            .O(N__7835),
            .I(N__7832));
    LocalMux I__1740 (
            .O(N__7832),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__1739 (
            .O(N__7829),
            .I(N__7826));
    LocalMux I__1738 (
            .O(N__7826),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__1737 (
            .O(N__7823),
            .I(N__7820));
    LocalMux I__1736 (
            .O(N__7820),
            .I(N__7817));
    Span4Mux_v I__1735 (
            .O(N__7817),
            .I(N__7813));
    InMux I__1734 (
            .O(N__7816),
            .I(N__7810));
    Sp12to4 I__1733 (
            .O(N__7813),
            .I(N__7805));
    LocalMux I__1732 (
            .O(N__7810),
            .I(N__7805));
    Span12Mux_h I__1731 (
            .O(N__7805),
            .I(N__7802));
    Span12Mux_v I__1730 (
            .O(N__7802),
            .I(N__7799));
    Odrv12 I__1729 (
            .O(N__7799),
            .I(DRA_c_1));
    InMux I__1728 (
            .O(N__7796),
            .I(N__7793));
    LocalMux I__1727 (
            .O(N__7793),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__1726 (
            .O(N__7790),
            .I(N__7786));
    InMux I__1725 (
            .O(N__7789),
            .I(N__7783));
    LocalMux I__1724 (
            .O(N__7786),
            .I(N__7780));
    LocalMux I__1723 (
            .O(N__7783),
            .I(N__7777));
    Span4Mux_h I__1722 (
            .O(N__7780),
            .I(N__7774));
    Span12Mux_v I__1721 (
            .O(N__7777),
            .I(N__7771));
    Sp12to4 I__1720 (
            .O(N__7774),
            .I(N__7768));
    Span12Mux_h I__1719 (
            .O(N__7771),
            .I(N__7765));
    Span12Mux_v I__1718 (
            .O(N__7768),
            .I(N__7762));
    Odrv12 I__1717 (
            .O(N__7765),
            .I(DRA_c_2));
    Odrv12 I__1716 (
            .O(N__7762),
            .I(DRA_c_2));
    InMux I__1715 (
            .O(N__7757),
            .I(N__7754));
    LocalMux I__1714 (
            .O(N__7754),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__1713 (
            .O(N__7751),
            .I(N__7746));
    InMux I__1712 (
            .O(N__7750),
            .I(N__7743));
    InMux I__1711 (
            .O(N__7749),
            .I(N__7740));
    LocalMux I__1710 (
            .O(N__7746),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    LocalMux I__1709 (
            .O(N__7743),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    LocalMux I__1708 (
            .O(N__7740),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__1707 (
            .O(N__7733),
            .I(N__7729));
    InMux I__1706 (
            .O(N__7732),
            .I(N__7726));
    LocalMux I__1705 (
            .O(N__7729),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    LocalMux I__1704 (
            .O(N__7726),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__1703 (
            .O(N__7721),
            .I(N__7718));
    LocalMux I__1702 (
            .O(N__7718),
            .I(N__7714));
    InMux I__1701 (
            .O(N__7717),
            .I(N__7711));
    Span4Mux_v I__1700 (
            .O(N__7714),
            .I(N__7706));
    LocalMux I__1699 (
            .O(N__7711),
            .I(N__7706));
    Sp12to4 I__1698 (
            .O(N__7706),
            .I(N__7703));
    Span12Mux_v I__1697 (
            .O(N__7703),
            .I(N__7700));
    Span12Mux_h I__1696 (
            .O(N__7700),
            .I(N__7697));
    Odrv12 I__1695 (
            .O(N__7697),
            .I(DRA_c_0));
    CascadeMux I__1694 (
            .O(N__7694),
            .I(N__7691));
    InMux I__1693 (
            .O(N__7691),
            .I(N__7688));
    LocalMux I__1692 (
            .O(N__7688),
            .I(N__7685));
    Span4Mux_h I__1691 (
            .O(N__7685),
            .I(N__7682));
    Odrv4 I__1690 (
            .O(N__7682),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    IoInMux I__1689 (
            .O(N__7679),
            .I(N__7676));
    LocalMux I__1688 (
            .O(N__7676),
            .I(N__7673));
    Span4Mux_s3_v I__1687 (
            .O(N__7673),
            .I(N__7670));
    Span4Mux_v I__1686 (
            .O(N__7670),
            .I(N__7667));
    Sp12to4 I__1685 (
            .O(N__7667),
            .I(N__7664));
    Odrv12 I__1684 (
            .O(N__7664),
            .I(RASn_c));
    InMux I__1683 (
            .O(N__7661),
            .I(N__7658));
    LocalMux I__1682 (
            .O(N__7658),
            .I(N__7655));
    Span4Mux_v I__1681 (
            .O(N__7655),
            .I(N__7652));
    Odrv4 I__1680 (
            .O(N__7652),
            .I(\U712_BYTE_ENABLE.un2_CLMBEnZ0 ));
    IoInMux I__1679 (
            .O(N__7649),
            .I(N__7646));
    LocalMux I__1678 (
            .O(N__7646),
            .I(N__7643));
    Span4Mux_s3_h I__1677 (
            .O(N__7643),
            .I(N__7640));
    Span4Mux_v I__1676 (
            .O(N__7640),
            .I(N__7637));
    Sp12to4 I__1675 (
            .O(N__7637),
            .I(N__7634));
    Span12Mux_v I__1674 (
            .O(N__7634),
            .I(N__7631));
    Odrv12 I__1673 (
            .O(N__7631),
            .I(CLMBEn_c));
    InMux I__1672 (
            .O(N__7628),
            .I(N__7623));
    InMux I__1671 (
            .O(N__7627),
            .I(N__7618));
    InMux I__1670 (
            .O(N__7626),
            .I(N__7618));
    LocalMux I__1669 (
            .O(N__7623),
            .I(N__7613));
    LocalMux I__1668 (
            .O(N__7618),
            .I(N__7613));
    Span4Mux_v I__1667 (
            .O(N__7613),
            .I(N__7610));
    Sp12to4 I__1666 (
            .O(N__7610),
            .I(N__7607));
    Span12Mux_h I__1665 (
            .O(N__7607),
            .I(N__7604));
    Span12Mux_v I__1664 (
            .O(N__7604),
            .I(N__7601));
    Odrv12 I__1663 (
            .O(N__7601),
            .I(CASUn_c));
    IoInMux I__1662 (
            .O(N__7598),
            .I(N__7593));
    CascadeMux I__1661 (
            .O(N__7597),
            .I(N__7589));
    CascadeMux I__1660 (
            .O(N__7596),
            .I(N__7586));
    LocalMux I__1659 (
            .O(N__7593),
            .I(N__7583));
    InMux I__1658 (
            .O(N__7592),
            .I(N__7580));
    InMux I__1657 (
            .O(N__7589),
            .I(N__7575));
    InMux I__1656 (
            .O(N__7586),
            .I(N__7575));
    Span12Mux_s5_v I__1655 (
            .O(N__7583),
            .I(N__7572));
    LocalMux I__1654 (
            .O(N__7580),
            .I(N__7567));
    LocalMux I__1653 (
            .O(N__7575),
            .I(N__7567));
    Span12Mux_v I__1652 (
            .O(N__7572),
            .I(N__7562));
    Span4Mux_v I__1651 (
            .O(N__7567),
            .I(N__7559));
    InMux I__1650 (
            .O(N__7566),
            .I(N__7556));
    InMux I__1649 (
            .O(N__7565),
            .I(N__7553));
    Odrv12 I__1648 (
            .O(N__7562),
            .I(DBENn_c));
    Odrv4 I__1647 (
            .O(N__7559),
            .I(DBENn_c));
    LocalMux I__1646 (
            .O(N__7556),
            .I(DBENn_c));
    LocalMux I__1645 (
            .O(N__7553),
            .I(DBENn_c));
    InMux I__1644 (
            .O(N__7544),
            .I(N__7541));
    LocalMux I__1643 (
            .O(N__7541),
            .I(N__7538));
    Span4Mux_v I__1642 (
            .O(N__7538),
            .I(N__7535));
    Odrv4 I__1641 (
            .O(N__7535),
            .I(\U712_BYTE_ENABLE.un2_CUUBEnZ0 ));
    IoInMux I__1640 (
            .O(N__7532),
            .I(N__7529));
    LocalMux I__1639 (
            .O(N__7529),
            .I(N__7526));
    IoSpan4Mux I__1638 (
            .O(N__7526),
            .I(N__7523));
    IoSpan4Mux I__1637 (
            .O(N__7523),
            .I(N__7520));
    Span4Mux_s3_h I__1636 (
            .O(N__7520),
            .I(N__7517));
    Sp12to4 I__1635 (
            .O(N__7517),
            .I(N__7514));
    Odrv12 I__1634 (
            .O(N__7514),
            .I(CUUBEn_c));
    CascadeMux I__1633 (
            .O(N__7511),
            .I(N__7508));
    InMux I__1632 (
            .O(N__7508),
            .I(N__7504));
    InMux I__1631 (
            .O(N__7507),
            .I(N__7501));
    LocalMux I__1630 (
            .O(N__7504),
            .I(N__7497));
    LocalMux I__1629 (
            .O(N__7501),
            .I(N__7494));
    InMux I__1628 (
            .O(N__7500),
            .I(N__7491));
    Span4Mux_v I__1627 (
            .O(N__7497),
            .I(N__7487));
    Span12Mux_h I__1626 (
            .O(N__7494),
            .I(N__7482));
    LocalMux I__1625 (
            .O(N__7491),
            .I(N__7482));
    InMux I__1624 (
            .O(N__7490),
            .I(N__7479));
    Odrv4 I__1623 (
            .O(N__7487),
            .I(REG_CYCLEm));
    Odrv12 I__1622 (
            .O(N__7482),
            .I(REG_CYCLEm));
    LocalMux I__1621 (
            .O(N__7479),
            .I(REG_CYCLEm));
    InMux I__1620 (
            .O(N__7472),
            .I(N__7466));
    CascadeMux I__1619 (
            .O(N__7471),
            .I(N__7462));
    InMux I__1618 (
            .O(N__7470),
            .I(N__7457));
    InMux I__1617 (
            .O(N__7469),
            .I(N__7454));
    LocalMux I__1616 (
            .O(N__7466),
            .I(N__7451));
    InMux I__1615 (
            .O(N__7465),
            .I(N__7444));
    InMux I__1614 (
            .O(N__7462),
            .I(N__7444));
    InMux I__1613 (
            .O(N__7461),
            .I(N__7444));
    CascadeMux I__1612 (
            .O(N__7460),
            .I(N__7441));
    LocalMux I__1611 (
            .O(N__7457),
            .I(N__7434));
    LocalMux I__1610 (
            .O(N__7454),
            .I(N__7434));
    Span4Mux_v I__1609 (
            .O(N__7451),
            .I(N__7429));
    LocalMux I__1608 (
            .O(N__7444),
            .I(N__7429));
    InMux I__1607 (
            .O(N__7441),
            .I(N__7426));
    InMux I__1606 (
            .O(N__7440),
            .I(N__7423));
    InMux I__1605 (
            .O(N__7439),
            .I(N__7420));
    Span4Mux_h I__1604 (
            .O(N__7434),
            .I(N__7417));
    Odrv4 I__1603 (
            .O(N__7429),
            .I(DMA_CYCLEm));
    LocalMux I__1602 (
            .O(N__7426),
            .I(DMA_CYCLEm));
    LocalMux I__1601 (
            .O(N__7423),
            .I(DMA_CYCLEm));
    LocalMux I__1600 (
            .O(N__7420),
            .I(DMA_CYCLEm));
    Odrv4 I__1599 (
            .O(N__7417),
            .I(DMA_CYCLEm));
    IoInMux I__1598 (
            .O(N__7406),
            .I(N__7403));
    LocalMux I__1597 (
            .O(N__7403),
            .I(N__7400));
    Span4Mux_s2_v I__1596 (
            .O(N__7400),
            .I(N__7397));
    Sp12to4 I__1595 (
            .O(N__7397),
            .I(N__7394));
    Span12Mux_s7_h I__1594 (
            .O(N__7394),
            .I(N__7391));
    Span12Mux_v I__1593 (
            .O(N__7391),
            .I(N__7388));
    Odrv12 I__1592 (
            .O(N__7388),
            .I(N_52_i));
    InMux I__1591 (
            .O(N__7385),
            .I(N__7381));
    InMux I__1590 (
            .O(N__7384),
            .I(N__7378));
    LocalMux I__1589 (
            .O(N__7381),
            .I(N__7375));
    LocalMux I__1588 (
            .O(N__7378),
            .I(N__7372));
    Span4Mux_h I__1587 (
            .O(N__7375),
            .I(N__7369));
    Sp12to4 I__1586 (
            .O(N__7372),
            .I(N__7366));
    Span4Mux_v I__1585 (
            .O(N__7369),
            .I(N__7363));
    Span12Mux_v I__1584 (
            .O(N__7366),
            .I(N__7358));
    Sp12to4 I__1583 (
            .O(N__7363),
            .I(N__7358));
    Span12Mux_h I__1582 (
            .O(N__7358),
            .I(N__7355));
    Odrv12 I__1581 (
            .O(N__7355),
            .I(DRA_c_7));
    InMux I__1580 (
            .O(N__7352),
            .I(N__7349));
    LocalMux I__1579 (
            .O(N__7349),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__1578 (
            .O(N__7346),
            .I(N__7343));
    LocalMux I__1577 (
            .O(N__7343),
            .I(\U712_CHIP_RAM.N_37 ));
    IoInMux I__1576 (
            .O(N__7340),
            .I(N__7337));
    LocalMux I__1575 (
            .O(N__7337),
            .I(N__7334));
    Span4Mux_s3_h I__1574 (
            .O(N__7334),
            .I(N__7331));
    Span4Mux_v I__1573 (
            .O(N__7331),
            .I(N__7328));
    Sp12to4 I__1572 (
            .O(N__7328),
            .I(N__7325));
    Span12Mux_h I__1571 (
            .O(N__7325),
            .I(N__7322));
    Odrv12 I__1570 (
            .O(N__7322),
            .I(CMA_c_5));
    InMux I__1569 (
            .O(N__7319),
            .I(N__7316));
    LocalMux I__1568 (
            .O(N__7316),
            .I(\U712_CHIP_RAM.N_39 ));
    IoInMux I__1567 (
            .O(N__7313),
            .I(N__7310));
    LocalMux I__1566 (
            .O(N__7310),
            .I(N__7307));
    IoSpan4Mux I__1565 (
            .O(N__7307),
            .I(N__7304));
    Span4Mux_s2_h I__1564 (
            .O(N__7304),
            .I(N__7301));
    Span4Mux_v I__1563 (
            .O(N__7301),
            .I(N__7298));
    Sp12to4 I__1562 (
            .O(N__7298),
            .I(N__7295));
    Odrv12 I__1561 (
            .O(N__7295),
            .I(CMA_c_7));
    InMux I__1560 (
            .O(N__7292),
            .I(N__7289));
    LocalMux I__1559 (
            .O(N__7289),
            .I(N__7286));
    Span4Mux_v I__1558 (
            .O(N__7286),
            .I(N__7283));
    Span4Mux_v I__1557 (
            .O(N__7283),
            .I(N__7280));
    Sp12to4 I__1556 (
            .O(N__7280),
            .I(N__7277));
    Span12Mux_h I__1555 (
            .O(N__7277),
            .I(N__7274));
    Odrv12 I__1554 (
            .O(N__7274),
            .I(A_c_19));
    IoInMux I__1553 (
            .O(N__7271),
            .I(N__7268));
    LocalMux I__1552 (
            .O(N__7268),
            .I(N__7265));
    IoSpan4Mux I__1551 (
            .O(N__7265),
            .I(N__7262));
    IoSpan4Mux I__1550 (
            .O(N__7262),
            .I(N__7259));
    Span4Mux_s2_h I__1549 (
            .O(N__7259),
            .I(N__7256));
    Sp12to4 I__1548 (
            .O(N__7256),
            .I(N__7253));
    Odrv12 I__1547 (
            .O(N__7253),
            .I(CMA_c_9));
    InMux I__1546 (
            .O(N__7250),
            .I(N__7247));
    LocalMux I__1545 (
            .O(N__7247),
            .I(N__7244));
    Odrv4 I__1544 (
            .O(N__7244),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    InMux I__1543 (
            .O(N__7241),
            .I(N__7238));
    LocalMux I__1542 (
            .O(N__7238),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__1541 (
            .O(N__7235),
            .I(N__7232));
    LocalMux I__1540 (
            .O(N__7232),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_3 ));
    InMux I__1539 (
            .O(N__7229),
            .I(N__7226));
    LocalMux I__1538 (
            .O(N__7226),
            .I(N__7223));
    Span12Mux_v I__1537 (
            .O(N__7223),
            .I(N__7220));
    Span12Mux_h I__1536 (
            .O(N__7220),
            .I(N__7217));
    Odrv12 I__1535 (
            .O(N__7217),
            .I(A_c_3));
    InMux I__1534 (
            .O(N__7214),
            .I(N__7211));
    LocalMux I__1533 (
            .O(N__7211),
            .I(N__7208));
    Span12Mux_v I__1532 (
            .O(N__7208),
            .I(N__7205));
    Span12Mux_h I__1531 (
            .O(N__7205),
            .I(N__7202));
    Odrv12 I__1530 (
            .O(N__7202),
            .I(A_c_10));
    CascadeMux I__1529 (
            .O(N__7199),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_ ));
    InMux I__1528 (
            .O(N__7196),
            .I(N__7193));
    LocalMux I__1527 (
            .O(N__7193),
            .I(N__7190));
    Odrv4 I__1526 (
            .O(N__7190),
            .I(\U712_CHIP_RAM.N_33 ));
    InMux I__1525 (
            .O(N__7187),
            .I(N__7184));
    LocalMux I__1524 (
            .O(N__7184),
            .I(N__7181));
    Span4Mux_v I__1523 (
            .O(N__7181),
            .I(N__7178));
    Sp12to4 I__1522 (
            .O(N__7178),
            .I(N__7175));
    Span12Mux_h I__1521 (
            .O(N__7175),
            .I(N__7172));
    Odrv12 I__1520 (
            .O(N__7172),
            .I(A_c_9));
    InMux I__1519 (
            .O(N__7169),
            .I(N__7166));
    LocalMux I__1518 (
            .O(N__7166),
            .I(N__7163));
    Span4Mux_v I__1517 (
            .O(N__7163),
            .I(N__7160));
    Sp12to4 I__1516 (
            .O(N__7160),
            .I(N__7157));
    Span12Mux_h I__1515 (
            .O(N__7157),
            .I(N__7154));
    Span12Mux_v I__1514 (
            .O(N__7154),
            .I(N__7151));
    Odrv12 I__1513 (
            .O(N__7151),
            .I(A_c_2));
    CascadeMux I__1512 (
            .O(N__7148),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_ ));
    InMux I__1511 (
            .O(N__7145),
            .I(N__7142));
    LocalMux I__1510 (
            .O(N__7142),
            .I(N__7139));
    Odrv12 I__1509 (
            .O(N__7139),
            .I(\U712_CHIP_RAM.N_32 ));
    InMux I__1508 (
            .O(N__7136),
            .I(N__7129));
    InMux I__1507 (
            .O(N__7135),
            .I(N__7126));
    CascadeMux I__1506 (
            .O(N__7134),
            .I(N__7123));
    InMux I__1505 (
            .O(N__7133),
            .I(N__7120));
    CascadeMux I__1504 (
            .O(N__7132),
            .I(N__7117));
    LocalMux I__1503 (
            .O(N__7129),
            .I(N__7112));
    LocalMux I__1502 (
            .O(N__7126),
            .I(N__7112));
    InMux I__1501 (
            .O(N__7123),
            .I(N__7109));
    LocalMux I__1500 (
            .O(N__7120),
            .I(N__7106));
    InMux I__1499 (
            .O(N__7117),
            .I(N__7103));
    Span4Mux_h I__1498 (
            .O(N__7112),
            .I(N__7100));
    LocalMux I__1497 (
            .O(N__7109),
            .I(N__7095));
    Span4Mux_h I__1496 (
            .O(N__7106),
            .I(N__7095));
    LocalMux I__1495 (
            .O(N__7103),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1494 (
            .O(N__7100),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1493 (
            .O(N__7095),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    InMux I__1492 (
            .O(N__7088),
            .I(N__7085));
    LocalMux I__1491 (
            .O(N__7085),
            .I(N__7082));
    Odrv12 I__1490 (
            .O(N__7082),
            .I(\U712_BYTE_ENABLE.un2_CUMBEnZ0 ));
    InMux I__1489 (
            .O(N__7079),
            .I(N__7075));
    InMux I__1488 (
            .O(N__7078),
            .I(N__7071));
    LocalMux I__1487 (
            .O(N__7075),
            .I(N__7068));
    InMux I__1486 (
            .O(N__7074),
            .I(N__7065));
    LocalMux I__1485 (
            .O(N__7071),
            .I(N__7062));
    Span4Mux_h I__1484 (
            .O(N__7068),
            .I(N__7057));
    LocalMux I__1483 (
            .O(N__7065),
            .I(N__7057));
    Sp12to4 I__1482 (
            .O(N__7062),
            .I(N__7054));
    Sp12to4 I__1481 (
            .O(N__7057),
            .I(N__7051));
    Span12Mux_v I__1480 (
            .O(N__7054),
            .I(N__7048));
    Span12Mux_h I__1479 (
            .O(N__7051),
            .I(N__7045));
    Span12Mux_h I__1478 (
            .O(N__7048),
            .I(N__7040));
    Span12Mux_v I__1477 (
            .O(N__7045),
            .I(N__7040));
    Odrv12 I__1476 (
            .O(N__7040),
            .I(CASLn_c));
    IoInMux I__1475 (
            .O(N__7037),
            .I(N__7034));
    LocalMux I__1474 (
            .O(N__7034),
            .I(N__7031));
    Span4Mux_s2_h I__1473 (
            .O(N__7031),
            .I(N__7028));
    Sp12to4 I__1472 (
            .O(N__7028),
            .I(N__7025));
    Span12Mux_s5_v I__1471 (
            .O(N__7025),
            .I(N__7022));
    Span12Mux_h I__1470 (
            .O(N__7022),
            .I(N__7019));
    Odrv12 I__1469 (
            .O(N__7019),
            .I(CUMBEn_c));
    InMux I__1468 (
            .O(N__7016),
            .I(N__7011));
    InMux I__1467 (
            .O(N__7015),
            .I(N__7008));
    InMux I__1466 (
            .O(N__7014),
            .I(N__7005));
    LocalMux I__1465 (
            .O(N__7011),
            .I(N__7000));
    LocalMux I__1464 (
            .O(N__7008),
            .I(N__7000));
    LocalMux I__1463 (
            .O(N__7005),
            .I(N__6996));
    Span4Mux_h I__1462 (
            .O(N__7000),
            .I(N__6993));
    InMux I__1461 (
            .O(N__6999),
            .I(N__6990));
    Odrv4 I__1460 (
            .O(N__6996),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0 ));
    Odrv4 I__1459 (
            .O(N__6993),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0 ));
    LocalMux I__1458 (
            .O(N__6990),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0 ));
    InMux I__1457 (
            .O(N__6983),
            .I(N__6978));
    InMux I__1456 (
            .O(N__6982),
            .I(N__6973));
    InMux I__1455 (
            .O(N__6981),
            .I(N__6967));
    LocalMux I__1454 (
            .O(N__6978),
            .I(N__6964));
    InMux I__1453 (
            .O(N__6977),
            .I(N__6961));
    InMux I__1452 (
            .O(N__6976),
            .I(N__6958));
    LocalMux I__1451 (
            .O(N__6973),
            .I(N__6955));
    InMux I__1450 (
            .O(N__6972),
            .I(N__6952));
    InMux I__1449 (
            .O(N__6971),
            .I(N__6947));
    InMux I__1448 (
            .O(N__6970),
            .I(N__6947));
    LocalMux I__1447 (
            .O(N__6967),
            .I(\U712_CHIP_RAM.N_45 ));
    Odrv4 I__1446 (
            .O(N__6964),
            .I(\U712_CHIP_RAM.N_45 ));
    LocalMux I__1445 (
            .O(N__6961),
            .I(\U712_CHIP_RAM.N_45 ));
    LocalMux I__1444 (
            .O(N__6958),
            .I(\U712_CHIP_RAM.N_45 ));
    Odrv4 I__1443 (
            .O(N__6955),
            .I(\U712_CHIP_RAM.N_45 ));
    LocalMux I__1442 (
            .O(N__6952),
            .I(\U712_CHIP_RAM.N_45 ));
    LocalMux I__1441 (
            .O(N__6947),
            .I(\U712_CHIP_RAM.N_45 ));
    InMux I__1440 (
            .O(N__6932),
            .I(N__6929));
    LocalMux I__1439 (
            .O(N__6929),
            .I(N__6926));
    Span12Mux_v I__1438 (
            .O(N__6926),
            .I(N__6923));
    Span12Mux_h I__1437 (
            .O(N__6923),
            .I(N__6920));
    Odrv12 I__1436 (
            .O(N__6920),
            .I(A_c_16));
    CascadeMux I__1435 (
            .O(N__6917),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_7_cascade_ ));
    InMux I__1434 (
            .O(N__6914),
            .I(N__6911));
    LocalMux I__1433 (
            .O(N__6911),
            .I(N__6908));
    Span12Mux_v I__1432 (
            .O(N__6908),
            .I(N__6905));
    Span12Mux_h I__1431 (
            .O(N__6905),
            .I(N__6902));
    Odrv12 I__1430 (
            .O(N__6902),
            .I(A_c_18));
    IoInMux I__1429 (
            .O(N__6899),
            .I(N__6896));
    LocalMux I__1428 (
            .O(N__6896),
            .I(N__6893));
    Span4Mux_s2_v I__1427 (
            .O(N__6893),
            .I(N__6890));
    Span4Mux_v I__1426 (
            .O(N__6890),
            .I(N__6887));
    Span4Mux_v I__1425 (
            .O(N__6887),
            .I(N__6884));
    Odrv4 I__1424 (
            .O(N__6884),
            .I(CMA_c_0));
    IoInMux I__1423 (
            .O(N__6881),
            .I(N__6878));
    LocalMux I__1422 (
            .O(N__6878),
            .I(N__6875));
    IoSpan4Mux I__1421 (
            .O(N__6875),
            .I(N__6872));
    Span4Mux_s3_h I__1420 (
            .O(N__6872),
            .I(N__6869));
    Span4Mux_v I__1419 (
            .O(N__6869),
            .I(N__6866));
    Span4Mux_v I__1418 (
            .O(N__6866),
            .I(N__6863));
    Sp12to4 I__1417 (
            .O(N__6863),
            .I(N__6860));
    Odrv12 I__1416 (
            .O(N__6860),
            .I(CMA_c_3));
    InMux I__1415 (
            .O(N__6857),
            .I(N__6854));
    LocalMux I__1414 (
            .O(N__6854),
            .I(N__6851));
    Span4Mux_h I__1413 (
            .O(N__6851),
            .I(N__6848));
    Sp12to4 I__1412 (
            .O(N__6848),
            .I(N__6845));
    Span12Mux_v I__1411 (
            .O(N__6845),
            .I(N__6842));
    Span12Mux_h I__1410 (
            .O(N__6842),
            .I(N__6839));
    Odrv12 I__1409 (
            .O(N__6839),
            .I(A_c_5));
    CascadeMux I__1408 (
            .O(N__6836),
            .I(N__6833));
    InMux I__1407 (
            .O(N__6833),
            .I(N__6830));
    LocalMux I__1406 (
            .O(N__6830),
            .I(N__6827));
    Span12Mux_v I__1405 (
            .O(N__6827),
            .I(N__6824));
    Span12Mux_h I__1404 (
            .O(N__6824),
            .I(N__6821));
    Odrv12 I__1403 (
            .O(N__6821),
            .I(A_c_12));
    InMux I__1402 (
            .O(N__6818),
            .I(N__6815));
    LocalMux I__1401 (
            .O(N__6815),
            .I(\U712_CHIP_RAM.N_35 ));
    CascadeMux I__1400 (
            .O(N__6812),
            .I(N__6809));
    InMux I__1399 (
            .O(N__6809),
            .I(N__6806));
    LocalMux I__1398 (
            .O(N__6806),
            .I(N__6803));
    Span4Mux_v I__1397 (
            .O(N__6803),
            .I(N__6800));
    Span4Mux_v I__1396 (
            .O(N__6800),
            .I(N__6797));
    Sp12to4 I__1395 (
            .O(N__6797),
            .I(N__6794));
    Span12Mux_h I__1394 (
            .O(N__6794),
            .I(N__6791));
    Odrv12 I__1393 (
            .O(N__6791),
            .I(A_c_7));
    InMux I__1392 (
            .O(N__6788),
            .I(N__6785));
    LocalMux I__1391 (
            .O(N__6785),
            .I(N__6782));
    Span12Mux_v I__1390 (
            .O(N__6782),
            .I(N__6779));
    Span12Mux_h I__1389 (
            .O(N__6779),
            .I(N__6776));
    Odrv12 I__1388 (
            .O(N__6776),
            .I(A_c_14));
    InMux I__1387 (
            .O(N__6773),
            .I(N__6770));
    LocalMux I__1386 (
            .O(N__6770),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_5 ));
    CEMux I__1385 (
            .O(N__6767),
            .I(N__6764));
    LocalMux I__1384 (
            .O(N__6764),
            .I(N__6761));
    Odrv12 I__1383 (
            .O(N__6761),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0 ));
    InMux I__1382 (
            .O(N__6758),
            .I(N__6753));
    InMux I__1381 (
            .O(N__6757),
            .I(N__6750));
    InMux I__1380 (
            .O(N__6756),
            .I(N__6747));
    LocalMux I__1379 (
            .O(N__6753),
            .I(N__6740));
    LocalMux I__1378 (
            .O(N__6750),
            .I(N__6740));
    LocalMux I__1377 (
            .O(N__6747),
            .I(N__6737));
    InMux I__1376 (
            .O(N__6746),
            .I(N__6731));
    InMux I__1375 (
            .O(N__6745),
            .I(N__6731));
    Span4Mux_v I__1374 (
            .O(N__6740),
            .I(N__6728));
    Span4Mux_v I__1373 (
            .O(N__6737),
            .I(N__6725));
    InMux I__1372 (
            .O(N__6736),
            .I(N__6722));
    LocalMux I__1371 (
            .O(N__6731),
            .I(N__6719));
    Sp12to4 I__1370 (
            .O(N__6728),
            .I(N__6712));
    Sp12to4 I__1369 (
            .O(N__6725),
            .I(N__6712));
    LocalMux I__1368 (
            .O(N__6722),
            .I(N__6712));
    Span12Mux_h I__1367 (
            .O(N__6719),
            .I(N__6709));
    Span12Mux_h I__1366 (
            .O(N__6712),
            .I(N__6706));
    Span12Mux_v I__1365 (
            .O(N__6709),
            .I(N__6703));
    Span12Mux_v I__1364 (
            .O(N__6706),
            .I(N__6700));
    Odrv12 I__1363 (
            .O(N__6703),
            .I(RnW_c));
    Odrv12 I__1362 (
            .O(N__6700),
            .I(RnW_c));
    IoInMux I__1361 (
            .O(N__6695),
            .I(N__6692));
    LocalMux I__1360 (
            .O(N__6692),
            .I(N__6689));
    Span4Mux_s3_v I__1359 (
            .O(N__6689),
            .I(N__6686));
    Span4Mux_h I__1358 (
            .O(N__6686),
            .I(N__6683));
    Sp12to4 I__1357 (
            .O(N__6683),
            .I(N__6679));
    CascadeMux I__1356 (
            .O(N__6682),
            .I(N__6675));
    Span12Mux_s10_v I__1355 (
            .O(N__6679),
            .I(N__6672));
    InMux I__1354 (
            .O(N__6678),
            .I(N__6669));
    InMux I__1353 (
            .O(N__6675),
            .I(N__6666));
    Odrv12 I__1352 (
            .O(N__6672),
            .I(DBDIR_c));
    LocalMux I__1351 (
            .O(N__6669),
            .I(DBDIR_c));
    LocalMux I__1350 (
            .O(N__6666),
            .I(DBDIR_c));
    IoInMux I__1349 (
            .O(N__6659),
            .I(N__6656));
    LocalMux I__1348 (
            .O(N__6656),
            .I(N__6653));
    IoSpan4Mux I__1347 (
            .O(N__6653),
            .I(N__6650));
    IoSpan4Mux I__1346 (
            .O(N__6650),
            .I(N__6647));
    Span4Mux_s2_v I__1345 (
            .O(N__6647),
            .I(N__6644));
    Sp12to4 I__1344 (
            .O(N__6644),
            .I(N__6641));
    Span12Mux_v I__1343 (
            .O(N__6641),
            .I(N__6638));
    Odrv12 I__1342 (
            .O(N__6638),
            .I(DRDDIR_0_i));
    CascadeMux I__1341 (
            .O(N__6635),
            .I(N__6632));
    InMux I__1340 (
            .O(N__6632),
            .I(N__6621));
    InMux I__1339 (
            .O(N__6631),
            .I(N__6618));
    InMux I__1338 (
            .O(N__6630),
            .I(N__6609));
    InMux I__1337 (
            .O(N__6629),
            .I(N__6609));
    InMux I__1336 (
            .O(N__6628),
            .I(N__6609));
    InMux I__1335 (
            .O(N__6627),
            .I(N__6609));
    InMux I__1334 (
            .O(N__6626),
            .I(N__6606));
    InMux I__1333 (
            .O(N__6625),
            .I(N__6603));
    InMux I__1332 (
            .O(N__6624),
            .I(N__6600));
    LocalMux I__1331 (
            .O(N__6621),
            .I(N__6591));
    LocalMux I__1330 (
            .O(N__6618),
            .I(N__6591));
    LocalMux I__1329 (
            .O(N__6609),
            .I(N__6591));
    LocalMux I__1328 (
            .O(N__6606),
            .I(N__6591));
    LocalMux I__1327 (
            .O(N__6603),
            .I(N__6588));
    LocalMux I__1326 (
            .O(N__6600),
            .I(N__6584));
    Span4Mux_v I__1325 (
            .O(N__6591),
            .I(N__6581));
    Span4Mux_v I__1324 (
            .O(N__6588),
            .I(N__6578));
    InMux I__1323 (
            .O(N__6587),
            .I(N__6575));
    Span12Mux_v I__1322 (
            .O(N__6584),
            .I(N__6570));
    Sp12to4 I__1321 (
            .O(N__6581),
            .I(N__6570));
    Sp12to4 I__1320 (
            .O(N__6578),
            .I(N__6565));
    LocalMux I__1319 (
            .O(N__6575),
            .I(N__6565));
    Span12Mux_h I__1318 (
            .O(N__6570),
            .I(N__6562));
    Span12Mux_h I__1317 (
            .O(N__6565),
            .I(N__6559));
    Odrv12 I__1316 (
            .O(N__6562),
            .I(RESETn_c));
    Odrv12 I__1315 (
            .O(N__6559),
            .I(RESETn_c));
    IoInMux I__1314 (
            .O(N__6554),
            .I(N__6551));
    LocalMux I__1313 (
            .O(N__6551),
            .I(N__6548));
    Span12Mux_s2_v I__1312 (
            .O(N__6548),
            .I(N__6545));
    Odrv12 I__1311 (
            .O(N__6545),
            .I(RESETn_c_i));
    IoInMux I__1310 (
            .O(N__6542),
            .I(N__6539));
    LocalMux I__1309 (
            .O(N__6539),
            .I(N__6536));
    Span4Mux_s0_v I__1308 (
            .O(N__6536),
            .I(N__6533));
    Span4Mux_v I__1307 (
            .O(N__6533),
            .I(N__6530));
    Span4Mux_v I__1306 (
            .O(N__6530),
            .I(N__6527));
    Span4Mux_h I__1305 (
            .O(N__6527),
            .I(N__6524));
    Odrv4 I__1304 (
            .O(N__6524),
            .I(CRCSn_c));
    InMux I__1303 (
            .O(N__6521),
            .I(N__6517));
    InMux I__1302 (
            .O(N__6520),
            .I(N__6514));
    LocalMux I__1301 (
            .O(N__6517),
            .I(N__6511));
    LocalMux I__1300 (
            .O(N__6514),
            .I(N__6508));
    Span4Mux_v I__1299 (
            .O(N__6511),
            .I(N__6502));
    Span4Mux_v I__1298 (
            .O(N__6508),
            .I(N__6502));
    InMux I__1297 (
            .O(N__6507),
            .I(N__6497));
    Span4Mux_h I__1296 (
            .O(N__6502),
            .I(N__6494));
    InMux I__1295 (
            .O(N__6501),
            .I(N__6489));
    InMux I__1294 (
            .O(N__6500),
            .I(N__6489));
    LocalMux I__1293 (
            .O(N__6497),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__1292 (
            .O(N__6494),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1291 (
            .O(N__6489),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__1290 (
            .O(N__6482),
            .I(N__6479));
    LocalMux I__1289 (
            .O(N__6479),
            .I(N__6476));
    IoSpan4Mux I__1288 (
            .O(N__6476),
            .I(N__6473));
    Sp12to4 I__1287 (
            .O(N__6473),
            .I(N__6470));
    Span12Mux_s9_v I__1286 (
            .O(N__6470),
            .I(N__6467));
    Odrv12 I__1285 (
            .O(N__6467),
            .I(CMA_c_10));
    IoInMux I__1284 (
            .O(N__6464),
            .I(N__6461));
    LocalMux I__1283 (
            .O(N__6461),
            .I(N__6458));
    Span4Mux_s2_v I__1282 (
            .O(N__6458),
            .I(N__6455));
    Span4Mux_v I__1281 (
            .O(N__6455),
            .I(N__6452));
    Span4Mux_v I__1280 (
            .O(N__6452),
            .I(N__6449));
    Odrv4 I__1279 (
            .O(N__6449),
            .I(CMA_c_1));
    InMux I__1278 (
            .O(N__6446),
            .I(N__6443));
    LocalMux I__1277 (
            .O(N__6443),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__1276 (
            .O(N__6440),
            .I(N__6437));
    LocalMux I__1275 (
            .O(N__6437),
            .I(N__6433));
    InMux I__1274 (
            .O(N__6436),
            .I(N__6430));
    Span4Mux_v I__1273 (
            .O(N__6433),
            .I(N__6427));
    LocalMux I__1272 (
            .O(N__6430),
            .I(N__6424));
    Sp12to4 I__1271 (
            .O(N__6427),
            .I(N__6421));
    Sp12to4 I__1270 (
            .O(N__6424),
            .I(N__6418));
    Span12Mux_h I__1269 (
            .O(N__6421),
            .I(N__6415));
    Span12Mux_v I__1268 (
            .O(N__6418),
            .I(N__6412));
    Span12Mux_v I__1267 (
            .O(N__6415),
            .I(N__6409));
    Span12Mux_h I__1266 (
            .O(N__6412),
            .I(N__6406));
    Odrv12 I__1265 (
            .O(N__6409),
            .I(DRA_c_3));
    Odrv12 I__1264 (
            .O(N__6406),
            .I(DRA_c_3));
    InMux I__1263 (
            .O(N__6401),
            .I(N__6398));
    LocalMux I__1262 (
            .O(N__6398),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    CascadeMux I__1261 (
            .O(N__6395),
            .I(\U712_CHIP_RAM.N_47_cascade_ ));
    InMux I__1260 (
            .O(N__6392),
            .I(N__6389));
    LocalMux I__1259 (
            .O(N__6389),
            .I(N__6386));
    Odrv4 I__1258 (
            .O(N__6386),
            .I(\U712_CHIP_RAM.N_89 ));
    InMux I__1257 (
            .O(N__6383),
            .I(N__6379));
    InMux I__1256 (
            .O(N__6382),
            .I(N__6376));
    LocalMux I__1255 (
            .O(N__6379),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_a2_6_0 ));
    LocalMux I__1254 (
            .O(N__6376),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_a2_6_0 ));
    InMux I__1253 (
            .O(N__6371),
            .I(N__6368));
    LocalMux I__1252 (
            .O(N__6368),
            .I(\U712_CHIP_RAM.N_100 ));
    CascadeMux I__1251 (
            .O(N__6365),
            .I(\U712_CHIP_RAM.N_100_cascade_ ));
    InMux I__1250 (
            .O(N__6362),
            .I(N__6358));
    InMux I__1249 (
            .O(N__6361),
            .I(N__6355));
    LocalMux I__1248 (
            .O(N__6358),
            .I(\U712_CHIP_RAM.N_101 ));
    LocalMux I__1247 (
            .O(N__6355),
            .I(\U712_CHIP_RAM.N_101 ));
    CascadeMux I__1246 (
            .O(N__6350),
            .I(N__6347));
    InMux I__1245 (
            .O(N__6347),
            .I(N__6344));
    LocalMux I__1244 (
            .O(N__6344),
            .I(N__6340));
    InMux I__1243 (
            .O(N__6343),
            .I(N__6337));
    Span4Mux_v I__1242 (
            .O(N__6340),
            .I(N__6334));
    LocalMux I__1241 (
            .O(N__6337),
            .I(N__6331));
    Span4Mux_v I__1240 (
            .O(N__6334),
            .I(N__6328));
    Span4Mux_v I__1239 (
            .O(N__6331),
            .I(N__6325));
    Sp12to4 I__1238 (
            .O(N__6328),
            .I(N__6320));
    Sp12to4 I__1237 (
            .O(N__6325),
            .I(N__6320));
    Span12Mux_h I__1236 (
            .O(N__6320),
            .I(N__6317));
    Odrv12 I__1235 (
            .O(N__6317),
            .I(AWEn_c));
    InMux I__1234 (
            .O(N__6314),
            .I(N__6311));
    LocalMux I__1233 (
            .O(N__6311),
            .I(N__6308));
    Odrv4 I__1232 (
            .O(N__6308),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_0_a2_1 ));
    CascadeMux I__1231 (
            .O(N__6305),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_0_cascade_ ));
    InMux I__1230 (
            .O(N__6302),
            .I(N__6298));
    InMux I__1229 (
            .O(N__6301),
            .I(N__6295));
    LocalMux I__1228 (
            .O(N__6298),
            .I(N__6292));
    LocalMux I__1227 (
            .O(N__6295),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    Odrv4 I__1226 (
            .O(N__6292),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    CascadeMux I__1225 (
            .O(N__6287),
            .I(N__6284));
    InMux I__1224 (
            .O(N__6284),
            .I(N__6279));
    CascadeMux I__1223 (
            .O(N__6283),
            .I(N__6276));
    InMux I__1222 (
            .O(N__6282),
            .I(N__6265));
    LocalMux I__1221 (
            .O(N__6279),
            .I(N__6262));
    InMux I__1220 (
            .O(N__6276),
            .I(N__6259));
    InMux I__1219 (
            .O(N__6275),
            .I(N__6256));
    InMux I__1218 (
            .O(N__6274),
            .I(N__6249));
    InMux I__1217 (
            .O(N__6273),
            .I(N__6249));
    InMux I__1216 (
            .O(N__6272),
            .I(N__6249));
    InMux I__1215 (
            .O(N__6271),
            .I(N__6246));
    InMux I__1214 (
            .O(N__6270),
            .I(N__6243));
    InMux I__1213 (
            .O(N__6269),
            .I(N__6238));
    InMux I__1212 (
            .O(N__6268),
            .I(N__6238));
    LocalMux I__1211 (
            .O(N__6265),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv12 I__1210 (
            .O(N__6262),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1209 (
            .O(N__6259),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1208 (
            .O(N__6256),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1207 (
            .O(N__6249),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1206 (
            .O(N__6246),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1205 (
            .O(N__6243),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1204 (
            .O(N__6238),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    CascadeMux I__1203 (
            .O(N__6221),
            .I(N__6217));
    CascadeMux I__1202 (
            .O(N__6220),
            .I(N__6214));
    InMux I__1201 (
            .O(N__6217),
            .I(N__6211));
    InMux I__1200 (
            .O(N__6214),
            .I(N__6208));
    LocalMux I__1199 (
            .O(N__6211),
            .I(N__6205));
    LocalMux I__1198 (
            .O(N__6208),
            .I(N__6194));
    Span4Mux_v I__1197 (
            .O(N__6205),
            .I(N__6191));
    InMux I__1196 (
            .O(N__6204),
            .I(N__6188));
    InMux I__1195 (
            .O(N__6203),
            .I(N__6185));
    InMux I__1194 (
            .O(N__6202),
            .I(N__6182));
    InMux I__1193 (
            .O(N__6201),
            .I(N__6179));
    InMux I__1192 (
            .O(N__6200),
            .I(N__6176));
    InMux I__1191 (
            .O(N__6199),
            .I(N__6173));
    InMux I__1190 (
            .O(N__6198),
            .I(N__6168));
    InMux I__1189 (
            .O(N__6197),
            .I(N__6168));
    Odrv4 I__1188 (
            .O(N__6194),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1187 (
            .O(N__6191),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1186 (
            .O(N__6188),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1185 (
            .O(N__6185),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1184 (
            .O(N__6182),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1183 (
            .O(N__6179),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1182 (
            .O(N__6176),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1181 (
            .O(N__6173),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1180 (
            .O(N__6168),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__1179 (
            .O(N__6149),
            .I(N__6144));
    CascadeMux I__1178 (
            .O(N__6148),
            .I(N__6140));
    CascadeMux I__1177 (
            .O(N__6147),
            .I(N__6137));
    LocalMux I__1176 (
            .O(N__6144),
            .I(N__6134));
    InMux I__1175 (
            .O(N__6143),
            .I(N__6128));
    InMux I__1174 (
            .O(N__6140),
            .I(N__6125));
    InMux I__1173 (
            .O(N__6137),
            .I(N__6122));
    Span4Mux_v I__1172 (
            .O(N__6134),
            .I(N__6119));
    InMux I__1171 (
            .O(N__6133),
            .I(N__6114));
    InMux I__1170 (
            .O(N__6132),
            .I(N__6114));
    InMux I__1169 (
            .O(N__6131),
            .I(N__6111));
    LocalMux I__1168 (
            .O(N__6128),
            .I(\U712_CHIP_RAM.N_56 ));
    LocalMux I__1167 (
            .O(N__6125),
            .I(\U712_CHIP_RAM.N_56 ));
    LocalMux I__1166 (
            .O(N__6122),
            .I(\U712_CHIP_RAM.N_56 ));
    Odrv4 I__1165 (
            .O(N__6119),
            .I(\U712_CHIP_RAM.N_56 ));
    LocalMux I__1164 (
            .O(N__6114),
            .I(\U712_CHIP_RAM.N_56 ));
    LocalMux I__1163 (
            .O(N__6111),
            .I(\U712_CHIP_RAM.N_56 ));
    CascadeMux I__1162 (
            .O(N__6098),
            .I(N__6094));
    InMux I__1161 (
            .O(N__6097),
            .I(N__6090));
    InMux I__1160 (
            .O(N__6094),
            .I(N__6087));
    InMux I__1159 (
            .O(N__6093),
            .I(N__6082));
    LocalMux I__1158 (
            .O(N__6090),
            .I(N__6079));
    LocalMux I__1157 (
            .O(N__6087),
            .I(N__6076));
    InMux I__1156 (
            .O(N__6086),
            .I(N__6071));
    InMux I__1155 (
            .O(N__6085),
            .I(N__6071));
    LocalMux I__1154 (
            .O(N__6082),
            .I(\U712_CHIP_RAM.N_42 ));
    Odrv4 I__1153 (
            .O(N__6079),
            .I(\U712_CHIP_RAM.N_42 ));
    Odrv4 I__1152 (
            .O(N__6076),
            .I(\U712_CHIP_RAM.N_42 ));
    LocalMux I__1151 (
            .O(N__6071),
            .I(\U712_CHIP_RAM.N_42 ));
    CascadeMux I__1150 (
            .O(N__6062),
            .I(N__6053));
    InMux I__1149 (
            .O(N__6061),
            .I(N__6046));
    InMux I__1148 (
            .O(N__6060),
            .I(N__6046));
    InMux I__1147 (
            .O(N__6059),
            .I(N__6035));
    InMux I__1146 (
            .O(N__6058),
            .I(N__6030));
    InMux I__1145 (
            .O(N__6057),
            .I(N__6030));
    InMux I__1144 (
            .O(N__6056),
            .I(N__6027));
    InMux I__1143 (
            .O(N__6053),
            .I(N__6024));
    InMux I__1142 (
            .O(N__6052),
            .I(N__6019));
    InMux I__1141 (
            .O(N__6051),
            .I(N__6019));
    LocalMux I__1140 (
            .O(N__6046),
            .I(N__6016));
    InMux I__1139 (
            .O(N__6045),
            .I(N__6011));
    InMux I__1138 (
            .O(N__6044),
            .I(N__6011));
    InMux I__1137 (
            .O(N__6043),
            .I(N__6006));
    InMux I__1136 (
            .O(N__6042),
            .I(N__6006));
    InMux I__1135 (
            .O(N__6041),
            .I(N__6003));
    InMux I__1134 (
            .O(N__6040),
            .I(N__5996));
    InMux I__1133 (
            .O(N__6039),
            .I(N__5996));
    InMux I__1132 (
            .O(N__6038),
            .I(N__5996));
    LocalMux I__1131 (
            .O(N__6035),
            .I(N__5991));
    LocalMux I__1130 (
            .O(N__6030),
            .I(N__5991));
    LocalMux I__1129 (
            .O(N__6027),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1128 (
            .O(N__6024),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1127 (
            .O(N__6019),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1126 (
            .O(N__6016),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1125 (
            .O(N__6011),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1124 (
            .O(N__6006),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1123 (
            .O(N__6003),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1122 (
            .O(N__5996),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1121 (
            .O(N__5991),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    CascadeMux I__1120 (
            .O(N__5972),
            .I(N__5959));
    InMux I__1119 (
            .O(N__5971),
            .I(N__5953));
    InMux I__1118 (
            .O(N__5970),
            .I(N__5953));
    InMux I__1117 (
            .O(N__5969),
            .I(N__5946));
    InMux I__1116 (
            .O(N__5968),
            .I(N__5946));
    InMux I__1115 (
            .O(N__5967),
            .I(N__5940));
    InMux I__1114 (
            .O(N__5966),
            .I(N__5933));
    InMux I__1113 (
            .O(N__5965),
            .I(N__5933));
    InMux I__1112 (
            .O(N__5964),
            .I(N__5933));
    InMux I__1111 (
            .O(N__5963),
            .I(N__5929));
    InMux I__1110 (
            .O(N__5962),
            .I(N__5924));
    InMux I__1109 (
            .O(N__5959),
            .I(N__5924));
    InMux I__1108 (
            .O(N__5958),
            .I(N__5921));
    LocalMux I__1107 (
            .O(N__5953),
            .I(N__5918));
    InMux I__1106 (
            .O(N__5952),
            .I(N__5913));
    InMux I__1105 (
            .O(N__5951),
            .I(N__5913));
    LocalMux I__1104 (
            .O(N__5946),
            .I(N__5910));
    InMux I__1103 (
            .O(N__5945),
            .I(N__5907));
    InMux I__1102 (
            .O(N__5944),
            .I(N__5902));
    InMux I__1101 (
            .O(N__5943),
            .I(N__5902));
    LocalMux I__1100 (
            .O(N__5940),
            .I(N__5897));
    LocalMux I__1099 (
            .O(N__5933),
            .I(N__5897));
    InMux I__1098 (
            .O(N__5932),
            .I(N__5894));
    LocalMux I__1097 (
            .O(N__5929),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1096 (
            .O(N__5924),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1095 (
            .O(N__5921),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1094 (
            .O(N__5918),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1093 (
            .O(N__5913),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1092 (
            .O(N__5910),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1091 (
            .O(N__5907),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1090 (
            .O(N__5902),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1089 (
            .O(N__5897),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1088 (
            .O(N__5894),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    CascadeMux I__1087 (
            .O(N__5873),
            .I(\U712_CHIP_RAM.N_42_cascade_ ));
    CascadeMux I__1086 (
            .O(N__5870),
            .I(N__5867));
    InMux I__1085 (
            .O(N__5867),
            .I(N__5863));
    InMux I__1084 (
            .O(N__5866),
            .I(N__5856));
    LocalMux I__1083 (
            .O(N__5863),
            .I(N__5853));
    InMux I__1082 (
            .O(N__5862),
            .I(N__5850));
    InMux I__1081 (
            .O(N__5861),
            .I(N__5843));
    InMux I__1080 (
            .O(N__5860),
            .I(N__5843));
    InMux I__1079 (
            .O(N__5859),
            .I(N__5843));
    LocalMux I__1078 (
            .O(N__5856),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1077 (
            .O(N__5853),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1076 (
            .O(N__5850),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1075 (
            .O(N__5843),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__1074 (
            .O(N__5834),
            .I(N__5831));
    LocalMux I__1073 (
            .O(N__5831),
            .I(N__5828));
    Span4Mux_h I__1072 (
            .O(N__5828),
            .I(N__5824));
    InMux I__1071 (
            .O(N__5827),
            .I(N__5821));
    Odrv4 I__1070 (
            .O(N__5824),
            .I(\U712_CHIP_RAM.N_98 ));
    LocalMux I__1069 (
            .O(N__5821),
            .I(\U712_CHIP_RAM.N_98 ));
    InMux I__1068 (
            .O(N__5816),
            .I(N__5813));
    LocalMux I__1067 (
            .O(N__5813),
            .I(N__5810));
    Span12Mux_v I__1066 (
            .O(N__5810),
            .I(N__5807));
    Span12Mux_h I__1065 (
            .O(N__5807),
            .I(N__5804));
    Odrv12 I__1064 (
            .O(N__5804),
            .I(A_c_15));
    CascadeMux I__1063 (
            .O(N__5801),
            .I(N__5798));
    InMux I__1062 (
            .O(N__5798),
            .I(N__5795));
    LocalMux I__1061 (
            .O(N__5795),
            .I(N__5792));
    Span4Mux_v I__1060 (
            .O(N__5792),
            .I(N__5789));
    Span4Mux_v I__1059 (
            .O(N__5789),
            .I(N__5786));
    Sp12to4 I__1058 (
            .O(N__5786),
            .I(N__5783));
    Span12Mux_h I__1057 (
            .O(N__5783),
            .I(N__5780));
    Odrv12 I__1056 (
            .O(N__5780),
            .I(A_c_8));
    InMux I__1055 (
            .O(N__5777),
            .I(N__5774));
    LocalMux I__1054 (
            .O(N__5774),
            .I(\U712_CHIP_RAM.N_38 ));
    InMux I__1053 (
            .O(N__5771),
            .I(N__5768));
    LocalMux I__1052 (
            .O(N__5768),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_6 ));
    InMux I__1051 (
            .O(N__5765),
            .I(N__5759));
    InMux I__1050 (
            .O(N__5764),
            .I(N__5752));
    InMux I__1049 (
            .O(N__5763),
            .I(N__5749));
    InMux I__1048 (
            .O(N__5762),
            .I(N__5746));
    LocalMux I__1047 (
            .O(N__5759),
            .I(N__5743));
    InMux I__1046 (
            .O(N__5758),
            .I(N__5740));
    InMux I__1045 (
            .O(N__5757),
            .I(N__5737));
    InMux I__1044 (
            .O(N__5756),
            .I(N__5732));
    InMux I__1043 (
            .O(N__5755),
            .I(N__5732));
    LocalMux I__1042 (
            .O(N__5752),
            .I(\U712_CHIP_RAM.N_44 ));
    LocalMux I__1041 (
            .O(N__5749),
            .I(\U712_CHIP_RAM.N_44 ));
    LocalMux I__1040 (
            .O(N__5746),
            .I(\U712_CHIP_RAM.N_44 ));
    Odrv4 I__1039 (
            .O(N__5743),
            .I(\U712_CHIP_RAM.N_44 ));
    LocalMux I__1038 (
            .O(N__5740),
            .I(\U712_CHIP_RAM.N_44 ));
    LocalMux I__1037 (
            .O(N__5737),
            .I(\U712_CHIP_RAM.N_44 ));
    LocalMux I__1036 (
            .O(N__5732),
            .I(\U712_CHIP_RAM.N_44 ));
    InMux I__1035 (
            .O(N__5717),
            .I(N__5714));
    LocalMux I__1034 (
            .O(N__5714),
            .I(N__5710));
    InMux I__1033 (
            .O(N__5713),
            .I(N__5707));
    Span4Mux_v I__1032 (
            .O(N__5710),
            .I(N__5704));
    LocalMux I__1031 (
            .O(N__5707),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    Odrv4 I__1030 (
            .O(N__5704),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__1029 (
            .O(N__5699),
            .I(N__5696));
    LocalMux I__1028 (
            .O(N__5696),
            .I(N__5693));
    Span4Mux_h I__1027 (
            .O(N__5693),
            .I(N__5690));
    Odrv4 I__1026 (
            .O(N__5690),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ));
    CascadeMux I__1025 (
            .O(N__5687),
            .I(N__5684));
    InMux I__1024 (
            .O(N__5684),
            .I(N__5681));
    LocalMux I__1023 (
            .O(N__5681),
            .I(N__5677));
    InMux I__1022 (
            .O(N__5680),
            .I(N__5674));
    Span4Mux_h I__1021 (
            .O(N__5677),
            .I(N__5671));
    LocalMux I__1020 (
            .O(N__5674),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    Odrv4 I__1019 (
            .O(N__5671),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__1018 (
            .O(N__5666),
            .I(N__5663));
    LocalMux I__1017 (
            .O(N__5663),
            .I(N__5660));
    Span4Mux_h I__1016 (
            .O(N__5660),
            .I(N__5657));
    Odrv4 I__1015 (
            .O(N__5657),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ));
    InMux I__1014 (
            .O(N__5654),
            .I(N__5651));
    LocalMux I__1013 (
            .O(N__5651),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    CascadeMux I__1012 (
            .O(N__5648),
            .I(N__5645));
    InMux I__1011 (
            .O(N__5645),
            .I(N__5641));
    InMux I__1010 (
            .O(N__5644),
            .I(N__5638));
    LocalMux I__1009 (
            .O(N__5641),
            .I(N__5635));
    LocalMux I__1008 (
            .O(N__5638),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_0 ));
    Odrv4 I__1007 (
            .O(N__5635),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_0 ));
    InMux I__1006 (
            .O(N__5630),
            .I(N__5626));
    InMux I__1005 (
            .O(N__5629),
            .I(N__5623));
    LocalMux I__1004 (
            .O(N__5626),
            .I(\U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ));
    LocalMux I__1003 (
            .O(N__5623),
            .I(\U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ));
    InMux I__1002 (
            .O(N__5618),
            .I(N__5613));
    InMux I__1001 (
            .O(N__5617),
            .I(N__5608));
    InMux I__1000 (
            .O(N__5616),
            .I(N__5608));
    LocalMux I__999 (
            .O(N__5613),
            .I(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ));
    LocalMux I__998 (
            .O(N__5608),
            .I(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ));
    InMux I__997 (
            .O(N__5603),
            .I(N__5599));
    InMux I__996 (
            .O(N__5602),
            .I(N__5596));
    LocalMux I__995 (
            .O(N__5599),
            .I(\U712_CHIP_RAM.N_47 ));
    LocalMux I__994 (
            .O(N__5596),
            .I(\U712_CHIP_RAM.N_47 ));
    InMux I__993 (
            .O(N__5591),
            .I(N__5588));
    LocalMux I__992 (
            .O(N__5588),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6 ));
    InMux I__991 (
            .O(N__5585),
            .I(N__5580));
    InMux I__990 (
            .O(N__5584),
            .I(N__5575));
    InMux I__989 (
            .O(N__5583),
            .I(N__5575));
    LocalMux I__988 (
            .O(N__5580),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__987 (
            .O(N__5575),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    CascadeMux I__986 (
            .O(N__5570),
            .I(N__5566));
    InMux I__985 (
            .O(N__5569),
            .I(N__5563));
    InMux I__984 (
            .O(N__5566),
            .I(N__5560));
    LocalMux I__983 (
            .O(N__5563),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__982 (
            .O(N__5560),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__981 (
            .O(N__5555),
            .I(N__5552));
    LocalMux I__980 (
            .O(N__5552),
            .I(N__5548));
    InMux I__979 (
            .O(N__5551),
            .I(N__5545));
    Odrv4 I__978 (
            .O(N__5548),
            .I(\U712_CHIP_RAM.N_57 ));
    LocalMux I__977 (
            .O(N__5545),
            .I(\U712_CHIP_RAM.N_57 ));
    InMux I__976 (
            .O(N__5540),
            .I(N__5537));
    LocalMux I__975 (
            .O(N__5537),
            .I(\U712_BYTE_ENABLE.un2_CLLBEnZ0 ));
    IoInMux I__974 (
            .O(N__5534),
            .I(N__5531));
    LocalMux I__973 (
            .O(N__5531),
            .I(N__5528));
    IoSpan4Mux I__972 (
            .O(N__5528),
            .I(N__5525));
    Span4Mux_s2_v I__971 (
            .O(N__5525),
            .I(N__5522));
    Sp12to4 I__970 (
            .O(N__5522),
            .I(N__5519));
    Span12Mux_v I__969 (
            .O(N__5519),
            .I(N__5516));
    Odrv12 I__968 (
            .O(N__5516),
            .I(CLLBEn_c));
    InMux I__967 (
            .O(N__5513),
            .I(N__5510));
    LocalMux I__966 (
            .O(N__5510),
            .I(\U712_CHIP_RAM.DMA_CYCLE_7 ));
    InMux I__965 (
            .O(N__5507),
            .I(N__5504));
    LocalMux I__964 (
            .O(N__5504),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_0 ));
    IoInMux I__963 (
            .O(N__5501),
            .I(N__5498));
    LocalMux I__962 (
            .O(N__5498),
            .I(N__5495));
    IoSpan4Mux I__961 (
            .O(N__5495),
            .I(N__5492));
    IoSpan4Mux I__960 (
            .O(N__5492),
            .I(N__5489));
    Sp12to4 I__959 (
            .O(N__5489),
            .I(N__5486));
    Span12Mux_s9_h I__958 (
            .O(N__5486),
            .I(N__5483));
    Odrv12 I__957 (
            .O(N__5483),
            .I(CMA_c_6));
    InMux I__956 (
            .O(N__5480),
            .I(N__5477));
    LocalMux I__955 (
            .O(N__5477),
            .I(N__5474));
    Odrv4 I__954 (
            .O(N__5474),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i ));
    CascadeMux I__953 (
            .O(N__5471),
            .I(\U712_CHIP_RAM.N_44_cascade_ ));
    InMux I__952 (
            .O(N__5468),
            .I(N__5463));
    InMux I__951 (
            .O(N__5467),
            .I(N__5460));
    InMux I__950 (
            .O(N__5466),
            .I(N__5457));
    LocalMux I__949 (
            .O(N__5463),
            .I(\U712_CHIP_RAM.N_93 ));
    LocalMux I__948 (
            .O(N__5460),
            .I(\U712_CHIP_RAM.N_93 ));
    LocalMux I__947 (
            .O(N__5457),
            .I(\U712_CHIP_RAM.N_93 ));
    InMux I__946 (
            .O(N__5450),
            .I(N__5446));
    InMux I__945 (
            .O(N__5449),
            .I(N__5443));
    LocalMux I__944 (
            .O(N__5446),
            .I(\U712_CHIP_RAM.N_13 ));
    LocalMux I__943 (
            .O(N__5443),
            .I(\U712_CHIP_RAM.N_13 ));
    InMux I__942 (
            .O(N__5438),
            .I(N__5435));
    LocalMux I__941 (
            .O(N__5435),
            .I(\U712_CHIP_RAM.N_65 ));
    CascadeMux I__940 (
            .O(N__5432),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_i_1_0_cascade_ ));
    InMux I__939 (
            .O(N__5429),
            .I(N__5426));
    LocalMux I__938 (
            .O(N__5426),
            .I(\U712_CHIP_RAM.N_62 ));
    InMux I__937 (
            .O(N__5423),
            .I(N__5417));
    InMux I__936 (
            .O(N__5422),
            .I(N__5414));
    InMux I__935 (
            .O(N__5421),
            .I(N__5409));
    InMux I__934 (
            .O(N__5420),
            .I(N__5409));
    LocalMux I__933 (
            .O(N__5417),
            .I(N__5402));
    LocalMux I__932 (
            .O(N__5414),
            .I(N__5402));
    LocalMux I__931 (
            .O(N__5409),
            .I(N__5402));
    Odrv4 I__930 (
            .O(N__5402),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3 ));
    InMux I__929 (
            .O(N__5399),
            .I(N__5394));
    InMux I__928 (
            .O(N__5398),
            .I(N__5389));
    InMux I__927 (
            .O(N__5397),
            .I(N__5389));
    LocalMux I__926 (
            .O(N__5394),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__925 (
            .O(N__5389),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__924 (
            .O(N__5384),
            .I(N__5381));
    InMux I__923 (
            .O(N__5381),
            .I(N__5375));
    InMux I__922 (
            .O(N__5380),
            .I(N__5368));
    InMux I__921 (
            .O(N__5379),
            .I(N__5368));
    InMux I__920 (
            .O(N__5378),
            .I(N__5368));
    LocalMux I__919 (
            .O(N__5375),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__918 (
            .O(N__5368),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    CascadeMux I__917 (
            .O(N__5363),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6_cascade_ ));
    InMux I__916 (
            .O(N__5360),
            .I(N__5350));
    InMux I__915 (
            .O(N__5359),
            .I(N__5350));
    InMux I__914 (
            .O(N__5358),
            .I(N__5350));
    InMux I__913 (
            .O(N__5357),
            .I(N__5347));
    LocalMux I__912 (
            .O(N__5350),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ));
    LocalMux I__911 (
            .O(N__5347),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ));
    InMux I__910 (
            .O(N__5342),
            .I(N__5339));
    LocalMux I__909 (
            .O(N__5339),
            .I(\U712_CHIP_RAM.N_75 ));
    InMux I__908 (
            .O(N__5336),
            .I(N__5332));
    InMux I__907 (
            .O(N__5335),
            .I(N__5329));
    LocalMux I__906 (
            .O(N__5332),
            .I(\U712_CHIP_RAM.N_60 ));
    LocalMux I__905 (
            .O(N__5329),
            .I(\U712_CHIP_RAM.N_60 ));
    InMux I__904 (
            .O(N__5324),
            .I(N__5321));
    LocalMux I__903 (
            .O(N__5321),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_1 ));
    InMux I__902 (
            .O(N__5318),
            .I(N__5315));
    LocalMux I__901 (
            .O(N__5315),
            .I(\U712_CHIP_RAM.N_77 ));
    InMux I__900 (
            .O(N__5312),
            .I(N__5309));
    LocalMux I__899 (
            .O(N__5309),
            .I(\U712_CHIP_RAM.N_40 ));
    CascadeMux I__898 (
            .O(N__5306),
            .I(\U712_CHIP_RAM.N_62_cascade_ ));
    CascadeMux I__897 (
            .O(N__5303),
            .I(\U712_CHIP_RAM.N_13_cascade_ ));
    InMux I__896 (
            .O(N__5300),
            .I(N__5297));
    LocalMux I__895 (
            .O(N__5297),
            .I(N__5294));
    Span4Mux_v I__894 (
            .O(N__5294),
            .I(N__5291));
    Sp12to4 I__893 (
            .O(N__5291),
            .I(N__5288));
    Span12Mux_h I__892 (
            .O(N__5288),
            .I(N__5285));
    Span12Mux_v I__891 (
            .O(N__5285),
            .I(N__5282));
    Odrv12 I__890 (
            .O(N__5282),
            .I(A_c_4));
    CascadeMux I__889 (
            .O(N__5279),
            .I(N__5276));
    InMux I__888 (
            .O(N__5276),
            .I(N__5273));
    LocalMux I__887 (
            .O(N__5273),
            .I(N__5270));
    Span4Mux_v I__886 (
            .O(N__5270),
            .I(N__5267));
    Sp12to4 I__885 (
            .O(N__5267),
            .I(N__5264));
    Span12Mux_h I__884 (
            .O(N__5264),
            .I(N__5261));
    Odrv12 I__883 (
            .O(N__5261),
            .I(A_c_11));
    InMux I__882 (
            .O(N__5258),
            .I(N__5255));
    LocalMux I__881 (
            .O(N__5255),
            .I(\U712_CHIP_RAM.N_34 ));
    InMux I__880 (
            .O(N__5252),
            .I(N__5249));
    LocalMux I__879 (
            .O(N__5249),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__878 (
            .O(N__5246),
            .I(N__5243));
    LocalMux I__877 (
            .O(N__5243),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_2 ));
    InMux I__876 (
            .O(N__5240),
            .I(N__5237));
    LocalMux I__875 (
            .O(N__5237),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    SRMux I__874 (
            .O(N__5234),
            .I(N__5231));
    LocalMux I__873 (
            .O(N__5231),
            .I(N__5228));
    Odrv4 I__872 (
            .O(N__5228),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    CascadeMux I__871 (
            .O(N__5225),
            .I(\U712_CHIP_RAM.N_74_cascade_ ));
    CascadeMux I__870 (
            .O(N__5222),
            .I(\U712_CHIP_RAM.N_50_cascade_ ));
    CascadeMux I__869 (
            .O(N__5219),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_ ));
    InMux I__868 (
            .O(N__5216),
            .I(N__5213));
    LocalMux I__867 (
            .O(N__5213),
            .I(\U712_CHIP_RAM.N_58 ));
    CascadeMux I__866 (
            .O(N__5210),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_a2_0_cascade_ ));
    InMux I__865 (
            .O(N__5207),
            .I(N__5204));
    LocalMux I__864 (
            .O(N__5204),
            .I(N__5200));
    InMux I__863 (
            .O(N__5203),
            .I(N__5197));
    Span12Mux_h I__862 (
            .O(N__5200),
            .I(N__5192));
    LocalMux I__861 (
            .O(N__5197),
            .I(N__5192));
    Span12Mux_h I__860 (
            .O(N__5192),
            .I(N__5189));
    Span12Mux_v I__859 (
            .O(N__5189),
            .I(N__5186));
    Odrv12 I__858 (
            .O(N__5186),
            .I(SIZ_c_1));
    InMux I__857 (
            .O(N__5183),
            .I(N__5173));
    InMux I__856 (
            .O(N__5182),
            .I(N__5173));
    InMux I__855 (
            .O(N__5181),
            .I(N__5173));
    InMux I__854 (
            .O(N__5180),
            .I(N__5170));
    LocalMux I__853 (
            .O(N__5173),
            .I(N__5165));
    LocalMux I__852 (
            .O(N__5170),
            .I(N__5165));
    Span4Mux_h I__851 (
            .O(N__5165),
            .I(N__5161));
    InMux I__850 (
            .O(N__5164),
            .I(N__5158));
    Span4Mux_v I__849 (
            .O(N__5161),
            .I(N__5155));
    LocalMux I__848 (
            .O(N__5158),
            .I(N__5152));
    Sp12to4 I__847 (
            .O(N__5155),
            .I(N__5147));
    Span12Mux_v I__846 (
            .O(N__5152),
            .I(N__5147));
    Odrv12 I__845 (
            .O(N__5147),
            .I(A_c_0));
    InMux I__844 (
            .O(N__5144),
            .I(N__5141));
    LocalMux I__843 (
            .O(N__5141),
            .I(\U712_BYTE_ENABLE.LLBE_0_0_tz ));
    InMux I__842 (
            .O(N__5138),
            .I(N__5132));
    InMux I__841 (
            .O(N__5137),
            .I(N__5125));
    InMux I__840 (
            .O(N__5136),
            .I(N__5125));
    InMux I__839 (
            .O(N__5135),
            .I(N__5125));
    LocalMux I__838 (
            .O(N__5132),
            .I(\U712_BYTE_ENABLE.LW_TRANS_0 ));
    LocalMux I__837 (
            .O(N__5125),
            .I(\U712_BYTE_ENABLE.LW_TRANS_0 ));
    CascadeMux I__836 (
            .O(N__5120),
            .I(\U712_BYTE_ENABLE.LLBE_0_0_tz_cascade_ ));
    CascadeMux I__835 (
            .O(N__5117),
            .I(N__5114));
    InMux I__834 (
            .O(N__5114),
            .I(N__5110));
    CascadeMux I__833 (
            .O(N__5113),
            .I(N__5106));
    LocalMux I__832 (
            .O(N__5110),
            .I(N__5102));
    InMux I__831 (
            .O(N__5109),
            .I(N__5095));
    InMux I__830 (
            .O(N__5106),
            .I(N__5095));
    InMux I__829 (
            .O(N__5105),
            .I(N__5095));
    Span4Mux_h I__828 (
            .O(N__5102),
            .I(N__5090));
    LocalMux I__827 (
            .O(N__5095),
            .I(N__5090));
    Span4Mux_v I__826 (
            .O(N__5090),
            .I(N__5087));
    Span4Mux_v I__825 (
            .O(N__5087),
            .I(N__5084));
    Sp12to4 I__824 (
            .O(N__5084),
            .I(N__5081));
    Span12Mux_h I__823 (
            .O(N__5081),
            .I(N__5078));
    Odrv12 I__822 (
            .O(N__5078),
            .I(A_c_1));
    IoInMux I__821 (
            .O(N__5075),
            .I(N__5072));
    LocalMux I__820 (
            .O(N__5072),
            .I(N__5069));
    Odrv12 I__819 (
            .O(N__5069),
            .I(CMA_c_2));
    CascadeMux I__818 (
            .O(N__5066),
            .I(\U712_CHIP_RAM.N_58_cascade_ ));
    CascadeMux I__817 (
            .O(N__5063),
            .I(\U712_CHIP_RAM.N_40_cascade_ ));
    InMux I__816 (
            .O(N__5060),
            .I(N__5057));
    LocalMux I__815 (
            .O(N__5057),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_0 ));
    CascadeMux I__814 (
            .O(N__5054),
            .I(\U712_CHIP_RAM.N_99_cascade_ ));
    InMux I__813 (
            .O(N__5051),
            .I(N__5048));
    LocalMux I__812 (
            .O(N__5048),
            .I(\U712_CHIP_RAM.N_85 ));
    CascadeMux I__811 (
            .O(N__5045),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_a2_0_cascade_ ));
    InMux I__810 (
            .O(N__5042),
            .I(N__5039));
    LocalMux I__809 (
            .O(N__5039),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_a2_0_0 ));
    CascadeMux I__808 (
            .O(N__5036),
            .I(\U712_CHIP_RAM.N_65_cascade_ ));
    InMux I__807 (
            .O(N__5033),
            .I(N__5030));
    LocalMux I__806 (
            .O(N__5030),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0 ));
    CascadeMux I__805 (
            .O(N__5027),
            .I(\U712_CHIP_RAM.N_49_cascade_ ));
    InMux I__804 (
            .O(N__5024),
            .I(N__5020));
    InMux I__803 (
            .O(N__5023),
            .I(N__5017));
    LocalMux I__802 (
            .O(N__5020),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    LocalMux I__801 (
            .O(N__5017),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    InMux I__800 (
            .O(N__5012),
            .I(N__5008));
    InMux I__799 (
            .O(N__5011),
            .I(N__5005));
    LocalMux I__798 (
            .O(N__5008),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__797 (
            .O(N__5005),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    CascadeMux I__796 (
            .O(N__5000),
            .I(N__4996));
    InMux I__795 (
            .O(N__4999),
            .I(N__4993));
    InMux I__794 (
            .O(N__4996),
            .I(N__4990));
    LocalMux I__793 (
            .O(N__4993),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__792 (
            .O(N__4990),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__791 (
            .O(N__4985),
            .I(N__4981));
    InMux I__790 (
            .O(N__4984),
            .I(N__4978));
    LocalMux I__789 (
            .O(N__4981),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ));
    LocalMux I__788 (
            .O(N__4978),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ));
    InMux I__787 (
            .O(N__4973),
            .I(N__4969));
    InMux I__786 (
            .O(N__4972),
            .I(N__4966));
    LocalMux I__785 (
            .O(N__4969),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__784 (
            .O(N__4966),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__783 (
            .O(N__4961),
            .I(N__4957));
    InMux I__782 (
            .O(N__4960),
            .I(N__4954));
    LocalMux I__781 (
            .O(N__4957),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__780 (
            .O(N__4954),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    CascadeMux I__779 (
            .O(N__4949),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_a2_0_0_cascade_ ));
    InMux I__778 (
            .O(N__4946),
            .I(N__4943));
    LocalMux I__777 (
            .O(N__4943),
            .I(N__4939));
    IoInMux I__776 (
            .O(N__4942),
            .I(N__4936));
    Span12Mux_h I__775 (
            .O(N__4939),
            .I(N__4933));
    LocalMux I__774 (
            .O(N__4936),
            .I(N__4930));
    Span12Mux_v I__773 (
            .O(N__4933),
            .I(N__4927));
    IoSpan4Mux I__772 (
            .O(N__4930),
            .I(N__4924));
    Odrv12 I__771 (
            .O(N__4927),
            .I(RAMENn_c));
    Odrv4 I__770 (
            .O(N__4924),
            .I(RAMENn_c));
    CascadeMux I__769 (
            .O(N__4919),
            .I(N__4916));
    InMux I__768 (
            .O(N__4916),
            .I(N__4913));
    LocalMux I__767 (
            .O(N__4913),
            .I(N__4909));
    InMux I__766 (
            .O(N__4912),
            .I(N__4906));
    Span4Mux_v I__765 (
            .O(N__4909),
            .I(N__4900));
    LocalMux I__764 (
            .O(N__4906),
            .I(N__4900));
    InMux I__763 (
            .O(N__4905),
            .I(N__4897));
    Span4Mux_v I__762 (
            .O(N__4900),
            .I(N__4894));
    LocalMux I__761 (
            .O(N__4897),
            .I(N__4891));
    Sp12to4 I__760 (
            .O(N__4894),
            .I(N__4888));
    Span12Mux_h I__759 (
            .O(N__4891),
            .I(N__4885));
    Span12Mux_h I__758 (
            .O(N__4888),
            .I(N__4882));
    Span12Mux_v I__757 (
            .O(N__4885),
            .I(N__4879));
    Span12Mux_v I__756 (
            .O(N__4882),
            .I(N__4876));
    Odrv12 I__755 (
            .O(N__4879),
            .I(TSn_c));
    Odrv12 I__754 (
            .O(N__4876),
            .I(TSn_c));
    InMux I__753 (
            .O(N__4871),
            .I(N__4867));
    InMux I__752 (
            .O(N__4870),
            .I(N__4863));
    LocalMux I__751 (
            .O(N__4867),
            .I(N__4860));
    InMux I__750 (
            .O(N__4866),
            .I(N__4857));
    LocalMux I__749 (
            .O(N__4863),
            .I(U712_REG_SM_DBR_SYNC_1));
    Odrv4 I__748 (
            .O(N__4860),
            .I(U712_REG_SM_DBR_SYNC_1));
    LocalMux I__747 (
            .O(N__4857),
            .I(U712_REG_SM_DBR_SYNC_1));
    CascadeMux I__746 (
            .O(N__4850),
            .I(N__4846));
    InMux I__745 (
            .O(N__4849),
            .I(N__4840));
    InMux I__744 (
            .O(N__4846),
            .I(N__4840));
    CascadeMux I__743 (
            .O(N__4845),
            .I(N__4836));
    LocalMux I__742 (
            .O(N__4840),
            .I(N__4833));
    InMux I__741 (
            .O(N__4839),
            .I(N__4830));
    InMux I__740 (
            .O(N__4836),
            .I(N__4827));
    Odrv12 I__739 (
            .O(N__4833),
            .I(U712_REG_SM_DBR_SYNC_0));
    LocalMux I__738 (
            .O(N__4830),
            .I(U712_REG_SM_DBR_SYNC_0));
    LocalMux I__737 (
            .O(N__4827),
            .I(U712_REG_SM_DBR_SYNC_0));
    InMux I__736 (
            .O(N__4820),
            .I(N__4814));
    InMux I__735 (
            .O(N__4819),
            .I(N__4814));
    LocalMux I__734 (
            .O(N__4814),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    CascadeMux I__733 (
            .O(N__4811),
            .I(\U712_CHIP_RAM.N_57_cascade_ ));
    InMux I__732 (
            .O(N__4808),
            .I(bfn_10_7_0_));
    InMux I__731 (
            .O(N__4805),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__730 (
            .O(N__4802),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__729 (
            .O(N__4799),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__728 (
            .O(N__4796),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__727 (
            .O(N__4793),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__726 (
            .O(N__4790),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__725 (
            .O(N__4787),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    ClkMux I__724 (
            .O(N__4784),
            .I(N__4781));
    GlobalMux I__723 (
            .O(N__4781),
            .I(N__4778));
    gio2CtrlBuf I__722 (
            .O(N__4778),
            .I(C1_c_g));
    InMux I__721 (
            .O(N__4775),
            .I(N__4772));
    LocalMux I__720 (
            .O(N__4772),
            .I(N__4769));
    Span4Mux_v I__719 (
            .O(N__4769),
            .I(N__4766));
    Sp12to4 I__718 (
            .O(N__4766),
            .I(N__4763));
    Span12Mux_h I__717 (
            .O(N__4763),
            .I(N__4760));
    Span12Mux_v I__716 (
            .O(N__4760),
            .I(N__4757));
    Odrv12 I__715 (
            .O(N__4757),
            .I(DBRn_c));
    InMux I__714 (
            .O(N__4754),
            .I(N__4749));
    InMux I__713 (
            .O(N__4753),
            .I(N__4746));
    InMux I__712 (
            .O(N__4752),
            .I(N__4743));
    LocalMux I__711 (
            .O(N__4749),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__710 (
            .O(N__4746),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__709 (
            .O(N__4743),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    CascadeMux I__708 (
            .O(N__4736),
            .I(N__4731));
    InMux I__707 (
            .O(N__4735),
            .I(N__4728));
    InMux I__706 (
            .O(N__4734),
            .I(N__4723));
    InMux I__705 (
            .O(N__4731),
            .I(N__4723));
    LocalMux I__704 (
            .O(N__4728),
            .I(N__4720));
    LocalMux I__703 (
            .O(N__4723),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    Odrv4 I__702 (
            .O(N__4720),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    CEMux I__701 (
            .O(N__4715),
            .I(N__4712));
    LocalMux I__700 (
            .O(N__4712),
            .I(N__4709));
    Span4Mux_h I__699 (
            .O(N__4709),
            .I(N__4706));
    Odrv4 I__698 (
            .O(N__4706),
            .I(\U712_CYCLE_TERM.N_45_0_0_en_0 ));
    InMux I__697 (
            .O(N__4703),
            .I(N__4700));
    LocalMux I__696 (
            .O(N__4700),
            .I(\U712_REG_SM.LDS_OUT_2_0_0 ));
    InMux I__695 (
            .O(N__4697),
            .I(N__4694));
    LocalMux I__694 (
            .O(N__4694),
            .I(N__4690));
    InMux I__693 (
            .O(N__4693),
            .I(N__4686));
    Span4Mux_h I__692 (
            .O(N__4690),
            .I(N__4683));
    InMux I__691 (
            .O(N__4689),
            .I(N__4680));
    LocalMux I__690 (
            .O(N__4686),
            .I(N__4677));
    Odrv4 I__689 (
            .O(N__4683),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__688 (
            .O(N__4680),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    Odrv4 I__687 (
            .O(N__4677),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    InMux I__686 (
            .O(N__4670),
            .I(N__4666));
    InMux I__685 (
            .O(N__4669),
            .I(N__4663));
    LocalMux I__684 (
            .O(N__4666),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    LocalMux I__683 (
            .O(N__4663),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    InMux I__682 (
            .O(N__4658),
            .I(N__4655));
    LocalMux I__681 (
            .O(N__4655),
            .I(N__4652));
    Odrv4 I__680 (
            .O(N__4652),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0 ));
    CascadeMux I__679 (
            .O(N__4649),
            .I(N__4645));
    CascadeMux I__678 (
            .O(N__4648),
            .I(N__4641));
    InMux I__677 (
            .O(N__4645),
            .I(N__4638));
    InMux I__676 (
            .O(N__4644),
            .I(N__4635));
    InMux I__675 (
            .O(N__4641),
            .I(N__4632));
    LocalMux I__674 (
            .O(N__4638),
            .I(N__4629));
    LocalMux I__673 (
            .O(N__4635),
            .I(N__4624));
    LocalMux I__672 (
            .O(N__4632),
            .I(N__4624));
    Sp12to4 I__671 (
            .O(N__4629),
            .I(N__4621));
    Span12Mux_h I__670 (
            .O(N__4624),
            .I(N__4618));
    Span12Mux_v I__669 (
            .O(N__4621),
            .I(N__4615));
    Span12Mux_v I__668 (
            .O(N__4618),
            .I(N__4612));
    Odrv12 I__667 (
            .O(N__4615),
            .I(SIZ_c_0));
    Odrv12 I__666 (
            .O(N__4612),
            .I(SIZ_c_0));
    InMux I__665 (
            .O(N__4607),
            .I(N__4604));
    LocalMux I__664 (
            .O(N__4604),
            .I(N__4601));
    Odrv4 I__663 (
            .O(N__4601),
            .I(TACK_EN_i_ess));
    IoInMux I__662 (
            .O(N__4598),
            .I(N__4595));
    LocalMux I__661 (
            .O(N__4595),
            .I(N__4592));
    Span4Mux_s0_h I__660 (
            .O(N__4592),
            .I(N__4589));
    Sp12to4 I__659 (
            .O(N__4589),
            .I(N__4586));
    Span12Mux_v I__658 (
            .O(N__4586),
            .I(N__4583));
    Span12Mux_h I__657 (
            .O(N__4583),
            .I(N__4580));
    Odrv12 I__656 (
            .O(N__4580),
            .I(N_614_i));
    InMux I__655 (
            .O(N__4577),
            .I(N__4574));
    LocalMux I__654 (
            .O(N__4574),
            .I(\U712_CHIP_RAM.N_36 ));
    IoInMux I__653 (
            .O(N__4571),
            .I(N__4568));
    LocalMux I__652 (
            .O(N__4568),
            .I(N__4565));
    Span4Mux_s3_h I__651 (
            .O(N__4565),
            .I(N__4562));
    Span4Mux_v I__650 (
            .O(N__4562),
            .I(N__4559));
    Span4Mux_v I__649 (
            .O(N__4559),
            .I(N__4556));
    Span4Mux_h I__648 (
            .O(N__4556),
            .I(N__4553));
    Sp12to4 I__647 (
            .O(N__4553),
            .I(N__4550));
    Odrv12 I__646 (
            .O(N__4550),
            .I(CMA_c_4));
    InMux I__645 (
            .O(N__4547),
            .I(N__4544));
    LocalMux I__644 (
            .O(N__4544),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__643 (
            .O(N__4541),
            .I(N__4537));
    InMux I__642 (
            .O(N__4540),
            .I(N__4534));
    LocalMux I__641 (
            .O(N__4537),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__640 (
            .O(N__4534),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    InMux I__639 (
            .O(N__4529),
            .I(N__4526));
    LocalMux I__638 (
            .O(N__4526),
            .I(\U712_REG_SM.N_188 ));
    InMux I__637 (
            .O(N__4523),
            .I(N__4519));
    InMux I__636 (
            .O(N__4522),
            .I(N__4516));
    LocalMux I__635 (
            .O(N__4519),
            .I(N__4511));
    LocalMux I__634 (
            .O(N__4516),
            .I(N__4511));
    Odrv4 I__633 (
            .O(N__4511),
            .I(REG_TACK));
    CascadeMux I__632 (
            .O(N__4508),
            .I(\U712_CYCLE_TERM.TACK_EN6_0_cascade_ ));
    CascadeMux I__631 (
            .O(N__4505),
            .I(\U712_CYCLE_TERM.N_45_0_0_en_cascade_ ));
    InMux I__630 (
            .O(N__4502),
            .I(N__4499));
    LocalMux I__629 (
            .O(N__4499),
            .I(N__4495));
    InMux I__628 (
            .O(N__4498),
            .I(N__4492));
    Span4Mux_v I__627 (
            .O(N__4495),
            .I(N__4487));
    LocalMux I__626 (
            .O(N__4492),
            .I(N__4487));
    Span4Mux_v I__625 (
            .O(N__4487),
            .I(N__4484));
    Sp12to4 I__624 (
            .O(N__4484),
            .I(N__4481));
    Span12Mux_h I__623 (
            .O(N__4481),
            .I(N__4478));
    Odrv12 I__622 (
            .O(N__4478),
            .I(REGSPACEn_c));
    InMux I__621 (
            .O(N__4475),
            .I(N__4471));
    InMux I__620 (
            .O(N__4474),
            .I(N__4468));
    LocalMux I__619 (
            .O(N__4471),
            .I(N__4464));
    LocalMux I__618 (
            .O(N__4468),
            .I(N__4461));
    InMux I__617 (
            .O(N__4467),
            .I(N__4458));
    Odrv4 I__616 (
            .O(N__4464),
            .I(\U712_REG_SM.DS_EN_0_sqmuxa_1 ));
    Odrv4 I__615 (
            .O(N__4461),
            .I(\U712_REG_SM.DS_EN_0_sqmuxa_1 ));
    LocalMux I__614 (
            .O(N__4458),
            .I(\U712_REG_SM.DS_EN_0_sqmuxa_1 ));
    CascadeMux I__613 (
            .O(N__4451),
            .I(N__4446));
    InMux I__612 (
            .O(N__4450),
            .I(N__4443));
    CascadeMux I__611 (
            .O(N__4449),
            .I(N__4440));
    InMux I__610 (
            .O(N__4446),
            .I(N__4437));
    LocalMux I__609 (
            .O(N__4443),
            .I(N__4434));
    InMux I__608 (
            .O(N__4440),
            .I(N__4431));
    LocalMux I__607 (
            .O(N__4437),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    Odrv4 I__606 (
            .O(N__4434),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    LocalMux I__605 (
            .O(N__4431),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    InMux I__604 (
            .O(N__4424),
            .I(N__4420));
    InMux I__603 (
            .O(N__4423),
            .I(N__4417));
    LocalMux I__602 (
            .O(N__4420),
            .I(CPU_TACKm));
    LocalMux I__601 (
            .O(N__4417),
            .I(CPU_TACKm));
    CascadeMux I__600 (
            .O(N__4412),
            .I(N__4406));
    InMux I__599 (
            .O(N__4411),
            .I(N__4403));
    InMux I__598 (
            .O(N__4410),
            .I(N__4400));
    InMux I__597 (
            .O(N__4409),
            .I(N__4395));
    InMux I__596 (
            .O(N__4406),
            .I(N__4395));
    LocalMux I__595 (
            .O(N__4403),
            .I(N__4392));
    LocalMux I__594 (
            .O(N__4400),
            .I(N__4389));
    LocalMux I__593 (
            .O(N__4395),
            .I(N__4386));
    Span4Mux_v I__592 (
            .O(N__4392),
            .I(N__4383));
    Span4Mux_v I__591 (
            .O(N__4389),
            .I(N__4378));
    Span4Mux_v I__590 (
            .O(N__4386),
            .I(N__4378));
    Sp12to4 I__589 (
            .O(N__4383),
            .I(N__4375));
    Span4Mux_h I__588 (
            .O(N__4378),
            .I(N__4372));
    Span12Mux_h I__587 (
            .O(N__4375),
            .I(N__4367));
    Sp12to4 I__586 (
            .O(N__4372),
            .I(N__4367));
    Span12Mux_v I__585 (
            .O(N__4367),
            .I(N__4364));
    Odrv12 I__584 (
            .O(N__4364),
            .I(CLK40_OUT_i));
    InMux I__583 (
            .O(N__4361),
            .I(N__4355));
    InMux I__582 (
            .O(N__4360),
            .I(N__4355));
    LocalMux I__581 (
            .O(N__4355),
            .I(N__4350));
    InMux I__580 (
            .O(N__4354),
            .I(N__4345));
    InMux I__579 (
            .O(N__4353),
            .I(N__4345));
    Odrv4 I__578 (
            .O(N__4350),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__577 (
            .O(N__4345),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    CascadeMux I__576 (
            .O(N__4340),
            .I(N__4337));
    InMux I__575 (
            .O(N__4337),
            .I(N__4333));
    InMux I__574 (
            .O(N__4336),
            .I(N__4330));
    LocalMux I__573 (
            .O(N__4333),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    LocalMux I__572 (
            .O(N__4330),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    InMux I__571 (
            .O(N__4325),
            .I(N__4322));
    LocalMux I__570 (
            .O(N__4322),
            .I(N__4319));
    Odrv4 I__569 (
            .O(N__4319),
            .I(\U712_REG_SM.UDS_OUT_2_0_0 ));
    InMux I__568 (
            .O(N__4316),
            .I(N__4312));
    InMux I__567 (
            .O(N__4315),
            .I(N__4309));
    LocalMux I__566 (
            .O(N__4312),
            .I(\U712_REG_SM.LDS_OUTZ0 ));
    LocalMux I__565 (
            .O(N__4309),
            .I(\U712_REG_SM.LDS_OUTZ0 ));
    IoInMux I__564 (
            .O(N__4304),
            .I(N__4301));
    LocalMux I__563 (
            .O(N__4301),
            .I(N__4298));
    IoSpan4Mux I__562 (
            .O(N__4298),
            .I(N__4295));
    IoSpan4Mux I__561 (
            .O(N__4295),
            .I(N__4292));
    Span4Mux_s2_v I__560 (
            .O(N__4292),
            .I(N__4289));
    Sp12to4 I__559 (
            .O(N__4289),
            .I(N__4286));
    Span12Mux_v I__558 (
            .O(N__4286),
            .I(N__4283));
    Odrv12 I__557 (
            .O(N__4283),
            .I(U712_REG_SM_un1_LDSn_i));
    InMux I__556 (
            .O(N__4280),
            .I(N__4277));
    LocalMux I__555 (
            .O(N__4277),
            .I(N__4273));
    InMux I__554 (
            .O(N__4276),
            .I(N__4270));
    Odrv4 I__553 (
            .O(N__4273),
            .I(\U712_REG_SM.UDS_OUTZ0 ));
    LocalMux I__552 (
            .O(N__4270),
            .I(\U712_REG_SM.UDS_OUTZ0 ));
    InMux I__551 (
            .O(N__4265),
            .I(N__4261));
    InMux I__550 (
            .O(N__4264),
            .I(N__4258));
    LocalMux I__549 (
            .O(N__4261),
            .I(N__4252));
    LocalMux I__548 (
            .O(N__4258),
            .I(N__4252));
    InMux I__547 (
            .O(N__4257),
            .I(N__4249));
    Odrv12 I__546 (
            .O(N__4252),
            .I(\U712_REG_SM.DS_ENZ0 ));
    LocalMux I__545 (
            .O(N__4249),
            .I(\U712_REG_SM.DS_ENZ0 ));
    IoInMux I__544 (
            .O(N__4244),
            .I(N__4241));
    LocalMux I__543 (
            .O(N__4241),
            .I(N__4238));
    IoSpan4Mux I__542 (
            .O(N__4238),
            .I(N__4235));
    IoSpan4Mux I__541 (
            .O(N__4235),
            .I(N__4232));
    Sp12to4 I__540 (
            .O(N__4232),
            .I(N__4229));
    Span12Mux_v I__539 (
            .O(N__4229),
            .I(N__4226));
    Odrv12 I__538 (
            .O(N__4226),
            .I(U712_REG_SM_un1_UDSn_i));
    InMux I__537 (
            .O(N__4223),
            .I(N__4220));
    LocalMux I__536 (
            .O(N__4220),
            .I(N__4217));
    Span4Mux_v I__535 (
            .O(N__4217),
            .I(N__4214));
    Sp12to4 I__534 (
            .O(N__4214),
            .I(N__4211));
    Odrv12 I__533 (
            .O(N__4211),
            .I(A_c_13));
    CascadeMux I__532 (
            .O(N__4208),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_4_cascade_ ));
    InMux I__531 (
            .O(N__4205),
            .I(N__4202));
    LocalMux I__530 (
            .O(N__4202),
            .I(N__4199));
    Span4Mux_h I__529 (
            .O(N__4199),
            .I(N__4196));
    Sp12to4 I__528 (
            .O(N__4196),
            .I(N__4193));
    Span12Mux_v I__527 (
            .O(N__4193),
            .I(N__4190));
    Odrv12 I__526 (
            .O(N__4190),
            .I(A_c_6));
    InMux I__525 (
            .O(N__4187),
            .I(N__4184));
    LocalMux I__524 (
            .O(N__4184),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    CascadeMux I__523 (
            .O(N__4181),
            .I(N__4175));
    InMux I__522 (
            .O(N__4180),
            .I(N__4172));
    InMux I__521 (
            .O(N__4179),
            .I(N__4169));
    InMux I__520 (
            .O(N__4178),
            .I(N__4166));
    InMux I__519 (
            .O(N__4175),
            .I(N__4163));
    LocalMux I__518 (
            .O(N__4172),
            .I(N__4160));
    LocalMux I__517 (
            .O(N__4169),
            .I(\U712_REG_SM.N_163_0 ));
    LocalMux I__516 (
            .O(N__4166),
            .I(\U712_REG_SM.N_163_0 ));
    LocalMux I__515 (
            .O(N__4163),
            .I(\U712_REG_SM.N_163_0 ));
    Odrv4 I__514 (
            .O(N__4160),
            .I(\U712_REG_SM.N_163_0 ));
    CascadeMux I__513 (
            .O(N__4151),
            .I(N__4147));
    InMux I__512 (
            .O(N__4150),
            .I(N__4144));
    InMux I__511 (
            .O(N__4147),
            .I(N__4141));
    LocalMux I__510 (
            .O(N__4144),
            .I(N__4135));
    LocalMux I__509 (
            .O(N__4141),
            .I(N__4129));
    InMux I__508 (
            .O(N__4140),
            .I(N__4126));
    InMux I__507 (
            .O(N__4139),
            .I(N__4121));
    InMux I__506 (
            .O(N__4138),
            .I(N__4121));
    Span4Mux_h I__505 (
            .O(N__4135),
            .I(N__4118));
    InMux I__504 (
            .O(N__4134),
            .I(N__4111));
    InMux I__503 (
            .O(N__4133),
            .I(N__4111));
    InMux I__502 (
            .O(N__4132),
            .I(N__4111));
    Odrv4 I__501 (
            .O(N__4129),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__500 (
            .O(N__4126),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__499 (
            .O(N__4121),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    Odrv4 I__498 (
            .O(N__4118),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__497 (
            .O(N__4111),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    InMux I__496 (
            .O(N__4100),
            .I(N__4097));
    LocalMux I__495 (
            .O(N__4097),
            .I(\U712_REG_SM.N_186 ));
    CascadeMux I__494 (
            .O(N__4094),
            .I(\U712_REG_SM.N_176_0_cascade_ ));
    InMux I__493 (
            .O(N__4091),
            .I(N__4085));
    InMux I__492 (
            .O(N__4090),
            .I(N__4080));
    InMux I__491 (
            .O(N__4089),
            .I(N__4080));
    InMux I__490 (
            .O(N__4088),
            .I(N__4077));
    LocalMux I__489 (
            .O(N__4085),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__488 (
            .O(N__4080),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__487 (
            .O(N__4077),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    InMux I__486 (
            .O(N__4070),
            .I(N__4063));
    InMux I__485 (
            .O(N__4069),
            .I(N__4063));
    InMux I__484 (
            .O(N__4068),
            .I(N__4060));
    LocalMux I__483 (
            .O(N__4063),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    LocalMux I__482 (
            .O(N__4060),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    CascadeMux I__481 (
            .O(N__4055),
            .I(N__4052));
    InMux I__480 (
            .O(N__4052),
            .I(N__4049));
    LocalMux I__479 (
            .O(N__4049),
            .I(N__4045));
    InMux I__478 (
            .O(N__4048),
            .I(N__4042));
    Odrv4 I__477 (
            .O(N__4045),
            .I(\U712_REG_SM.N_157_0 ));
    LocalMux I__476 (
            .O(N__4042),
            .I(\U712_REG_SM.N_157_0 ));
    InMux I__475 (
            .O(N__4037),
            .I(N__4029));
    InMux I__474 (
            .O(N__4036),
            .I(N__4024));
    InMux I__473 (
            .O(N__4035),
            .I(N__4024));
    CascadeMux I__472 (
            .O(N__4034),
            .I(N__4021));
    InMux I__471 (
            .O(N__4033),
            .I(N__4017));
    InMux I__470 (
            .O(N__4032),
            .I(N__4014));
    LocalMux I__469 (
            .O(N__4029),
            .I(N__4009));
    LocalMux I__468 (
            .O(N__4024),
            .I(N__4009));
    InMux I__467 (
            .O(N__4021),
            .I(N__4006));
    InMux I__466 (
            .O(N__4020),
            .I(N__4003));
    LocalMux I__465 (
            .O(N__4017),
            .I(N__4000));
    LocalMux I__464 (
            .O(N__4014),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    Odrv4 I__463 (
            .O(N__4009),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__462 (
            .O(N__4006),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__461 (
            .O(N__4003),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    Odrv4 I__460 (
            .O(N__4000),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    CascadeMux I__459 (
            .O(N__3989),
            .I(N__3982));
    InMux I__458 (
            .O(N__3988),
            .I(N__3979));
    InMux I__457 (
            .O(N__3987),
            .I(N__3976));
    InMux I__456 (
            .O(N__3986),
            .I(N__3973));
    InMux I__455 (
            .O(N__3985),
            .I(N__3968));
    InMux I__454 (
            .O(N__3982),
            .I(N__3968));
    LocalMux I__453 (
            .O(N__3979),
            .I(\U712_REG_SM.C1_SYNCZ0Z_2 ));
    LocalMux I__452 (
            .O(N__3976),
            .I(\U712_REG_SM.C1_SYNCZ0Z_2 ));
    LocalMux I__451 (
            .O(N__3973),
            .I(\U712_REG_SM.C1_SYNCZ0Z_2 ));
    LocalMux I__450 (
            .O(N__3968),
            .I(\U712_REG_SM.C1_SYNCZ0Z_2 ));
    CascadeMux I__449 (
            .O(N__3959),
            .I(\U712_REG_SM.N_157_0_cascade_ ));
    CascadeMux I__448 (
            .O(N__3956),
            .I(N__3953));
    InMux I__447 (
            .O(N__3953),
            .I(N__3945));
    InMux I__446 (
            .O(N__3952),
            .I(N__3942));
    InMux I__445 (
            .O(N__3951),
            .I(N__3939));
    InMux I__444 (
            .O(N__3950),
            .I(N__3932));
    InMux I__443 (
            .O(N__3949),
            .I(N__3932));
    InMux I__442 (
            .O(N__3948),
            .I(N__3932));
    LocalMux I__441 (
            .O(N__3945),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__440 (
            .O(N__3942),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__439 (
            .O(N__3939),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__438 (
            .O(N__3932),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    InMux I__437 (
            .O(N__3923),
            .I(N__3920));
    LocalMux I__436 (
            .O(N__3920),
            .I(\U712_REG_SM.N_176_0 ));
    CascadeMux I__435 (
            .O(N__3917),
            .I(N__3912));
    CascadeMux I__434 (
            .O(N__3916),
            .I(N__3909));
    InMux I__433 (
            .O(N__3915),
            .I(N__3906));
    InMux I__432 (
            .O(N__3912),
            .I(N__3901));
    InMux I__431 (
            .O(N__3909),
            .I(N__3901));
    LocalMux I__430 (
            .O(N__3906),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__429 (
            .O(N__3901),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    InMux I__428 (
            .O(N__3896),
            .I(N__3893));
    LocalMux I__427 (
            .O(N__3893),
            .I(N__3887));
    InMux I__426 (
            .O(N__3892),
            .I(N__3880));
    InMux I__425 (
            .O(N__3891),
            .I(N__3880));
    InMux I__424 (
            .O(N__3890),
            .I(N__3880));
    Odrv4 I__423 (
            .O(N__3887),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    LocalMux I__422 (
            .O(N__3880),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    CascadeMux I__421 (
            .O(N__3875),
            .I(N__3871));
    CascadeMux I__420 (
            .O(N__3874),
            .I(N__3868));
    InMux I__419 (
            .O(N__3871),
            .I(N__3865));
    InMux I__418 (
            .O(N__3868),
            .I(N__3861));
    LocalMux I__417 (
            .O(N__3865),
            .I(N__3858));
    InMux I__416 (
            .O(N__3864),
            .I(N__3855));
    LocalMux I__415 (
            .O(N__3861),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    Odrv4 I__414 (
            .O(N__3858),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__413 (
            .O(N__3855),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    InMux I__412 (
            .O(N__3848),
            .I(N__3845));
    LocalMux I__411 (
            .O(N__3845),
            .I(\U712_REG_SM.N_192 ));
    IoInMux I__410 (
            .O(N__3842),
            .I(N__3839));
    LocalMux I__409 (
            .O(N__3839),
            .I(N__3836));
    Span4Mux_s0_h I__408 (
            .O(N__3836),
            .I(N__3833));
    Span4Mux_h I__407 (
            .O(N__3833),
            .I(N__3830));
    Sp12to4 I__406 (
            .O(N__3830),
            .I(N__3827));
    Span12Mux_v I__405 (
            .O(N__3827),
            .I(N__3823));
    InMux I__404 (
            .O(N__3826),
            .I(N__3820));
    Odrv12 I__403 (
            .O(N__3823),
            .I(TACK_OUTn));
    LocalMux I__402 (
            .O(N__3820),
            .I(TACK_OUTn));
    InMux I__401 (
            .O(N__3815),
            .I(N__3811));
    InMux I__400 (
            .O(N__3814),
            .I(N__3807));
    LocalMux I__399 (
            .O(N__3811),
            .I(N__3803));
    InMux I__398 (
            .O(N__3810),
            .I(N__3800));
    LocalMux I__397 (
            .O(N__3807),
            .I(N__3797));
    InMux I__396 (
            .O(N__3806),
            .I(N__3794));
    Odrv12 I__395 (
            .O(N__3803),
            .I(\U712_REG_SM.N_171_0 ));
    LocalMux I__394 (
            .O(N__3800),
            .I(\U712_REG_SM.N_171_0 ));
    Odrv4 I__393 (
            .O(N__3797),
            .I(\U712_REG_SM.N_171_0 ));
    LocalMux I__392 (
            .O(N__3794),
            .I(\U712_REG_SM.N_171_0 ));
    IoInMux I__391 (
            .O(N__3785),
            .I(N__3782));
    LocalMux I__390 (
            .O(N__3782),
            .I(N__3779));
    Span12Mux_s4_v I__389 (
            .O(N__3779),
            .I(N__3776));
    Odrv12 I__388 (
            .O(N__3776),
            .I(VBENn_c));
    InMux I__387 (
            .O(N__3773),
            .I(N__3770));
    LocalMux I__386 (
            .O(N__3770),
            .I(N__3766));
    InMux I__385 (
            .O(N__3769),
            .I(N__3763));
    Odrv4 I__384 (
            .O(N__3766),
            .I(\U712_REG_SM.N_162_0 ));
    LocalMux I__383 (
            .O(N__3763),
            .I(\U712_REG_SM.N_162_0 ));
    CascadeMux I__382 (
            .O(N__3758),
            .I(\U712_REG_SM.N_171_0_cascade_ ));
    InMux I__381 (
            .O(N__3755),
            .I(N__3752));
    LocalMux I__380 (
            .O(N__3752),
            .I(\U712_REG_SM.RnW_m ));
    CascadeMux I__379 (
            .O(N__3749),
            .I(\U712_REG_SM.un1_LDS_OUT_0_sqmuxa_1_0_cascade_ ));
    CascadeMux I__378 (
            .O(N__3746),
            .I(N__3742));
    InMux I__377 (
            .O(N__3745),
            .I(N__3738));
    InMux I__376 (
            .O(N__3742),
            .I(N__3735));
    InMux I__375 (
            .O(N__3741),
            .I(N__3732));
    LocalMux I__374 (
            .O(N__3738),
            .I(\U712_REG_SM.N_165_0 ));
    LocalMux I__373 (
            .O(N__3735),
            .I(\U712_REG_SM.N_165_0 ));
    LocalMux I__372 (
            .O(N__3732),
            .I(\U712_REG_SM.N_165_0 ));
    CascadeMux I__371 (
            .O(N__3725),
            .I(\U712_REG_SM.N_167_0_cascade_ ));
    InMux I__370 (
            .O(N__3722),
            .I(N__3713));
    InMux I__369 (
            .O(N__3721),
            .I(N__3713));
    InMux I__368 (
            .O(N__3720),
            .I(N__3713));
    LocalMux I__367 (
            .O(N__3713),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    InMux I__366 (
            .O(N__3710),
            .I(N__3704));
    InMux I__365 (
            .O(N__3709),
            .I(N__3704));
    LocalMux I__364 (
            .O(N__3704),
            .I(\U712_REG_SM.N_167_0 ));
    InMux I__363 (
            .O(N__3701),
            .I(N__3696));
    InMux I__362 (
            .O(N__3700),
            .I(N__3693));
    InMux I__361 (
            .O(N__3699),
            .I(N__3690));
    LocalMux I__360 (
            .O(N__3696),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    LocalMux I__359 (
            .O(N__3693),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    LocalMux I__358 (
            .O(N__3690),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    CascadeMux I__357 (
            .O(N__3683),
            .I(\U712_REG_SM.DS_EN_0_sqmuxa_1_0_a3_0_cascade_ ));
    InMux I__356 (
            .O(N__3680),
            .I(N__3677));
    LocalMux I__355 (
            .O(N__3677),
            .I(N__3673));
    IoInMux I__354 (
            .O(N__3676),
            .I(N__3670));
    Span4Mux_v I__353 (
            .O(N__3673),
            .I(N__3667));
    LocalMux I__352 (
            .O(N__3670),
            .I(N__3664));
    Sp12to4 I__351 (
            .O(N__3667),
            .I(N__3661));
    Span4Mux_s3_h I__350 (
            .O(N__3664),
            .I(N__3658));
    Span12Mux_h I__349 (
            .O(N__3661),
            .I(N__3653));
    Sp12to4 I__348 (
            .O(N__3658),
            .I(N__3653));
    Span12Mux_v I__347 (
            .O(N__3653),
            .I(N__3650));
    Odrv12 I__346 (
            .O(N__3650),
            .I(C1_c));
    CascadeMux I__345 (
            .O(N__3647),
            .I(\U712_REG_SM.N_162_0_cascade_ ));
    InMux I__344 (
            .O(N__3644),
            .I(N__3641));
    LocalMux I__343 (
            .O(N__3641),
            .I(N__3636));
    InMux I__342 (
            .O(N__3640),
            .I(N__3631));
    InMux I__341 (
            .O(N__3639),
            .I(N__3631));
    Odrv4 I__340 (
            .O(N__3636),
            .I(\U712_REG_SM.N_166_0 ));
    LocalMux I__339 (
            .O(N__3631),
            .I(\U712_REG_SM.N_166_0 ));
    InMux I__338 (
            .O(N__3626),
            .I(N__3623));
    LocalMux I__337 (
            .O(N__3623),
            .I(N__3620));
    Span12Mux_h I__336 (
            .O(N__3620),
            .I(N__3617));
    Span12Mux_v I__335 (
            .O(N__3617),
            .I(N__3614));
    Odrv12 I__334 (
            .O(N__3614),
            .I(C3_c));
    CascadeMux I__333 (
            .O(N__3611),
            .I(\U712_REG_SM.REG_TACK_7_0_cascade_ ));
    InMux I__332 (
            .O(N__3608),
            .I(N__3604));
    InMux I__331 (
            .O(N__3607),
            .I(N__3601));
    LocalMux I__330 (
            .O(N__3604),
            .I(\U712_REG_SM.un1_STATE_COUNT_5_0_1 ));
    LocalMux I__329 (
            .O(N__3601),
            .I(\U712_REG_SM.un1_STATE_COUNT_5_0_1 ));
    CascadeMux I__328 (
            .O(N__3596),
            .I(\U712_REG_SM.N_183_cascade_ ));
    IoInMux I__327 (
            .O(N__3593),
            .I(N__3590));
    LocalMux I__326 (
            .O(N__3590),
            .I(N__3587));
    Odrv12 I__325 (
            .O(N__3587),
            .I(CLK40_OUT_i_i));
    IoInMux I__324 (
            .O(N__3584),
            .I(N__3581));
    LocalMux I__323 (
            .O(N__3581),
            .I(N__3578));
    Span4Mux_s2_v I__322 (
            .O(N__3578),
            .I(N__3575));
    Span4Mux_v I__321 (
            .O(N__3575),
            .I(N__3572));
    Span4Mux_h I__320 (
            .O(N__3572),
            .I(N__3569));
    Odrv4 I__319 (
            .O(N__3569),
            .I(CLK80_OUT_i_i));
    IoInMux I__318 (
            .O(N__3566),
            .I(N__3563));
    LocalMux I__317 (
            .O(N__3563),
            .I(N__3559));
    IoInMux I__316 (
            .O(N__3562),
            .I(N__3556));
    IoSpan4Mux I__315 (
            .O(N__3559),
            .I(N__3553));
    LocalMux I__314 (
            .O(N__3556),
            .I(N__3550));
    Sp12to4 I__313 (
            .O(N__3553),
            .I(N__3547));
    IoSpan4Mux I__312 (
            .O(N__3550),
            .I(N__3544));
    Span12Mux_s6_v I__311 (
            .O(N__3547),
            .I(N__3541));
    Sp12to4 I__310 (
            .O(N__3544),
            .I(N__3538));
    Span12Mux_v I__309 (
            .O(N__3541),
            .I(N__3535));
    Span12Mux_s6_v I__308 (
            .O(N__3538),
            .I(N__3532));
    Span12Mux_h I__307 (
            .O(N__3535),
            .I(N__3526));
    Span12Mux_v I__306 (
            .O(N__3532),
            .I(N__3526));
    InMux I__305 (
            .O(N__3531),
            .I(N__3523));
    Odrv12 I__304 (
            .O(N__3526),
            .I(ASn_c));
    LocalMux I__303 (
            .O(N__3523),
            .I(ASn_c));
    IoInMux I__302 (
            .O(N__3518),
            .I(N__3515));
    LocalMux I__301 (
            .O(N__3515),
            .I(N__3512));
    IoSpan4Mux I__300 (
            .O(N__3512),
            .I(N__3509));
    Span4Mux_s2_v I__299 (
            .O(N__3509),
            .I(N__3506));
    Sp12to4 I__298 (
            .O(N__3506),
            .I(N__3503));
    Span12Mux_v I__297 (
            .O(N__3503),
            .I(N__3500));
    Odrv12 I__296 (
            .O(N__3500),
            .I(CLK40_IN_c));
    defparam IN_MUX_bfv_10_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_7_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__6554),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__3676),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CLK40C_obuf_RNO_LC_3_10_4.C_ON=1'b0;
    defparam CLK40C_obuf_RNO_LC_3_10_4.SEQ_MODE=4'b0000;
    defparam CLK40C_obuf_RNO_LC_3_10_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLK40C_obuf_RNO_LC_3_10_4 (
            .in0(N__4411),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_OUT_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_5_1_2.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_5_1_2.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_5_1_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLKRAM_obuf_RNO_LC_5_1_2 (
            .in0(N__9287),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK80_OUT_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REGENn_1_LC_7_8_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_1_LC_7_8_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_1_LC_7_8_1 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \U712_REG_SM.REGENn_1_LC_7_8_1  (
            .in0(N__3810),
            .in1(N__3531),
            .in2(_gnd_net_),
            .in3(N__4474),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9270),
            .ce(),
            .sr(N__9064));
    defparam \U712_REG_SM.STATE_COUNT_5_LC_7_8_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_7_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_7_8_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_REG_SM.STATE_COUNT_5_LC_7_8_5  (
            .in0(_gnd_net_),
            .in1(N__3607),
            .in2(_gnd_net_),
            .in3(N__3644),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9270),
            .ce(),
            .sr(N__9064));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_7_9_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_7_9_0 .LUT_INIT=16'b0001110100111111;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_7_9_0  (
            .in0(N__3891),
            .in1(N__6746),
            .in2(N__3917),
            .in3(N__3639),
            .lcout(),
            .ltout(\U712_REG_SM.REG_TACK_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_LC_7_9_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_7_9_1 .LUT_INIT=16'b0010111000001111;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_7_9_1  (
            .in0(N__4523),
            .in1(N__3701),
            .in2(N__3611),
            .in3(N__3608),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9274),
            .ce(),
            .sr(N__9058));
    defparam \U712_REG_SM.STATE_COUNT_RNIFFKI2_4_LC_7_9_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIFFKI2_4_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIFFKI2_4_LC_7_9_2 .LUT_INIT=16'b0100010101010101;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIFFKI2_4_LC_7_9_2  (
            .in0(N__3890),
            .in1(N__4139),
            .in2(N__3916),
            .in3(N__4178),
            .lcout(\U712_REG_SM.un1_STATE_COUNT_5_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_7_9_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_7_9_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_7_9_3  (
            .in0(N__4037),
            .in1(N__3745),
            .in2(N__3956),
            .in3(N__3988),
            .lcout(),
            .ltout(\U712_REG_SM.N_183_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_6_LC_7_9_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_7_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_7_9_4 .LUT_INIT=16'b0000111000001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_6_LC_7_9_4  (
            .in0(N__3892),
            .in1(N__3700),
            .in2(N__3596),
            .in3(N__3640),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9274),
            .ce(),
            .sr(N__9058));
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_7_9_6 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_7_9_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_0_LC_7_9_6  (
            .in0(_gnd_net_),
            .in1(N__6745),
            .in2(_gnd_net_),
            .in3(N__4138),
            .lcout(\U712_REG_SM.RnW_m ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIQU741_2_LC_7_10_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIQU741_2_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIQU741_2_LC_7_10_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIQU741_2_LC_7_10_0  (
            .in0(N__4089),
            .in1(N__4069),
            .in2(_gnd_net_),
            .in3(N__4133),
            .lcout(\U712_REG_SM.N_165_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_1_LC_7_10_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_7_10_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_7_10_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_7_10_1  (
            .in0(N__4134),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9278),
            .ce(),
            .sr(N__9051));
    defparam \U712_REG_SM.C1_SYNC_2_LC_7_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_2_LC_7_10_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_2_LC_7_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_2_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3950),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9278),
            .ce(),
            .sr(N__9051));
    defparam \U712_REG_SM.STATE_COUNT_RNI81E81_6_LC_7_10_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI81E81_6_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI81E81_6_LC_7_10_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI81E81_6_LC_7_10_3  (
            .in0(N__3949),
            .in1(N__3699),
            .in2(N__4034),
            .in3(N__3985),
            .lcout(),
            .ltout(\U712_REG_SM.DS_EN_0_sqmuxa_1_0_a3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_7_10_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_7_10_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_7_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3683),
            .in3(N__3741),
            .lcout(\U712_REG_SM.DS_EN_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_0_LC_7_10_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_7_10_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_7_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_7_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3680),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9278),
            .ce(),
            .sr(N__9051));
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_7_10_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_7_10_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_7_10_6  (
            .in0(N__4033),
            .in1(N__4132),
            .in2(N__3989),
            .in3(N__3948),
            .lcout(\U712_REG_SM.N_162_0 ),
            .ltout(\U712_REG_SM.N_162_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_7_10_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_7_10_7 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_7_10_7  (
            .in0(N__4070),
            .in1(_gnd_net_),
            .in2(N__3647),
            .in3(N__4090),
            .lcout(\U712_REG_SM.N_166_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_2_LC_7_11_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_2_LC_7_11_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_2_LC_7_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_2_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4091),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9281),
            .ce(),
            .sr(N__9041));
    defparam \U712_REG_SM.C3_SYNC_0_LC_7_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_7_11_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_7_11_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_7_11_4  (
            .in0(N__3626),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9281),
            .ce(),
            .sr(N__9041));
    defparam \U712_REG_SM.C3_SYNC_1_LC_7_11_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_7_11_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_7_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4032),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9281),
            .ce(),
            .sr(N__9041));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_7_12_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_7_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_7_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4670),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9283),
            .ce(),
            .sr(N__9033));
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_6_5 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_6_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a2_LC_8_6_5  (
            .in0(N__7500),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8861),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_8_8_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_8_8_1 .LUT_INIT=16'b0101010100010101;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_8_8_1  (
            .in0(N__4529),
            .in1(N__3773),
            .in2(N__4055),
            .in3(N__4450),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9265),
            .ce(),
            .sr(N__9059));
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_8_9_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_8_9_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_8_9_0  (
            .in0(N__4540),
            .in1(N__3769),
            .in2(_gnd_net_),
            .in3(N__4048),
            .lcout(\U712_REG_SM.N_171_0 ),
            .ltout(\U712_REG_SM.N_171_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_8_9_1 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_8_9_1 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_1_LC_8_9_1  (
            .in0(N__3720),
            .in1(N__3709),
            .in2(N__3758),
            .in3(N__4467),
            .lcout(),
            .ltout(\U712_REG_SM.un1_LDS_OUT_0_sqmuxa_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_LC_8_9_2 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DS_EN_LC_8_9_2 .LUT_INIT=16'b1111111000001110;
    LogicCell40 \U712_REG_SM.DS_EN_LC_8_9_2  (
            .in0(N__3755),
            .in1(N__4036),
            .in2(N__3749),
            .in3(N__4257),
            .lcout(\U712_REG_SM.DS_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9271),
            .ce(),
            .sr(N__9052));
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_2_LC_8_9_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_2_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_2_LC_8_9_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNIIDN62_2_LC_8_9_3  (
            .in0(N__4035),
            .in1(N__3987),
            .in2(N__3746),
            .in3(N__3952),
            .lcout(\U712_REG_SM.N_167_0 ),
            .ltout(\U712_REG_SM.N_167_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_8_9_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_8_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_8_9_4 .LUT_INIT=16'b0000111100001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__3721),
            .in2(N__3725),
            .in3(N__3806),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9271),
            .ce(),
            .sr(N__9052));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_8_9_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_8_9_5 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_8_9_5  (
            .in0(N__3722),
            .in1(N__3710),
            .in2(N__3874),
            .in3(N__4100),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9271),
            .ce(),
            .sr(N__9052));
    defparam \U712_REG_SM.STATE_COUNT_RNIVAPS2_3_LC_8_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIVAPS2_3_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIVAPS2_3_LC_8_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIVAPS2_3_LC_8_10_2  (
            .in0(N__4871),
            .in1(N__4839),
            .in2(N__4181),
            .in3(N__3864),
            .lcout(\U712_REG_SM.N_176_0 ),
            .ltout(\U712_REG_SM.N_176_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_8_10_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_8_10_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_0_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4094),
            .in3(N__4140),
            .lcout(\U712_REG_SM.N_192 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_8_10_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_8_10_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_8_10_4  (
            .in0(N__4088),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4068),
            .lcout(\U712_REG_SM.N_157_0 ),
            .ltout(\U712_REG_SM.N_157_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI1FQR1_2_LC_8_10_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI1FQR1_2_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI1FQR1_2_LC_8_10_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI1FQR1_2_LC_8_10_5  (
            .in0(N__4020),
            .in1(N__3986),
            .in2(N__3959),
            .in3(N__3951),
            .lcout(\U712_REG_SM.N_163_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_8_10_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_8_10_7 .LUT_INIT=16'b1111010111000100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_8_10_7  (
            .in0(N__4179),
            .in1(N__3923),
            .in2(N__4151),
            .in3(N__3915),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9275),
            .ce(),
            .sr(N__9042));
    defparam \U712_REG_SM.REG_CYCLE_LC_8_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_8_11_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_8_11_1  (
            .in0(N__3896),
            .in1(N__7490),
            .in2(N__3875),
            .in3(N__3848),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9279),
            .ce(),
            .sr(N__9034));
    defparam \U712_REG_SM.UDS_OUT_LC_8_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.UDS_OUT_LC_8_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.UDS_OUT_LC_8_11_6 .LUT_INIT=16'b0101111111001100;
    LogicCell40 \U712_REG_SM.UDS_OUT_LC_8_11_6  (
            .in0(N__4325),
            .in1(N__4276),
            .in2(N__4649),
            .in3(N__3814),
            .lcout(\U712_REG_SM.UDS_OUTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9279),
            .ce(),
            .sr(N__9034));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_12_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_12_3 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_12_3 .LUT_INIT=16'b1111111111000100;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_8_12_3  (
            .in0(N__4361),
            .in1(N__3826),
            .in2(N__4412),
            .in3(N__4689),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9282),
            .ce(),
            .sr(N__9022));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_8_12_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_8_12_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(N__4409),
            .in2(_gnd_net_),
            .in3(N__4360),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9282),
            .ce(),
            .sr(N__9022));
    defparam \U712_REG_SM.LDS_OUT_LC_8_12_6 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.LDS_OUT_LC_8_12_6 .LUT_INIT=16'b0101111111001100;
    LogicCell40 \U712_REG_SM.LDS_OUT_LC_8_12_6  (
            .in0(N__4703),
            .in1(N__4315),
            .in2(N__4648),
            .in3(N__3815),
            .lcout(\U712_REG_SM.LDS_OUTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9282),
            .ce(),
            .sr(N__9022));
    defparam \U712_REG_SM.UDS_OUT_RNO_0_LC_8_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.UDS_OUT_RNO_0_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDS_OUT_RNO_0_LC_8_13_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_REG_SM.UDS_OUT_RNO_0_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__6736),
            .in2(_gnd_net_),
            .in3(N__5164),
            .lcout(\U712_REG_SM.UDS_OUT_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_8_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_8_13_7 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_REG_SM.LDS_OUT_RNIL31J_LC_8_13_7  (
            .in0(N__4264),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4316),
            .lcout(U712_REG_SM_un1_LDSn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_8_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_8_14_7 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_REG_SM.UDS_OUT_RNIUP9B_LC_8_14_7  (
            .in0(N__4280),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4265),
            .lcout(U712_REG_SM_un1_UDSn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_6_5 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_6_5  (
            .in0(N__4187),
            .in1(N__8856),
            .in2(N__8133),
            .in3(N__4547),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_9_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_9_6_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_9_6_6  (
            .in0(N__8857),
            .in1(N__4223),
            .in2(N__4208),
            .in3(N__4205),
            .lcout(\U712_CHIP_RAM.N_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_9_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_9_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_9_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7871),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9252),
            .ce(N__8285),
            .sr(N__9060));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_8_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_8_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_8_2  (
            .in0(N__4180),
            .in1(N__4870),
            .in2(N__4850),
            .in3(N__4150),
            .lcout(\U712_REG_SM.N_186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DBR_SYNC_1_LC_9_8_3 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_9_8_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_9_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.DBR_SYNC_1_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4849),
            .lcout(U712_REG_SM_DBR_SYNC_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9259),
            .ce(),
            .sr(N__9053));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_9_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_9_1 .LUT_INIT=16'b0000000011101111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_9_1  (
            .in0(N__4905),
            .in1(N__4498),
            .in2(N__4449),
            .in3(N__4541),
            .lcout(\U712_REG_SM.N_188 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_9_9_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_9_9_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN6_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__4522),
            .in2(_gnd_net_),
            .in3(N__4423),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(\U712_CYCLE_TERM.TACK_EN6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_9_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_9_5 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_9_5  (
            .in0(N__6625),
            .in1(N__4752),
            .in2(N__4508),
            .in3(N__4336),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_45_0_0_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_9_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_9_6 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_9_6  (
            .in0(N__9119),
            .in1(_gnd_net_),
            .in2(N__4505),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.N_45_0_0_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_9_10_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_9_10_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_9_10_0 .LUT_INIT=16'b0000000011111000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_9_10_0  (
            .in0(N__4658),
            .in1(N__4734),
            .in2(N__4340),
            .in3(N__4353),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9272),
            .ce(),
            .sr(N__9035));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_9_10_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_9_10_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_9_10_1 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_9_10_1  (
            .in0(N__4912),
            .in1(N__4502),
            .in2(N__4451),
            .in3(N__4475),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9272),
            .ce(),
            .sr(N__9035));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_9_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_9_10_2 .LUT_INIT=16'b0010111000100010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_9_10_2  (
            .in0(N__4424),
            .in1(N__5033),
            .in2(N__6221),
            .in3(N__8864),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9272),
            .ce(),
            .sr(N__9035));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_10_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_10_5 .LUT_INIT=16'b1010111010001100;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_9_10_5  (
            .in0(N__4354),
            .in1(N__4753),
            .in2(N__4736),
            .in3(N__4410),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9272),
            .ce(),
            .sr(N__9035));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_9_10_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_9_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_9_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4697),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9272),
            .ce(),
            .sr(N__9035));
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_9_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_9_10_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_9_10_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DBR_SYNC_0_LC_9_10_7  (
            .in0(N__4775),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(U712_REG_SM_DBR_SYNC_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9272),
            .ce(),
            .sr(N__9035));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_9_11_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_9_11_5 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_9_11_5 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_LC_9_11_5  (
            .in0(N__6587),
            .in1(N__4754),
            .in2(_gnd_net_),
            .in3(N__4735),
            .lcout(TACK_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9276),
            .ce(N__4715),
            .sr(N__9023));
    defparam \U712_REG_SM.LDS_OUT_RNO_0_LC_9_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_RNO_0_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDS_OUT_RNO_0_LC_9_12_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_REG_SM.LDS_OUT_RNO_0_LC_9_12_0  (
            .in0(N__5180),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6756),
            .lcout(\U712_REG_SM.LDS_OUT_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_9_12_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_9_12_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__4693),
            .in2(_gnd_net_),
            .in3(N__4669),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LW_TRANS_LC_9_12_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LW_TRANS_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LW_TRANS_LC_9_12_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \U712_BYTE_ENABLE.LW_TRANS_LC_9_12_4  (
            .in0(N__5203),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4644),
            .lcout(\U712_BYTE_ENABLE.LW_TRANS_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TACKn_obuft_RNO_LC_9_13_7.C_ON=1'b0;
    defparam TACKn_obuft_RNO_LC_9_13_7.SEQ_MODE=4'b0000;
    defparam TACKn_obuft_RNO_LC_9_13_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 TACKn_obuft_RNO_LC_9_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4607),
            .lcout(N_614_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_10_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_10_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_10_5_7 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_10_5_7  (
            .in0(N__8433),
            .in1(N__4577),
            .in2(_gnd_net_),
            .in3(N__8552),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9236),
            .ce(N__8646),
            .sr(N__9065));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_10_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_10_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_10_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_10_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7789),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9245),
            .ce(N__7961),
            .sr(N__9061));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_10_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_10_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_10_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_10_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8330),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9245),
            .ce(N__7961),
            .sr(N__9061));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_7_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_7_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_7_0  (
            .in0(_gnd_net_),
            .in1(N__4985),
            .in2(_gnd_net_),
            .in3(N__4808),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(bfn_10_7_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__4784),
            .ce(),
            .sr(N__5234));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_7_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_7_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_7_1  (
            .in0(_gnd_net_),
            .in1(N__5012),
            .in2(_gnd_net_),
            .in3(N__4805),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__4784),
            .ce(),
            .sr(N__5234));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_7_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_7_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_7_2  (
            .in0(_gnd_net_),
            .in1(N__5024),
            .in2(_gnd_net_),
            .in3(N__4802),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__4784),
            .ce(),
            .sr(N__5234));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_7_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_7_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_7_3  (
            .in0(_gnd_net_),
            .in1(N__5713),
            .in2(_gnd_net_),
            .in3(N__4799),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__4784),
            .ce(),
            .sr(N__5234));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_7_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_7_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_7_4  (
            .in0(_gnd_net_),
            .in1(N__4999),
            .in2(_gnd_net_),
            .in3(N__4796),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__4784),
            .ce(),
            .sr(N__5234));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_7_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_7_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_7_5  (
            .in0(_gnd_net_),
            .in1(N__4961),
            .in2(_gnd_net_),
            .in3(N__4793),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__4784),
            .ce(),
            .sr(N__5234));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_7_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_7_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_7_6  (
            .in0(_gnd_net_),
            .in1(N__4973),
            .in2(_gnd_net_),
            .in3(N__4790),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__4784),
            .ce(),
            .sr(N__5234));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_7_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_7_7  (
            .in0(_gnd_net_),
            .in1(N__5680),
            .in2(_gnd_net_),
            .in3(N__4787),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4784),
            .ce(),
            .sr(N__5234));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_8_0 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_8_0  (
            .in0(N__5966),
            .in1(N__5763),
            .in2(N__6635),
            .in3(N__5335),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_49_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_8_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_8_1  (
            .in0(N__5357),
            .in1(_gnd_net_),
            .in2(N__5027),
            .in3(N__6507),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9253),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_8_2 .LUT_INIT=16'b0001111101011111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_8_2  (
            .in0(N__5023),
            .in1(N__5011),
            .in2(N__5000),
            .in3(N__4984),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_8_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_8_3  (
            .in0(_gnd_net_),
            .in1(N__4972),
            .in2(_gnd_net_),
            .in3(N__4960),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_10_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_10_8_4 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_10_8_4  (
            .in0(N__5965),
            .in1(N__6058),
            .in2(_gnd_net_),
            .in3(N__6203),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISSMN4_3_LC_10_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISSMN4_3_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISSMN4_3_LC_10_8_5 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNISSMN4_3_LC_10_8_5  (
            .in0(N__6149),
            .in1(N__5467),
            .in2(N__4949),
            .in3(N__6275),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_0_2_LC_10_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_0_2_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_0_2_LC_10_8_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_0_2_LC_10_8_7  (
            .in0(N__6057),
            .in1(N__5964),
            .in2(_gnd_net_),
            .in3(N__6202),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_9_0 .LUT_INIT=16'b0000001110101011;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_9_0  (
            .in0(N__4820),
            .in1(N__4946),
            .in2(N__4919),
            .in3(N__8848),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9260),
            .ce(),
            .sr(N__9036));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_10_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_10_9_1 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_10_9_1  (
            .in0(N__4866),
            .in1(N__7133),
            .in2(N__4845),
            .in3(N__4819),
            .lcout(\U712_CHIP_RAM.N_57 ),
            .ltout(\U712_CHIP_RAM.N_57_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0V852_2_LC_10_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0V852_2_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0V852_2_LC_10_9_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI0V852_2_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4811),
            .in3(N__6199),
            .lcout(\U712_CHIP_RAM.N_58 ),
            .ltout(\U712_CHIP_RAM.N_58_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSC34_0_LC_10_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSC34_0_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSC34_0_LC_10_9_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSC34_0_LC_10_9_3  (
            .in0(N__5952),
            .in1(N__6044),
            .in2(N__5066),
            .in3(N__5466),
            .lcout(\U712_CHIP_RAM.N_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN7BL3_LC_10_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN7BL3_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN7BL3_LC_10_9_4 .LUT_INIT=16'b1111111100000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN7BL3_LC_10_9_4  (
            .in0(N__6382),
            .in1(N__5951),
            .in2(N__5870),
            .in3(N__6392),
            .lcout(\U712_CHIP_RAM.N_40 ),
            .ltout(\U712_CHIP_RAM.N_40_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUB006_0_LC_10_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUB006_0_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUB006_0_LC_10_9_5 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIUB006_0_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(N__6045),
            .in2(N__5063),
            .in3(N__6143),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_99_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3F0BF_0_LC_10_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3F0BF_0_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3F0BF_0_LC_10_9_6 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI3F0BF_0_LC_10_9_6  (
            .in0(N__6631),
            .in1(N__5060),
            .in2(N__5054),
            .in3(N__5051),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_10_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_10_0  (
            .in0(N__5756),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6039),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_1_2_LC_10_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_1_2_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_1_2_LC_10_10_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_1_2_LC_10_10_1  (
            .in0(N__6040),
            .in1(N__5958),
            .in2(_gnd_net_),
            .in3(N__6204),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_3_LC_10_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_3_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_3_LC_10_10_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_3_LC_10_10_2  (
            .in0(N__6133),
            .in1(N__5758),
            .in2(N__5045),
            .in3(N__6273),
            .lcout(\U712_CHIP_RAM.N_65 ),
            .ltout(\U712_CHIP_RAM.N_65_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_10_3 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_10_3  (
            .in0(N__5944),
            .in1(N__5042),
            .in2(N__5036),
            .in3(N__6097),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_5_LC_10_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_5_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_5_LC_10_10_4 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_5_LC_10_10_4  (
            .in0(N__5422),
            .in1(N__5399),
            .in2(N__5384),
            .in3(N__6274),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_10_5 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_10_5  (
            .in0(N__9116),
            .in1(_gnd_net_),
            .in2(N__5219),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9266),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITJ7E1_0_LC_10_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITJ7E1_0_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITJ7E1_0_LC_10_10_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITJ7E1_0_LC_10_10_6  (
            .in0(N__5755),
            .in1(N__6038),
            .in2(_gnd_net_),
            .in3(N__5943),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7Q5U5_3_LC_10_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7Q5U5_3_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7Q5U5_3_LC_10_10_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI7Q5U5_3_LC_10_10_7  (
            .in0(N__6272),
            .in1(N__5216),
            .in2(N__5210),
            .in3(N__6132),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un2_CUMBEn_LC_10_11_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un2_CUMBEn_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un2_CUMBEn_LC_10_11_0 .LUT_INIT=16'b0011011100000000;
    LogicCell40 \U712_BYTE_ENABLE.un2_CUMBEn_LC_10_11_0  (
            .in0(N__5144),
            .in1(N__5138),
            .in2(N__5117),
            .in3(N__8850),
            .lcout(\U712_BYTE_ENABLE.un2_CUMBEnZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un2_CLMBEn_LC_10_12_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un2_CLMBEn_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un2_CLMBEn_LC_10_12_1 .LUT_INIT=16'b0111010100000000;
    LogicCell40 \U712_BYTE_ENABLE.un2_CLMBEn_LC_10_12_1  (
            .in0(N__5136),
            .in1(N__5182),
            .in2(N__5113),
            .in3(N__8852),
            .lcout(\U712_BYTE_ENABLE.un2_CLMBEnZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un2_CUUBEn_LC_10_12_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un2_CUUBEn_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un2_CUUBEn_LC_10_12_2 .LUT_INIT=16'b0011000001110000;
    LogicCell40 \U712_BYTE_ENABLE.un2_CUUBEn_LC_10_12_2  (
            .in0(N__5183),
            .in1(N__5137),
            .in2(N__8863),
            .in3(N__5109),
            .lcout(\U712_BYTE_ENABLE.un2_CUUBEnZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LLBE_0_tz_LC_10_12_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LLBE_0_tz_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LLBE_0_tz_LC_10_12_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BYTE_ENABLE.LLBE_0_tz_LC_10_12_5  (
            .in0(N__5207),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5181),
            .lcout(\U712_BYTE_ENABLE.LLBE_0_0_tz ),
            .ltout(\U712_BYTE_ENABLE.LLBE_0_0_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un2_CLLBEn_LC_10_12_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un2_CLLBEn_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un2_CLLBEn_LC_10_12_6 .LUT_INIT=16'b0010101000100010;
    LogicCell40 \U712_BYTE_ENABLE.un2_CLLBEn_LC_10_12_6  (
            .in0(N__8851),
            .in1(N__5135),
            .in2(N__5120),
            .in3(N__5105),
            .lcout(\U712_BYTE_ENABLE.un2_CLLBEnZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_3_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_3_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_3_1 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_11_3_1  (
            .in0(N__8556),
            .in1(N__5258),
            .in2(_gnd_net_),
            .in3(N__8442),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9231),
            .ce(N__8645),
            .sr(N__9069));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_2 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_2  (
            .in0(N__5300),
            .in1(N__8862),
            .in2(N__5279),
            .in3(N__5246),
            .lcout(\U712_CHIP_RAM.N_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_5_3 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_5_3  (
            .in0(N__5240),
            .in1(N__8826),
            .in2(N__8118),
            .in3(N__5252),
            .lcout(\U712_CHIP_RAM.CMA_5_3_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_11_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_11_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6440),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9237),
            .ce(N__8281),
            .sr(N__9054));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_7_1 .LUT_INIT=16'b0001001000010011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_7_1  (
            .in0(N__8510),
            .in1(N__6501),
            .in2(N__8061),
            .in3(N__8389),
            .lcout(\U712_CHIP_RAM.un1_CMA31_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_7_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_7_2  (
            .in0(N__6500),
            .in1(N__8509),
            .in2(N__8417),
            .in3(N__8025),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_8_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_8_0  (
            .in0(N__6628),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5834),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_74_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_8_1 .LUT_INIT=16'b1010101100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_8_1  (
            .in0(N__5359),
            .in1(N__5342),
            .in2(N__5225),
            .in3(N__8416),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9249),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_11_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_11_8_2 .LUT_INIT=16'b1110111011101100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_11_8_2  (
            .in0(N__6629),
            .in1(N__5318),
            .in2(N__5648),
            .in3(N__6362),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_50_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_11_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_11_8_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_11_8_3  (
            .in0(N__5358),
            .in1(_gnd_net_),
            .in2(N__5222),
            .in3(N__8060),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9249),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_8_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_8_4  (
            .in0(N__6630),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6059),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_8_5 .LUT_INIT=16'b1011000111110101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_8_5  (
            .in0(N__5360),
            .in1(N__5336),
            .in2(N__8557),
            .in3(N__6627),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9249),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_11_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_11_8_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_11_8_6  (
            .in0(N__5967),
            .in1(N__6302),
            .in2(_gnd_net_),
            .in3(N__5468),
            .lcout(\U712_CHIP_RAM.N_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_11_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_11_8_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(N__6201),
            .in2(_gnd_net_),
            .in3(N__6270),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_a2_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI264TB_LC_11_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI264TB_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI264TB_LC_11_9_0 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI264TB_LC_11_9_0  (
            .in0(N__6361),
            .in1(N__5827),
            .in2(_gnd_net_),
            .in3(N__6970),
            .lcout(\U712_CHIP_RAM.N_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_9_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_9_1  (
            .in0(N__5602),
            .in1(N__5324),
            .in2(N__5972),
            .in3(N__6093),
            .lcout(\U712_CHIP_RAM.N_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIKLSF6_0_LC_11_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIKLSF6_0_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIKLSF6_0_LC_11_9_2 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIKLSF6_0_LC_11_9_2  (
            .in0(N__6051),
            .in1(N__5312),
            .in2(N__6148),
            .in3(N__9117),
            .lcout(\U712_CHIP_RAM.N_62 ),
            .ltout(\U712_CHIP_RAM.N_62_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI13TLG_0_LC_11_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI13TLG_0_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI13TLG_0_LC_11_9_3 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI13TLG_0_LC_11_9_3  (
            .in0(N__6971),
            .in1(N__5762),
            .in2(N__5306),
            .in3(N__7015),
            .lcout(\U712_CHIP_RAM.N_13 ),
            .ltout(\U712_CHIP_RAM.N_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_9_4 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_9_4  (
            .in0(N__5423),
            .in1(_gnd_net_),
            .in2(N__5303),
            .in3(N__6282),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9254),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_9_5 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_9_5  (
            .in0(N__5962),
            .in1(N__5449),
            .in2(N__6220),
            .in3(N__6052),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9254),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_11_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_11_9_6 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_11_9_6  (
            .in0(N__5862),
            .in1(N__5630),
            .in2(_gnd_net_),
            .in3(N__5618),
            .lcout(\U712_CHIP_RAM.N_44 ),
            .ltout(\U712_CHIP_RAM.N_44_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNIOG801_LC_11_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNIOG801_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNIOG801_LC_11_9_7 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_RNIOG801_LC_11_9_7  (
            .in0(N__6626),
            .in1(_gnd_net_),
            .in2(N__5471),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_10_0 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_10_0  (
            .in0(N__6056),
            .in1(N__5963),
            .in2(_gnd_net_),
            .in3(N__5450),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9261),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_10_1 .LUT_INIT=16'b1111000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_10_1  (
            .in0(N__5764),
            .in1(N__5551),
            .in2(N__6062),
            .in3(N__6976),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_0_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_11_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_11_10_2 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_11_10_2  (
            .in0(N__5438),
            .in1(_gnd_net_),
            .in2(N__5432),
            .in3(N__5429),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9261),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_10_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_10_3  (
            .in0(N__5583),
            .in1(N__5397),
            .in2(N__5570),
            .in3(N__5378),
            .lcout(\U712_CHIP_RAM.N_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_10_4 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_10_4  (
            .in0(N__5380),
            .in1(N__5421),
            .in2(N__6287),
            .in3(N__9111),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9261),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_11_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_11_10_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_11_10_5  (
            .in0(N__5420),
            .in1(N__5398),
            .in2(N__6283),
            .in3(N__5379),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_10_6 .LUT_INIT=16'b0000001100110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__9112),
            .in2(N__5363),
            .in3(N__5584),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9261),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_10_7 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_10_7  (
            .in0(N__5591),
            .in1(N__5585),
            .in2(N__9122),
            .in3(N__5569),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9261),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_11_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_11_11_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__9110),
            .in2(_gnd_net_),
            .in3(N__6999),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBDIR_RNO_0_LC_11_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_RNO_0_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBDIR_RNO_0_LC_11_11_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_RNO_0_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__5555),
            .in2(_gnd_net_),
            .in3(N__5765),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_LC_11_11_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_LC_11_11_4 .LUT_INIT=16'b0100010101010101;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_LC_11_11_4  (
            .in0(N__5540),
            .in1(N__7079),
            .in2(N__7460),
            .in3(N__7566),
            .lcout(CLLBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIH4474_LC_11_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIH4474_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIH4474_LC_11_11_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIH4474_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(N__7135),
            .in2(_gnd_net_),
            .in3(N__6972),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_LC_11_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_11_12_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_11_12_3 .LUT_INIT=16'b0100111011101110;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_11_12_3  (
            .in0(N__7014),
            .in1(N__7565),
            .in2(N__7694),
            .in3(N__5513),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9273),
            .ce(),
            .sr(N__9013));
    defparam \U712_CHIP_RAM.DBDIR_LC_11_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_11_12_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_11_12_5 .LUT_INIT=16'b1011000111110000;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_11_12_5  (
            .in0(N__6982),
            .in1(N__6343),
            .in2(N__6682),
            .in3(N__5507),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9273),
            .ce(),
            .sr(N__9013));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_12_4_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_12_4_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_12_4_1 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_12_4_1  (
            .in0(N__5777),
            .in1(N__8575),
            .in2(_gnd_net_),
            .in3(N__8454),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9230),
            .ce(N__8616),
            .sr(N__9057));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_5_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_5_2  (
            .in0(N__9120),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5480),
            .lcout(\U712_CHIP_RAM.un1_CMA31_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_5_5 .LUT_INIT=16'b1110001000110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_5_5  (
            .in0(N__5816),
            .in1(N__5771),
            .in2(N__5801),
            .in3(N__8838),
            .lcout(\U712_CHIP_RAM.N_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_6_5 .LUT_INIT=16'b0000101101011011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_6_5  (
            .in0(N__8787),
            .in1(N__6446),
            .in2(N__8114),
            .in3(N__6401),
            .lcout(\U712_CHIP_RAM.CMA_5_3_ns_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_12_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_12_8_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_12_8_0  (
            .in0(N__6060),
            .in1(N__5757),
            .in2(_gnd_net_),
            .in3(N__5970),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_0_LC_12_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_0_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_0_LC_12_8_6 .LUT_INIT=16'b0000001000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_0_LC_12_8_6  (
            .in0(N__6061),
            .in1(N__5603),
            .in2(N__6098),
            .in3(N__5971),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_12_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_12_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_12_9_0 .LUT_INIT=16'b1111001111111011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_12_9_0  (
            .in0(N__5717),
            .in1(N__5699),
            .in2(N__5687),
            .in3(N__5666),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9248),
            .ce(),
            .sr(N__9018));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_12_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_12_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_12_9_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_12_9_1  (
            .in0(N__8794),
            .in1(N__5654),
            .in2(_gnd_net_),
            .in3(N__7470),
            .lcout(\U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9248),
            .ce(),
            .sr(N__9018));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_LC_12_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_LC_12_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_LC_12_9_2 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_LC_12_9_2  (
            .in0(N__5617),
            .in1(N__5644),
            .in2(_gnd_net_),
            .in3(N__6983),
            .lcout(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9248),
            .ce(),
            .sr(N__9018));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_0_LC_12_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_0_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_0_LC_12_9_3 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_0_LC_12_9_3  (
            .in0(N__5859),
            .in1(N__5629),
            .in2(_gnd_net_),
            .in3(N__5616),
            .lcout(\U712_CHIP_RAM.N_47 ),
            .ltout(\U712_CHIP_RAM.N_47_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_2_LC_12_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_2_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_2_LC_12_9_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_2_LC_12_9_4  (
            .in0(N__6197),
            .in1(N__5932),
            .in2(N__6395),
            .in3(N__6268),
            .lcout(\U712_CHIP_RAM.N_89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_12_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_12_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_12_9_5 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_12_9_5  (
            .in0(N__5861),
            .in1(N__6371),
            .in2(_gnd_net_),
            .in3(N__6383),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9248),
            .ce(),
            .sr(N__9018));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI0CV43_LC_12_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI0CV43_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI0CV43_LC_12_9_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI0CV43_LC_12_9_6  (
            .in0(N__5945),
            .in1(N__6041),
            .in2(N__6147),
            .in3(N__5860),
            .lcout(\U712_CHIP_RAM.N_100 ),
            .ltout(\U712_CHIP_RAM.N_100_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_2_LC_12_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_2_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_2_LC_12_9_7 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_2_LC_12_9_7  (
            .in0(N__6269),
            .in1(_gnd_net_),
            .in2(N__6365),
            .in3(N__6198),
            .lcout(\U712_CHIP_RAM.N_101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_12_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_12_10_2 .LUT_INIT=16'b1100010011110101;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_12_10_2  (
            .in0(N__7439),
            .in1(N__6758),
            .in2(N__6350),
            .in3(N__8849),
            .lcout(),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_12_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_12_10_3 .LUT_INIT=16'b1100110001001110;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_12_10_3  (
            .in0(N__6314),
            .in1(N__6301),
            .in2(N__6305),
            .in3(N__6086),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9251),
            .ce(),
            .sr(N__9014));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_12_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_12_10_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_12_10_5  (
            .in0(N__6042),
            .in1(N__5968),
            .in2(_gnd_net_),
            .in3(N__6085),
            .lcout(\U712_CHIP_RAM.N_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_12_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_12_10_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_12_10_6  (
            .in0(N__6271),
            .in1(N__6200),
            .in2(_gnd_net_),
            .in3(N__6131),
            .lcout(\U712_CHIP_RAM.N_42 ),
            .ltout(\U712_CHIP_RAM.N_42_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_12_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_12_10_7 .LUT_INIT=16'b0000100000000101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_12_10_7  (
            .in0(N__6043),
            .in1(N__5969),
            .in2(N__5873),
            .in3(N__5866),
            .lcout(\U712_CHIP_RAM.N_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_12_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_12_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_12_11_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__7136),
            .in2(_gnd_net_),
            .in3(N__6977),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9258),
            .ce(N__6767),
            .sr(N__9012));
    defparam \U712_BUFFERS.DRDDIR_0_i_LC_12_12_4 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_0_i_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_0_i_LC_12_12_4 .LUT_INIT=16'b0111001101010000;
    LogicCell40 \U712_BUFFERS.DRDDIR_0_i_LC_12_12_4  (
            .in0(N__6757),
            .in1(N__6678),
            .in2(N__7511),
            .in3(N__7440),
            .lcout(DRDDIR_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_5.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_5.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_19_5 (
            .in0(N__6624),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CRCSn_LC_13_3_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_13_3_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_13_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_13_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6520),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9232),
            .ce(),
            .sr(N__9070));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_13_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_13_4_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_13_4_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_13_4_4  (
            .in0(N__8574),
            .in1(N__8119),
            .in2(N__8471),
            .in3(N__6521),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9233),
            .ce(N__8621),
            .sr(N__9066));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_13_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_13_5_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_13_5_1 .LUT_INIT=16'b1111110100000001;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_13_5_1  (
            .in0(N__8123),
            .in1(N__8576),
            .in2(N__8472),
            .in3(N__7196),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9234),
            .ce(N__8617),
            .sr(N__9062));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_13_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_13_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_13_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7385),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9238),
            .ce(N__8280),
            .sr(N__9055));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_7_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_7_0  (
            .in0(N__6436),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9246),
            .ce(N__7957),
            .sr(N__9043));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7904),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9246),
            .ce(N__7957),
            .sr(N__9043));
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_13_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_13_9_0 .LUT_INIT=16'b0100010001001110;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_LC_13_9_0  (
            .in0(N__7016),
            .in1(N__8768),
            .in2(N__7132),
            .in3(N__6981),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9255),
            .ce(),
            .sr(N__9024));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_14_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_14_4_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_14_4_0 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_14_4_0  (
            .in0(N__7250),
            .in1(N__8841),
            .in2(N__8134),
            .in3(N__7352),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_14_4_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_14_4_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_14_4_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_14_4_1  (
            .in0(N__8842),
            .in1(N__6932),
            .in2(N__6917),
            .in3(N__6914),
            .lcout(\U712_CHIP_RAM.N_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_14_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_14_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_14_5_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_14_5_2  (
            .in0(N__8583),
            .in1(N__7145),
            .in2(_gnd_net_),
            .in3(N__8461),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9239),
            .ce(N__8653),
            .sr(N__9067));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_14_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_14_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_14_5_6 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_14_5_6  (
            .in0(N__8584),
            .in1(N__6818),
            .in2(_gnd_net_),
            .in3(N__8462),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9239),
            .ce(N__8653),
            .sr(N__9067));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_14_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_14_6_3 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_14_6_3  (
            .in0(N__6857),
            .in1(N__8844),
            .in2(N__6836),
            .in3(N__7235),
            .lcout(\U712_CHIP_RAM.N_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_14_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_14_6_5 .LUT_INIT=16'b1101010110010001;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_14_6_5  (
            .in0(N__6773),
            .in1(N__8843),
            .in2(N__6812),
            .in3(N__6788),
            .lcout(\U712_CHIP_RAM.N_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_7_0 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_7_0  (
            .in0(N__7877),
            .in1(N__8795),
            .in2(N__8124),
            .in3(N__7841),
            .lcout(\U712_CHIP_RAM.CMA_5_3_ns_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_14_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_14_7_4 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_14_7_4  (
            .in0(N__8294),
            .in1(N__8796),
            .in2(N__8125),
            .in3(N__7241),
            .lcout(\U712_CHIP_RAM.CMA_5_3_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_14_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_14_8_3 .LUT_INIT=16'b0000101101011011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_14_8_3  (
            .in0(N__8765),
            .in1(N__7757),
            .in2(N__8116),
            .in3(N__7829),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_14_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_14_8_4 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_14_8_4  (
            .in0(N__7229),
            .in1(N__7214),
            .in2(N__7199),
            .in3(N__8766),
            .lcout(\U712_CHIP_RAM.N_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_14_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_14_8_6 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_14_8_6  (
            .in0(N__7796),
            .in1(N__8764),
            .in2(N__8115),
            .in3(N__7835),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_14_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_14_8_7 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_14_8_7  (
            .in0(N__7187),
            .in1(N__7169),
            .in2(N__7148),
            .in3(N__8767),
            .lcout(\U712_CHIP_RAM.N_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_14_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_14_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_14_9_6 .LUT_INIT=16'b0111010100110000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_14_9_6  (
            .in0(N__7751),
            .in1(N__7469),
            .in2(N__7134),
            .in3(N__7733),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9262),
            .ce(),
            .sr(N__9037));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_14_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_14_10_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_14_10_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_14_10_1  (
            .in0(N__7078),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7628),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9267),
            .ce(),
            .sr(N__9025));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_14_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_14_10_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_14_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_14_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7750),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9267),
            .ce(),
            .sr(N__9025));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_LC_14_11_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_LC_14_11_1 .LUT_INIT=16'b0101010101000101;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_LC_14_11_1  (
            .in0(N__7088),
            .in1(N__7592),
            .in2(N__7471),
            .in3(N__7074),
            .lcout(CUMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_LC_14_11_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_LC_14_11_5 .LUT_INIT=16'b0000000011011111;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_LC_14_11_5  (
            .in0(N__7461),
            .in1(N__7626),
            .in2(N__7596),
            .in3(N__7661),
            .lcout(CLMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_LC_14_11_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_LC_14_11_7 .LUT_INIT=16'b0000000011111101;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_LC_14_11_7  (
            .in0(N__7465),
            .in1(N__7627),
            .in2(N__7597),
            .in3(N__7544),
            .lcout(CUUBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.N_52_i_LC_14_12_1 .C_ON=1'b0;
    defparam \U712_BUFFERS.N_52_i_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.N_52_i_LC_14_12_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_BUFFERS.N_52_i_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(N__7507),
            .in2(_gnd_net_),
            .in3(N__7472),
            .lcout(N_52_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_4_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_4_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7384),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9240),
            .ce(N__7956),
            .sr(N__9076));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_15_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_15_5_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_15_5_1 .LUT_INIT=16'b1010101010100011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_15_5_1  (
            .in0(N__7346),
            .in1(N__8129),
            .in2(N__8473),
            .in3(N__8582),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9247),
            .ce(N__8633),
            .sr(N__9071));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_15_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_15_5_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_15_5_5 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_15_5_5  (
            .in0(N__7319),
            .in1(_gnd_net_),
            .in2(N__8474),
            .in3(N__8581),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9247),
            .ce(N__8633),
            .sr(N__9071));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_15_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_15_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_15_5_6 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_15_5_6  (
            .in0(N__7292),
            .in1(N__8342),
            .in2(N__9335),
            .in3(N__8839),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9247),
            .ce(N__8633),
            .sr(N__9071));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_15_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_15_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_15_7_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_15_7_3  (
            .in0(N__8180),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9256),
            .ce(N__8266),
            .sr(N__9063));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_15_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_15_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_15_7_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_15_7_6  (
            .in0(N__7900),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9256),
            .ce(N__8266),
            .sr(N__9063));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_8_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_8_2  (
            .in0(N__7864),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9263),
            .ce(N__7941),
            .sr(N__9056));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_8_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_8_3  (
            .in0(N__7721),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9263),
            .ce(N__7941),
            .sr(N__9056));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7823),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9263),
            .ce(N__7941),
            .sr(N__9056));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_15_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_15_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_15_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_15_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7816),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9268),
            .ce(N__8250),
            .sr(N__9044));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_15_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_15_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_15_9_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_15_9_4  (
            .in0(N__7790),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9268),
            .ce(N__8250),
            .sr(N__9044));
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_15_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_15_10_2 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_15_10_2  (
            .in0(N__9118),
            .in1(N__7749),
            .in2(_gnd_net_),
            .in3(N__7732),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_15_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_15_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_15_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_15_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7717),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9277),
            .ce(N__8251),
            .sr(N__9026));
    defparam \U712_CHIP_RAM.RASn_LC_16_2_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_16_2_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_16_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_16_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8585),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9235),
            .ce(),
            .sr(N__9080));
    defparam \U712_CHIP_RAM.WEn_LC_16_3_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_16_3_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_16_3_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_16_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8470),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9241),
            .ce(),
            .sr(N__9079));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_16_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_16_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_16_5_2 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_16_5_2  (
            .in0(N__8879),
            .in1(N__8341),
            .in2(N__8147),
            .in3(N__8840),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9250),
            .ce(N__8654),
            .sr(N__9077));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_16_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_16_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_16_6_7 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_16_6_7  (
            .in0(N__8577),
            .in1(N__8117),
            .in2(_gnd_net_),
            .in3(N__8463),
            .lcout(\U712_CHIP_RAM.CMA_5_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_16_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_16_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_16_7_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_16_7_7  (
            .in0(N__8323),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9264),
            .ce(N__8279),
            .sr(N__9068));
    defparam CONSTANT_ONE_LUT4_LC_17_5_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_17_5_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_17_5_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_17_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_17_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_17_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_17_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_17_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8176),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9269),
            .ce(N__7931),
            .sr(N__9072));
    defparam \U712_CHIP_RAM.CASn_LC_18_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_18_4_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_18_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_18_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8135),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9257),
            .ce(),
            .sr(N__9081));
    defparam \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_18_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_18_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_18_8_3 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_18_8_3  (
            .in0(N__9121),
            .in1(N__7910),
            .in2(_gnd_net_),
            .in3(N__9298),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_19_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_19_8_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_19_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_1_LC_19_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9299),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9280),
            .ce(),
            .sr(N__9078));
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_19_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_19_8_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_19_8_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_0_LC_19_8_7  (
            .in0(N__9328),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9308),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9280),
            .ce(),
            .sr(N__9078));
endmodule // U712_TOP

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Apr 28 2025 13:13:51

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DA : out std_logic_vector(2 downto 0);
    A : in std_logic_vector(20 downto 0);
    DBRn : in std_logic;
    RAMENn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    TCIn : out std_logic;
    TBIn : out std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__12519\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12382\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12211\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \REGENn_c\ : std_logic;
signal \U712_REG_SM.START_RSTZ0\ : std_logic;
signal \U712_REG_SM.un6_REG_CYCLE_START_cascade_\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_1_sqmuxa_1\ : std_logic;
signal \U712_REG_SM.N_188\ : std_logic;
signal \U712_REG_SM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\ : std_logic;
signal \U712_REG_SM.N_157_cascade_\ : std_logic;
signal \U712_REG_SM.N_109_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTc_0_0_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_0_sqmuxa_cascade_\ : std_logic;
signal \U712_REG_SM.N_185\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.N_109_0\ : std_logic;
signal \U712_REG_SM.N_105_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_1\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_166\ : std_logic;
signal \LDSn_c\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.un2_DBR_COUNT_cry_1\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.un2_DBR_COUNT_cry_2\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.un2_DBR_COUNT_cry_3\ : std_logic;
signal \U712_CHIP_RAM.un2_DBR_COUNT_cry_4\ : std_logic;
signal \U712_CHIP_RAM.un2_DBR_COUNT_cry_5\ : std_logic;
signal \U712_CHIP_RAM.un2_DBR_COUNT_cry_6\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_159\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_0\ : std_logic;
signal \U712_REG_SM.N_109\ : std_logic;
signal \U712_REG_SM.N_164\ : std_logic;
signal \U712_REG_SM.N_80\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_96\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.N_96_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \UDSn_c\ : std_logic;
signal \U712_BYTE_ENABLE_UDS_0\ : std_logic;
signal \U712_REG_SM.N_163\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \U712_CYCLE_TERM.N_51_cascade_\ : std_logic;
signal \U712_CHIP_RAM.BANK0_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_0_cascade_\ : std_logic;
signal \LATCH_CLK_c\ : std_logic;
signal \U712_CHIP_RAM.N_144_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_4\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_3\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.N_163_0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_CYCLE_TERM.N_47_0\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \bfn_10_9_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_START_2_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.N_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER18_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER33_1_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_i_0_68_i_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_64_cascade_\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER18\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_1\ : std_logic;
signal \U712_CHIP_RAM.LATCH_CLK_6\ : std_logic;
signal \bfn_10_13_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.N_64\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ1Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \CLMBEn_c\ : std_logic;
signal \U712_CHIP_RAM.LATCH_CLK_0_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.LATCH_CLK_0_sqmuxa_cascade_\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER42_7_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER42_7_0_cascade_\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_152\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_108_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_i_0_68_i_a3_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_i_0_68_i_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER42_0_cascade_\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER42_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.N_331_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER37_0_a3_1_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_7_2\ : std_logic;
signal \U712_CHIP_RAM.BANK0_7_0_cascade_\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.A_m_20\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_\ : std_logic;
signal \U712_CHIP_RAM.A_m_2_20\ : std_logic;
signal \U712_CHIP_RAM.N_94_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_187\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERlde_0_a3_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a3_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_155\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a3_1\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_cascade_\ : std_logic;
signal \U712_BYTE_ENABLE.N_58\ : std_logic;
signal \N_56_i\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \A_c_1\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \N_58_i\ : std_logic;
signal \DMA_LATCH_EN_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER42_7_0_0\ : std_logic;
signal \A_c_8\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_13\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_5_0\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_DISABLEZ0\ : std_logic;
signal \U712_CHIP_RAM.N_95\ : std_logic;
signal \U712_CHIP_RAM.N_119\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.N_95_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_3_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_3_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_cascade_\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_7\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER38_1_0\ : std_logic;
signal \U712_CHIP_RAM.N_94\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER42_4_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_7_0\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \A_c_7\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.N_173\ : std_logic;
signal \U712_CHIP_RAM.un3_CPU_CYCLE_START\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_177\ : std_logic;
signal \U712_CHIP_RAM.N_172\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_1_sqmuxa_1_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_186\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER34\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER34_cascade_\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER16_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER17_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER15\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER17_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_33\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER19_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER17_1_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.N_38_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_i_1_1\ : std_logic;
signal \U712_CHIP_RAM.N_151\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER19_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_i\ : std_logic;
signal \U712_CHIP_RAM.N_331_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_29_i_a2_i_1\ : std_logic;
signal \U712_CHIP_RAM.N_61_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_218\ : std_logic;
signal \U712_CHIP_RAM.N_154\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_29_i_a2_i_1_0\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \UMBEn_c\ : std_logic;
signal \U712_BYTE_ENABLE.un3_CUMBEnZ0Z_1_cascade_\ : std_logic;
signal \CUMBEn_c\ : std_logic;
signal \UUBEn_c\ : std_logic;
signal \U712_BYTE_ENABLE.un3_CUMBEnZ0Z_1\ : std_logic;
signal \CUUBEn_c\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_56\ : std_logic;
signal \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_0_cascade_\ : std_logic;
signal \CLLBEn_c\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.N_11_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_12\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_11\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z20\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A20C_net\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_0\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \RnW_c\ : std_logic;
signal \WRITE_CYCLEm\ : std_logic;
signal \DRDDIR_c\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \DA_wire\ : std_logic_vector(2 downto 0);
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    TBIn <= \TBIn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    ASn <= \ASn_wire\;
    DA <= \DA_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    TCIn <= \TCIn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__4259\,
            RESETB => \N__5831\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12519\,
            DIN => \N__12518\,
            DOUT => \N__12517\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12519\,
            PADOUT => \N__12518\,
            PADIN => \N__12517\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8723\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12510\,
            DIN => \N__12509\,
            DOUT => \N__12508\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12510\,
            PADOUT => \N__12509\,
            PADIN => \N__12508\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12501\,
            DIN => \N__12500\,
            DOUT => \N__12499\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12501\,
            PADOUT => \N__12500\,
            PADIN => \N__12499\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9554\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12492\,
            DIN => \N__12491\,
            DOUT => \N__12490\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12492\,
            PADOUT => \N__12491\,
            PADIN => \N__12490\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10682\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12483\,
            DIN => \N__12482\,
            DOUT => \N__12481\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12483\,
            PADOUT => \N__12482\,
            PADIN => \N__12481\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12474\,
            DIN => \N__12473\,
            DOUT => \N__12472\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12474\,
            PADOUT => \N__12473\,
            PADIN => \N__12472\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12465\,
            DIN => \N__12464\,
            DOUT => \N__12463\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12465\,
            PADOUT => \N__12464\,
            PADIN => \N__12463\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12456\,
            DIN => \N__12455\,
            DOUT => \N__12454\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12456\,
            PADOUT => \N__12455\,
            PADIN => \N__12454\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12447\,
            DIN => \N__12446\,
            DOUT => \N__12445\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12447\,
            PADOUT => \N__12446\,
            PADIN => \N__12445\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12438\,
            DIN => \N__12437\,
            DOUT => \N__12436\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12438\,
            PADOUT => \N__12437\,
            PADIN => \N__12436\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12429\,
            DIN => \N__12428\,
            DOUT => \N__12427\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12429\,
            PADOUT => \N__12428\,
            PADIN => \N__12427\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10364\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12420\,
            DIN => \N__12419\,
            DOUT => \N__12418\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12420\,
            PADOUT => \N__12419\,
            PADIN => \N__12418\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8779\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12411\,
            DIN => \N__12410\,
            DOUT => \N__12409\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12411\,
            PADOUT => \N__12410\,
            PADIN => \N__12409\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12402\,
            DIN => \N__12401\,
            DOUT => \N__12400\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12402\,
            PADOUT => \N__12401\,
            PADIN => \N__12400\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5371\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12393\,
            DIN => \N__12392\,
            DOUT => \N__12391\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12393\,
            PADOUT => \N__12392\,
            PADIN => \N__12391\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12384\,
            DIN => \N__12383\,
            DOUT => \N__12382\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12384\,
            PADOUT => \N__12383\,
            PADIN => \N__12382\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12375\,
            DIN => \N__12374\,
            DOUT => \N__12373\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12375\,
            PADOUT => \N__12374\,
            PADIN => \N__12373\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5348\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12366\,
            DIN => \N__12365\,
            DOUT => \N__12364\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12366\,
            PADOUT => \N__12365\,
            PADIN => \N__12364\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12357\,
            DIN => \N__12356\,
            DOUT => \N__12355\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12357\,
            PADOUT => \N__12356\,
            PADIN => \N__12355\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12348\,
            DIN => \N__12347\,
            DOUT => \N__12346\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12348\,
            PADOUT => \N__12347\,
            PADIN => \N__12346\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9143\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12339\,
            DIN => \N__12338\,
            DOUT => \N__12337\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12339\,
            PADOUT => \N__12338\,
            PADIN => \N__12337\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12330\,
            DIN => \N__12329\,
            DOUT => \N__12328\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12330\,
            PADOUT => \N__12329\,
            PADIN => \N__12328\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9455\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12321\,
            DIN => \N__12320\,
            DOUT => \N__12319\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12321\,
            PADOUT => \N__12320\,
            PADIN => \N__12319\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12312\,
            DIN => \N__12311\,
            DOUT => \N__12310\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12312\,
            PADOUT => \N__12311\,
            PADIN => \N__12310\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7031\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12303\,
            DIN => \N__12302\,
            DOUT => \N__12301\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12303\,
            PADOUT => \N__12302\,
            PADIN => \N__12301\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5319\,
            DIN0 => OPEN,
            DOUT0 => \N__5257\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12294\,
            DIN => \N__12293\,
            DOUT => \N__12292\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12294\,
            PADOUT => \N__12293\,
            PADIN => \N__12292\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12285\,
            DIN => \N__12284\,
            DOUT => \N__12283\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12285\,
            PADOUT => \N__12284\,
            PADIN => \N__12283\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12276\,
            DIN => \N__12275\,
            DOUT => \N__12274\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12276\,
            PADOUT => \N__12275\,
            PADIN => \N__12274\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12267\,
            DIN => \N__12266\,
            DOUT => \N__12265\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12267\,
            PADOUT => \N__12266\,
            PADIN => \N__12265\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12258\,
            DIN => \N__12257\,
            DOUT => \N__12256\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12258\,
            PADOUT => \N__12257\,
            PADIN => \N__12256\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12249\,
            DIN => \N__12248\,
            DOUT => \N__12247\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12249\,
            PADOUT => \N__12248\,
            PADIN => \N__12247\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6728\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12240\,
            DIN => \N__12239\,
            DOUT => \N__12238\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12240\,
            PADOUT => \N__12239\,
            PADIN => \N__12238\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12231\,
            DIN => \N__12230\,
            DOUT => \N__12229\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12231\,
            PADOUT => \N__12230\,
            PADIN => \N__12229\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12222\,
            DIN => \N__12221\,
            DOUT => \N__12220\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12222\,
            PADOUT => \N__12221\,
            PADIN => \N__12220\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12213\,
            DIN => \N__12212\,
            DOUT => \N__12211\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12213\,
            PADOUT => \N__12212\,
            PADIN => \N__12211\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12204\,
            DIN => \N__12203\,
            DOUT => \N__12202\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12204\,
            PADOUT => \N__12203\,
            PADIN => \N__12202\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12195\,
            DIN => \N__12194\,
            DOUT => \N__12193\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12195\,
            PADOUT => \N__12194\,
            PADIN => \N__12193\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9719\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12186\,
            DIN => \N__12185\,
            DOUT => \N__12184\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12186\,
            PADOUT => \N__12185\,
            PADIN => \N__12184\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6503\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12177\,
            DIN => \N__12176\,
            DOUT => \N__12175\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12177\,
            PADOUT => \N__12176\,
            PADIN => \N__12175\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12168\,
            DIN => \N__12167\,
            DOUT => \N__12166\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12168\,
            PADOUT => \N__12167\,
            PADIN => \N__12166\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5441\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12159\,
            DIN => \N__12158\,
            DOUT => \N__12157\,
            PACKAGEPIN => \DA_wire\(0)
        );

    \DA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12159\,
            PADOUT => \N__12158\,
            PADIN => \N__12157\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7442\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12150\,
            DIN => \N__12149\,
            DOUT => \N__12148\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12150\,
            PADOUT => \N__12149\,
            PADIN => \N__12148\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12141\,
            DIN => \N__12140\,
            DOUT => \N__12139\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12141\,
            PADOUT => \N__12140\,
            PADIN => \N__12139\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8849\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12132\,
            DIN => \N__12131\,
            DOUT => \N__12130\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12132\,
            PADOUT => \N__12131\,
            PADIN => \N__12130\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10487\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12123\,
            DIN => \N__12122\,
            DOUT => \N__12121\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12123\,
            PADOUT => \N__12122\,
            PADIN => \N__12121\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11618\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12114\,
            DIN => \N__12113\,
            DOUT => \N__12112\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12114\,
            PADOUT => \N__12113\,
            PADIN => \N__12112\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8627\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12105\,
            DIN => \N__12104\,
            DOUT => \N__12103\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12105\,
            PADOUT => \N__12104\,
            PADIN => \N__12103\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9383\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12096\,
            DIN => \N__12095\,
            DOUT => \N__12094\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12096\,
            PADOUT => \N__12095\,
            PADIN => \N__12094\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4412\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12087\,
            DIN => \N__12086\,
            DOUT => \N__12085\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12087\,
            PADOUT => \N__12086\,
            PADIN => \N__12085\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12078\,
            DIN => \N__12077\,
            DOUT => \N__12076\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12078\,
            PADOUT => \N__12077\,
            PADIN => \N__12076\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12069\,
            DIN => \N__12068\,
            DOUT => \N__12067\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12069\,
            PADOUT => \N__12068\,
            PADIN => \N__12067\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6014\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12060\,
            DIN => \N__12059\,
            DOUT => \N__12058\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12060\,
            PADOUT => \N__12059\,
            PADIN => \N__12058\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5323\,
            DIN0 => OPEN,
            DOUT0 => \N__5258\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12051\,
            DIN => \N__12050\,
            DOUT => \N__12049\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12051\,
            PADOUT => \N__12050\,
            PADIN => \N__12049\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9800\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12042\,
            DIN => \N__12041\,
            DOUT => \N__12040\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12042\,
            PADOUT => \N__12041\,
            PADIN => \N__12040\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4679\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12033\,
            DIN => \N__12032\,
            DOUT => \N__12031\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12033\,
            PADOUT => \N__12032\,
            PADIN => \N__12031\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8798\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12024\,
            DIN => \N__12023\,
            DOUT => \N__12022\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12024\,
            PADOUT => \N__12023\,
            PADIN => \N__12022\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12015\,
            DIN => \N__12014\,
            DOUT => \N__12013\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12015\,
            PADOUT => \N__12014\,
            PADIN => \N__12013\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12006\,
            DIN => \N__12005\,
            DOUT => \N__12004\,
            PACKAGEPIN => \DA_wire\(2)
        );

    \DA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12006\,
            PADOUT => \N__12005\,
            PADIN => \N__12004\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8897\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11997\,
            DIN => \N__11996\,
            DOUT => \N__11995\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11997\,
            PADOUT => \N__11996\,
            PADIN => \N__11995\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11988\,
            DIN => \N__11987\,
            DOUT => \N__11986\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11988\,
            PADOUT => \N__11987\,
            PADIN => \N__11986\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11979\,
            DIN => \N__11978\,
            DOUT => \N__11977\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11979\,
            PADOUT => \N__11978\,
            PADIN => \N__11977\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8606\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11970\,
            DIN => \N__11969\,
            DOUT => \N__11968\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11970\,
            PADOUT => \N__11969\,
            PADIN => \N__11968\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6746\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11961\,
            DIN => \N__11960\,
            DOUT => \N__11959\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11961\,
            PADOUT => \N__11960\,
            PADIN => \N__11959\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11952\,
            DIN => \N__11951\,
            DOUT => \N__11950\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11952\,
            PADOUT => \N__11951\,
            PADIN => \N__11950\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8744\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11943\,
            DIN => \N__11942\,
            DOUT => \N__11941\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11943\,
            PADOUT => \N__11942\,
            PADIN => \N__11941\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5324\,
            DIN0 => OPEN,
            DOUT0 => \N__5253\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11934\,
            DIN => \N__11933\,
            DOUT => \N__11932\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11934\,
            PADOUT => \N__11933\,
            PADIN => \N__11932\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9950\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11925\,
            DIN => \N__11924\,
            DOUT => \N__11923\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11925\,
            PADOUT => \N__11924\,
            PADIN => \N__11923\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11916\,
            DIN => \N__11915\,
            DOUT => \N__11914\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11916\,
            PADOUT => \N__11915\,
            PADIN => \N__11914\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11907\,
            DIN => \N__11906\,
            DOUT => \N__11905\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11907\,
            PADOUT => \N__11906\,
            PADIN => \N__11905\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9101\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11898\,
            DIN => \N__11897\,
            DOUT => \N__11896\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11898\,
            PADOUT => \N__11897\,
            PADIN => \N__11896\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11889\,
            DIN => \N__11888\,
            DOUT => \N__11887\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11889\,
            PADOUT => \N__11888\,
            PADIN => \N__11887\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11880\,
            DIN => \N__11879\,
            DOUT => \N__11878\,
            PACKAGEPIN => \DA_wire\(1)
        );

    \DA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11880\,
            PADOUT => \N__11879\,
            PADIN => \N__11878\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9002\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11871\,
            DIN => \N__11870\,
            DOUT => \N__11869\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11871\,
            PADOUT => \N__11870\,
            PADIN => \N__11869\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11862\,
            DIN => \N__11861\,
            DOUT => \N__11860\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11862\,
            PADOUT => \N__11861\,
            PADIN => \N__11860\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11853\,
            DIN => \N__11852\,
            DOUT => \N__11851\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11853\,
            PADOUT => \N__11852\,
            PADIN => \N__11851\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9062\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11844\,
            DIN => \N__11843\,
            DOUT => \N__11842\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11844\,
            PADOUT => \N__11843\,
            PADIN => \N__11842\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4757\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11835\,
            DIN => \N__11834\,
            DOUT => \N__11833\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11835\,
            PADOUT => \N__11834\,
            PADIN => \N__11833\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8837\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11826\,
            DIN => \N__11825\,
            DOUT => \N__11824\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11826\,
            PADOUT => \N__11825\,
            PADIN => \N__11824\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6419\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11817\,
            DIN => \N__11816\,
            DOUT => \N__11815\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11817\,
            PADOUT => \N__11816\,
            PADIN => \N__11815\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11808\,
            DIN => \N__11807\,
            DOUT => \N__11806\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11808\,
            PADOUT => \N__11807\,
            PADIN => \N__11806\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11799\,
            DIN => \N__11798\,
            DOUT => \N__11797\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11799\,
            PADOUT => \N__11798\,
            PADIN => \N__11797\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10508\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11790\,
            DIN => \N__11789\,
            DOUT => \N__11788\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11790\,
            PADOUT => \N__11789\,
            PADIN => \N__11788\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11781\,
            DIN => \N__11780\,
            DOUT => \N__11779\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11781\,
            PADOUT => \N__11780\,
            PADIN => \N__11779\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11772\,
            DIN => \N__11771\,
            DOUT => \N__11770\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11772\,
            PADOUT => \N__11771\,
            PADIN => \N__11770\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5156\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11763\,
            DIN => \N__11762\,
            DOUT => \N__11761\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11763\,
            PADOUT => \N__11762\,
            PADIN => \N__11761\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4709\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11754\,
            DIN => \N__11753\,
            DOUT => \N__11752\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11754\,
            PADOUT => \N__11753\,
            PADIN => \N__11752\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5102\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11745\,
            DIN => \N__11744\,
            DOUT => \N__11743\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11745\,
            PADOUT => \N__11744\,
            PADIN => \N__11743\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11736\,
            DIN => \N__11735\,
            DOUT => \N__11734\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11736\,
            PADOUT => \N__11735\,
            PADIN => \N__11734\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5101\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11727\,
            DIN => \N__11726\,
            DOUT => \N__11725\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11727\,
            PADOUT => \N__11726\,
            PADIN => \N__11725\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4280\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11718\,
            DIN => \N__11717\,
            DOUT => \N__11716\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11718\,
            PADOUT => \N__11717\,
            PADIN => \N__11716\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9926\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11709\,
            DIN => \N__11708\,
            DOUT => \N__11707\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11709\,
            PADOUT => \N__11708\,
            PADIN => \N__11707\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11700\,
            DIN => \N__11699\,
            DOUT => \N__11698\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11700\,
            PADOUT => \N__11699\,
            PADIN => \N__11698\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11691\,
            DIN => \N__11690\,
            DOUT => \N__11689\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11691\,
            PADOUT => \N__11690\,
            PADIN => \N__11689\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11682\,
            DIN => \N__11681\,
            DOUT => \N__11680\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11682\,
            PADOUT => \N__11681\,
            PADIN => \N__11680\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11673\,
            DIN => \N__11672\,
            DOUT => \N__11671\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11673\,
            PADOUT => \N__11672\,
            PADIN => \N__11671\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5088\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2838\ : InMux
    port map (
            O => \N__11654\,
            I => \N__11650\
        );

    \I__2837\ : InMux
    port map (
            O => \N__11653\,
            I => \N__11647\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__11650\,
            I => \N__11644\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__11647\,
            I => \N__11641\
        );

    \I__2834\ : Span12Mux_s9_h
    port map (
            O => \N__11644\,
            I => \N__11638\
        );

    \I__2833\ : Span4Mux_h
    port map (
            O => \N__11641\,
            I => \N__11635\
        );

    \I__2832\ : Span12Mux_h
    port map (
            O => \N__11638\,
            I => \N__11631\
        );

    \I__2831\ : Span4Mux_v
    port map (
            O => \N__11635\,
            I => \N__11628\
        );

    \I__2830\ : InMux
    port map (
            O => \N__11634\,
            I => \N__11625\
        );

    \I__2829\ : Odrv12
    port map (
            O => \N__11631\,
            I => \REG_CYCLEm\
        );

    \I__2828\ : Odrv4
    port map (
            O => \N__11628\,
            I => \REG_CYCLEm\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__11625\,
            I => \REG_CYCLEm\
        );

    \I__2826\ : IoInMux
    port map (
            O => \N__11618\,
            I => \N__11615\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__11615\,
            I => \N__11612\
        );

    \I__2824\ : Span4Mux_s2_v
    port map (
            O => \N__11612\,
            I => \N__11609\
        );

    \I__2823\ : Span4Mux_v
    port map (
            O => \N__11609\,
            I => \N__11606\
        );

    \I__2822\ : Odrv4
    port map (
            O => \N__11606\,
            I => \DRDENn_c\
        );

    \I__2821\ : InMux
    port map (
            O => \N__11603\,
            I => \N__11600\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__11600\,
            I => \N__11597\
        );

    \I__2819\ : Odrv12
    port map (
            O => \N__11597\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2818\ : InMux
    port map (
            O => \N__11594\,
            I => \N__11590\
        );

    \I__2817\ : InMux
    port map (
            O => \N__11593\,
            I => \N__11586\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__11590\,
            I => \N__11583\
        );

    \I__2815\ : InMux
    port map (
            O => \N__11589\,
            I => \N__11580\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__11586\,
            I => \N__11572\
        );

    \I__2813\ : Span4Mux_v
    port map (
            O => \N__11583\,
            I => \N__11572\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__11580\,
            I => \N__11572\
        );

    \I__2811\ : InMux
    port map (
            O => \N__11579\,
            I => \N__11569\
        );

    \I__2810\ : Span4Mux_h
    port map (
            O => \N__11572\,
            I => \N__11566\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__11569\,
            I => \N__11563\
        );

    \I__2808\ : Span4Mux_v
    port map (
            O => \N__11566\,
            I => \N__11560\
        );

    \I__2807\ : Sp12to4
    port map (
            O => \N__11563\,
            I => \N__11557\
        );

    \I__2806\ : Sp12to4
    port map (
            O => \N__11560\,
            I => \N__11552\
        );

    \I__2805\ : Span12Mux_v
    port map (
            O => \N__11557\,
            I => \N__11552\
        );

    \I__2804\ : Odrv12
    port map (
            O => \N__11552\,
            I => \DRA_c_2\
        );

    \I__2803\ : InMux
    port map (
            O => \N__11549\,
            I => \N__11543\
        );

    \I__2802\ : InMux
    port map (
            O => \N__11548\,
            I => \N__11543\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__11543\,
            I => \N__11540\
        );

    \I__2800\ : Span4Mux_h
    port map (
            O => \N__11540\,
            I => \N__11537\
        );

    \I__2799\ : Odrv4
    port map (
            O => \N__11537\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2798\ : InMux
    port map (
            O => \N__11534\,
            I => \N__11531\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__11531\,
            I => \N__11527\
        );

    \I__2796\ : InMux
    port map (
            O => \N__11530\,
            I => \N__11524\
        );

    \I__2795\ : Span4Mux_h
    port map (
            O => \N__11527\,
            I => \N__11517\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__11524\,
            I => \N__11517\
        );

    \I__2793\ : InMux
    port map (
            O => \N__11523\,
            I => \N__11514\
        );

    \I__2792\ : InMux
    port map (
            O => \N__11522\,
            I => \N__11511\
        );

    \I__2791\ : Span4Mux_h
    port map (
            O => \N__11517\,
            I => \N__11504\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__11514\,
            I => \N__11504\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__11511\,
            I => \N__11504\
        );

    \I__2788\ : Span4Mux_v
    port map (
            O => \N__11504\,
            I => \N__11501\
        );

    \I__2787\ : Span4Mux_v
    port map (
            O => \N__11501\,
            I => \N__11498\
        );

    \I__2786\ : Sp12to4
    port map (
            O => \N__11498\,
            I => \N__11495\
        );

    \I__2785\ : Odrv12
    port map (
            O => \N__11495\,
            I => \DRA_c_1\
        );

    \I__2784\ : InMux
    port map (
            O => \N__11492\,
            I => \N__11488\
        );

    \I__2783\ : InMux
    port map (
            O => \N__11491\,
            I => \N__11485\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__11488\,
            I => \N__11480\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__11485\,
            I => \N__11480\
        );

    \I__2780\ : Span4Mux_h
    port map (
            O => \N__11480\,
            I => \N__11477\
        );

    \I__2779\ : Sp12to4
    port map (
            O => \N__11477\,
            I => \N__11474\
        );

    \I__2778\ : Span12Mux_v
    port map (
            O => \N__11474\,
            I => \N__11471\
        );

    \I__2777\ : Odrv12
    port map (
            O => \N__11471\,
            I => \DRA_c_0\
        );

    \I__2776\ : InMux
    port map (
            O => \N__11468\,
            I => \N__11465\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__11465\,
            I => \N__11462\
        );

    \I__2774\ : Span4Mux_h
    port map (
            O => \N__11462\,
            I => \N__11459\
        );

    \I__2773\ : Odrv4
    port map (
            O => \N__11459\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2772\ : InMux
    port map (
            O => \N__11456\,
            I => \N__11452\
        );

    \I__2771\ : InMux
    port map (
            O => \N__11455\,
            I => \N__11448\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__11452\,
            I => \N__11444\
        );

    \I__2769\ : InMux
    port map (
            O => \N__11451\,
            I => \N__11441\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__11448\,
            I => \N__11438\
        );

    \I__2767\ : InMux
    port map (
            O => \N__11447\,
            I => \N__11435\
        );

    \I__2766\ : Span12Mux_v
    port map (
            O => \N__11444\,
            I => \N__11430\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__11441\,
            I => \N__11430\
        );

    \I__2764\ : Span4Mux_v
    port map (
            O => \N__11438\,
            I => \N__11427\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__11435\,
            I => \N__11424\
        );

    \I__2762\ : Span12Mux_h
    port map (
            O => \N__11430\,
            I => \N__11421\
        );

    \I__2761\ : Sp12to4
    port map (
            O => \N__11427\,
            I => \N__11416\
        );

    \I__2760\ : Span12Mux_v
    port map (
            O => \N__11424\,
            I => \N__11416\
        );

    \I__2759\ : Odrv12
    port map (
            O => \N__11421\,
            I => \DRA_c_8\
        );

    \I__2758\ : Odrv12
    port map (
            O => \N__11416\,
            I => \DRA_c_8\
        );

    \I__2757\ : InMux
    port map (
            O => \N__11411\,
            I => \N__11408\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__11408\,
            I => \N__11405\
        );

    \I__2755\ : Odrv4
    port map (
            O => \N__11405\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2754\ : InMux
    port map (
            O => \N__11402\,
            I => \N__11399\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__11399\,
            I => \N__11396\
        );

    \I__2752\ : Span4Mux_v
    port map (
            O => \N__11396\,
            I => \N__11390\
        );

    \I__2751\ : InMux
    port map (
            O => \N__11395\,
            I => \N__11387\
        );

    \I__2750\ : InMux
    port map (
            O => \N__11394\,
            I => \N__11382\
        );

    \I__2749\ : InMux
    port map (
            O => \N__11393\,
            I => \N__11382\
        );

    \I__2748\ : Span4Mux_h
    port map (
            O => \N__11390\,
            I => \N__11379\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__11387\,
            I => \N__11374\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__11382\,
            I => \N__11374\
        );

    \I__2745\ : Sp12to4
    port map (
            O => \N__11379\,
            I => \N__11369\
        );

    \I__2744\ : Span12Mux_h
    port map (
            O => \N__11374\,
            I => \N__11369\
        );

    \I__2743\ : Odrv12
    port map (
            O => \N__11369\,
            I => \DRA_c_7\
        );

    \I__2742\ : InMux
    port map (
            O => \N__11366\,
            I => \N__11362\
        );

    \I__2741\ : InMux
    port map (
            O => \N__11365\,
            I => \N__11359\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__11362\,
            I => \N__11353\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__11359\,
            I => \N__11353\
        );

    \I__2738\ : InMux
    port map (
            O => \N__11358\,
            I => \N__11349\
        );

    \I__2737\ : Span4Mux_v
    port map (
            O => \N__11353\,
            I => \N__11346\
        );

    \I__2736\ : InMux
    port map (
            O => \N__11352\,
            I => \N__11343\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__11349\,
            I => \N__11340\
        );

    \I__2734\ : Sp12to4
    port map (
            O => \N__11346\,
            I => \N__11337\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__11343\,
            I => \N__11334\
        );

    \I__2732\ : Span4Mux_v
    port map (
            O => \N__11340\,
            I => \N__11331\
        );

    \I__2731\ : Span12Mux_h
    port map (
            O => \N__11337\,
            I => \N__11328\
        );

    \I__2730\ : Span12Mux_v
    port map (
            O => \N__11334\,
            I => \N__11323\
        );

    \I__2729\ : Sp12to4
    port map (
            O => \N__11331\,
            I => \N__11323\
        );

    \I__2728\ : Odrv12
    port map (
            O => \N__11328\,
            I => \DRA_c_6\
        );

    \I__2727\ : Odrv12
    port map (
            O => \N__11323\,
            I => \DRA_c_6\
        );

    \I__2726\ : InMux
    port map (
            O => \N__11318\,
            I => \N__11315\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__11315\,
            I => \N__11312\
        );

    \I__2724\ : Odrv4
    port map (
            O => \N__11312\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2723\ : InMux
    port map (
            O => \N__11309\,
            I => \N__11306\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__11306\,
            I => \N__11303\
        );

    \I__2721\ : Span12Mux_v
    port map (
            O => \N__11303\,
            I => \N__11300\
        );

    \I__2720\ : Odrv12
    port map (
            O => \N__11300\,
            I => \RAS0n_c\
        );

    \I__2719\ : InMux
    port map (
            O => \N__11297\,
            I => \N__11294\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__11294\,
            I => \N__11276\
        );

    \I__2717\ : InMux
    port map (
            O => \N__11293\,
            I => \N__11269\
        );

    \I__2716\ : InMux
    port map (
            O => \N__11292\,
            I => \N__11269\
        );

    \I__2715\ : InMux
    port map (
            O => \N__11291\,
            I => \N__11262\
        );

    \I__2714\ : InMux
    port map (
            O => \N__11290\,
            I => \N__11262\
        );

    \I__2713\ : InMux
    port map (
            O => \N__11289\,
            I => \N__11262\
        );

    \I__2712\ : InMux
    port map (
            O => \N__11288\,
            I => \N__11259\
        );

    \I__2711\ : InMux
    port map (
            O => \N__11287\,
            I => \N__11256\
        );

    \I__2710\ : InMux
    port map (
            O => \N__11286\,
            I => \N__11253\
        );

    \I__2709\ : InMux
    port map (
            O => \N__11285\,
            I => \N__11250\
        );

    \I__2708\ : InMux
    port map (
            O => \N__11284\,
            I => \N__11247\
        );

    \I__2707\ : InMux
    port map (
            O => \N__11283\,
            I => \N__11244\
        );

    \I__2706\ : InMux
    port map (
            O => \N__11282\,
            I => \N__11241\
        );

    \I__2705\ : InMux
    port map (
            O => \N__11281\,
            I => \N__11238\
        );

    \I__2704\ : InMux
    port map (
            O => \N__11280\,
            I => \N__11235\
        );

    \I__2703\ : InMux
    port map (
            O => \N__11279\,
            I => \N__11230\
        );

    \I__2702\ : Span4Mux_v
    port map (
            O => \N__11276\,
            I => \N__11226\
        );

    \I__2701\ : InMux
    port map (
            O => \N__11275\,
            I => \N__11223\
        );

    \I__2700\ : InMux
    port map (
            O => \N__11274\,
            I => \N__11220\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__11269\,
            I => \N__11217\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__11262\,
            I => \N__11210\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__11259\,
            I => \N__11210\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__11256\,
            I => \N__11210\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__11253\,
            I => \N__11207\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__11250\,
            I => \N__11194\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__11247\,
            I => \N__11194\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__11244\,
            I => \N__11194\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__11241\,
            I => \N__11194\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__11238\,
            I => \N__11194\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__11235\,
            I => \N__11194\
        );

    \I__2688\ : InMux
    port map (
            O => \N__11234\,
            I => \N__11191\
        );

    \I__2687\ : InMux
    port map (
            O => \N__11233\,
            I => \N__11188\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__11230\,
            I => \N__11185\
        );

    \I__2685\ : InMux
    port map (
            O => \N__11229\,
            I => \N__11182\
        );

    \I__2684\ : Span4Mux_h
    port map (
            O => \N__11226\,
            I => \N__11171\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__11223\,
            I => \N__11171\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__11220\,
            I => \N__11171\
        );

    \I__2681\ : Span4Mux_v
    port map (
            O => \N__11217\,
            I => \N__11171\
        );

    \I__2680\ : Span4Mux_v
    port map (
            O => \N__11210\,
            I => \N__11171\
        );

    \I__2679\ : Span4Mux_v
    port map (
            O => \N__11207\,
            I => \N__11166\
        );

    \I__2678\ : Span4Mux_v
    port map (
            O => \N__11194\,
            I => \N__11166\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__11191\,
            I => \N__11161\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__11188\,
            I => \N__11161\
        );

    \I__2675\ : Span4Mux_h
    port map (
            O => \N__11185\,
            I => \N__11158\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__11182\,
            I => \N__11151\
        );

    \I__2673\ : Sp12to4
    port map (
            O => \N__11171\,
            I => \N__11151\
        );

    \I__2672\ : Sp12to4
    port map (
            O => \N__11166\,
            I => \N__11151\
        );

    \I__2671\ : Span12Mux_v
    port map (
            O => \N__11161\,
            I => \N__11148\
        );

    \I__2670\ : Sp12to4
    port map (
            O => \N__11158\,
            I => \N__11143\
        );

    \I__2669\ : Span12Mux_h
    port map (
            O => \N__11151\,
            I => \N__11143\
        );

    \I__2668\ : Span12Mux_h
    port map (
            O => \N__11148\,
            I => \N__11140\
        );

    \I__2667\ : Span12Mux_v
    port map (
            O => \N__11143\,
            I => \N__11137\
        );

    \I__2666\ : Odrv12
    port map (
            O => \N__11140\,
            I => \AGNUS_REV_c\
        );

    \I__2665\ : Odrv12
    port map (
            O => \N__11137\,
            I => \AGNUS_REV_c\
        );

    \I__2664\ : InMux
    port map (
            O => \N__11132\,
            I => \N__11128\
        );

    \I__2663\ : InMux
    port map (
            O => \N__11131\,
            I => \N__11125\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__11128\,
            I => \N__11118\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__11125\,
            I => \N__11118\
        );

    \I__2660\ : InMux
    port map (
            O => \N__11124\,
            I => \N__11115\
        );

    \I__2659\ : InMux
    port map (
            O => \N__11123\,
            I => \N__11112\
        );

    \I__2658\ : Span12Mux_v
    port map (
            O => \N__11118\,
            I => \N__11109\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__11115\,
            I => \N__11106\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__11112\,
            I => \N__11103\
        );

    \I__2655\ : Span12Mux_h
    port map (
            O => \N__11109\,
            I => \N__11100\
        );

    \I__2654\ : Span12Mux_v
    port map (
            O => \N__11106\,
            I => \N__11097\
        );

    \I__2653\ : Span12Mux_v
    port map (
            O => \N__11103\,
            I => \N__11094\
        );

    \I__2652\ : Span12Mux_v
    port map (
            O => \N__11100\,
            I => \N__11089\
        );

    \I__2651\ : Span12Mux_h
    port map (
            O => \N__11097\,
            I => \N__11089\
        );

    \I__2650\ : Span12Mux_v
    port map (
            O => \N__11094\,
            I => \N__11086\
        );

    \I__2649\ : Odrv12
    port map (
            O => \N__11089\,
            I => \DRA_c_9\
        );

    \I__2648\ : Odrv12
    port map (
            O => \N__11086\,
            I => \DRA_c_9\
        );

    \I__2647\ : InMux
    port map (
            O => \N__11081\,
            I => \N__11078\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__11078\,
            I => \N__11075\
        );

    \I__2645\ : Span12Mux_v
    port map (
            O => \N__11075\,
            I => \N__11072\
        );

    \I__2644\ : Odrv12
    port map (
            O => \N__11072\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2643\ : ClkMux
    port map (
            O => \N__11069\,
            I => \N__11042\
        );

    \I__2642\ : ClkMux
    port map (
            O => \N__11068\,
            I => \N__11042\
        );

    \I__2641\ : ClkMux
    port map (
            O => \N__11067\,
            I => \N__11042\
        );

    \I__2640\ : ClkMux
    port map (
            O => \N__11066\,
            I => \N__11042\
        );

    \I__2639\ : ClkMux
    port map (
            O => \N__11065\,
            I => \N__11042\
        );

    \I__2638\ : ClkMux
    port map (
            O => \N__11064\,
            I => \N__11042\
        );

    \I__2637\ : ClkMux
    port map (
            O => \N__11063\,
            I => \N__11042\
        );

    \I__2636\ : ClkMux
    port map (
            O => \N__11062\,
            I => \N__11042\
        );

    \I__2635\ : ClkMux
    port map (
            O => \N__11061\,
            I => \N__11042\
        );

    \I__2634\ : GlobalMux
    port map (
            O => \N__11042\,
            I => \N__11039\
        );

    \I__2633\ : gio2CtrlBuf
    port map (
            O => \N__11039\,
            I => \C3_c_g\
        );

    \I__2632\ : CEMux
    port map (
            O => \N__11036\,
            I => \N__10988\
        );

    \I__2631\ : CEMux
    port map (
            O => \N__11035\,
            I => \N__10988\
        );

    \I__2630\ : CEMux
    port map (
            O => \N__11034\,
            I => \N__10988\
        );

    \I__2629\ : CEMux
    port map (
            O => \N__11033\,
            I => \N__10988\
        );

    \I__2628\ : CEMux
    port map (
            O => \N__11032\,
            I => \N__10988\
        );

    \I__2627\ : CEMux
    port map (
            O => \N__11031\,
            I => \N__10988\
        );

    \I__2626\ : CEMux
    port map (
            O => \N__11030\,
            I => \N__10988\
        );

    \I__2625\ : CEMux
    port map (
            O => \N__11029\,
            I => \N__10988\
        );

    \I__2624\ : CEMux
    port map (
            O => \N__11028\,
            I => \N__10988\
        );

    \I__2623\ : CEMux
    port map (
            O => \N__11027\,
            I => \N__10988\
        );

    \I__2622\ : CEMux
    port map (
            O => \N__11026\,
            I => \N__10988\
        );

    \I__2621\ : CEMux
    port map (
            O => \N__11025\,
            I => \N__10988\
        );

    \I__2620\ : CEMux
    port map (
            O => \N__11024\,
            I => \N__10988\
        );

    \I__2619\ : CEMux
    port map (
            O => \N__11023\,
            I => \N__10988\
        );

    \I__2618\ : CEMux
    port map (
            O => \N__11022\,
            I => \N__10988\
        );

    \I__2617\ : CEMux
    port map (
            O => \N__11021\,
            I => \N__10988\
        );

    \I__2616\ : GlobalMux
    port map (
            O => \N__10988\,
            I => \N__10985\
        );

    \I__2615\ : gio2CtrlBuf
    port map (
            O => \N__10985\,
            I => \DBRn_c_i_0_g\
        );

    \I__2614\ : InMux
    port map (
            O => \N__10982\,
            I => \N__10976\
        );

    \I__2613\ : InMux
    port map (
            O => \N__10981\,
            I => \N__10973\
        );

    \I__2612\ : InMux
    port map (
            O => \N__10980\,
            I => \N__10970\
        );

    \I__2611\ : InMux
    port map (
            O => \N__10979\,
            I => \N__10967\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__10976\,
            I => \N__10959\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__10973\,
            I => \N__10935\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__10970\,
            I => \N__10919\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__10967\,
            I => \N__10914\
        );

    \I__2606\ : SRMux
    port map (
            O => \N__10966\,
            I => \N__10820\
        );

    \I__2605\ : SRMux
    port map (
            O => \N__10965\,
            I => \N__10820\
        );

    \I__2604\ : SRMux
    port map (
            O => \N__10964\,
            I => \N__10820\
        );

    \I__2603\ : SRMux
    port map (
            O => \N__10963\,
            I => \N__10820\
        );

    \I__2602\ : SRMux
    port map (
            O => \N__10962\,
            I => \N__10820\
        );

    \I__2601\ : Glb2LocalMux
    port map (
            O => \N__10959\,
            I => \N__10820\
        );

    \I__2600\ : SRMux
    port map (
            O => \N__10958\,
            I => \N__10820\
        );

    \I__2599\ : SRMux
    port map (
            O => \N__10957\,
            I => \N__10820\
        );

    \I__2598\ : SRMux
    port map (
            O => \N__10956\,
            I => \N__10820\
        );

    \I__2597\ : SRMux
    port map (
            O => \N__10955\,
            I => \N__10820\
        );

    \I__2596\ : SRMux
    port map (
            O => \N__10954\,
            I => \N__10820\
        );

    \I__2595\ : SRMux
    port map (
            O => \N__10953\,
            I => \N__10820\
        );

    \I__2594\ : SRMux
    port map (
            O => \N__10952\,
            I => \N__10820\
        );

    \I__2593\ : SRMux
    port map (
            O => \N__10951\,
            I => \N__10820\
        );

    \I__2592\ : SRMux
    port map (
            O => \N__10950\,
            I => \N__10820\
        );

    \I__2591\ : SRMux
    port map (
            O => \N__10949\,
            I => \N__10820\
        );

    \I__2590\ : SRMux
    port map (
            O => \N__10948\,
            I => \N__10820\
        );

    \I__2589\ : SRMux
    port map (
            O => \N__10947\,
            I => \N__10820\
        );

    \I__2588\ : SRMux
    port map (
            O => \N__10946\,
            I => \N__10820\
        );

    \I__2587\ : SRMux
    port map (
            O => \N__10945\,
            I => \N__10820\
        );

    \I__2586\ : SRMux
    port map (
            O => \N__10944\,
            I => \N__10820\
        );

    \I__2585\ : SRMux
    port map (
            O => \N__10943\,
            I => \N__10820\
        );

    \I__2584\ : SRMux
    port map (
            O => \N__10942\,
            I => \N__10820\
        );

    \I__2583\ : SRMux
    port map (
            O => \N__10941\,
            I => \N__10820\
        );

    \I__2582\ : SRMux
    port map (
            O => \N__10940\,
            I => \N__10820\
        );

    \I__2581\ : SRMux
    port map (
            O => \N__10939\,
            I => \N__10820\
        );

    \I__2580\ : SRMux
    port map (
            O => \N__10938\,
            I => \N__10820\
        );

    \I__2579\ : Glb2LocalMux
    port map (
            O => \N__10935\,
            I => \N__10820\
        );

    \I__2578\ : SRMux
    port map (
            O => \N__10934\,
            I => \N__10820\
        );

    \I__2577\ : SRMux
    port map (
            O => \N__10933\,
            I => \N__10820\
        );

    \I__2576\ : SRMux
    port map (
            O => \N__10932\,
            I => \N__10820\
        );

    \I__2575\ : SRMux
    port map (
            O => \N__10931\,
            I => \N__10820\
        );

    \I__2574\ : SRMux
    port map (
            O => \N__10930\,
            I => \N__10820\
        );

    \I__2573\ : SRMux
    port map (
            O => \N__10929\,
            I => \N__10820\
        );

    \I__2572\ : SRMux
    port map (
            O => \N__10928\,
            I => \N__10820\
        );

    \I__2571\ : SRMux
    port map (
            O => \N__10927\,
            I => \N__10820\
        );

    \I__2570\ : SRMux
    port map (
            O => \N__10926\,
            I => \N__10820\
        );

    \I__2569\ : SRMux
    port map (
            O => \N__10925\,
            I => \N__10820\
        );

    \I__2568\ : SRMux
    port map (
            O => \N__10924\,
            I => \N__10820\
        );

    \I__2567\ : SRMux
    port map (
            O => \N__10923\,
            I => \N__10820\
        );

    \I__2566\ : SRMux
    port map (
            O => \N__10922\,
            I => \N__10820\
        );

    \I__2565\ : Glb2LocalMux
    port map (
            O => \N__10919\,
            I => \N__10820\
        );

    \I__2564\ : SRMux
    port map (
            O => \N__10918\,
            I => \N__10820\
        );

    \I__2563\ : SRMux
    port map (
            O => \N__10917\,
            I => \N__10820\
        );

    \I__2562\ : Glb2LocalMux
    port map (
            O => \N__10914\,
            I => \N__10820\
        );

    \I__2561\ : SRMux
    port map (
            O => \N__10913\,
            I => \N__10820\
        );

    \I__2560\ : GlobalMux
    port map (
            O => \N__10820\,
            I => \N__10817\
        );

    \I__2559\ : gio2CtrlBuf
    port map (
            O => \N__10817\,
            I => \RESETn_c_i_g\
        );

    \I__2558\ : InMux
    port map (
            O => \N__10814\,
            I => \N__10810\
        );

    \I__2557\ : InMux
    port map (
            O => \N__10813\,
            I => \N__10807\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__10810\,
            I => \N__10802\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__10807\,
            I => \N__10798\
        );

    \I__2554\ : InMux
    port map (
            O => \N__10806\,
            I => \N__10795\
        );

    \I__2553\ : InMux
    port map (
            O => \N__10805\,
            I => \N__10792\
        );

    \I__2552\ : Span4Mux_v
    port map (
            O => \N__10802\,
            I => \N__10789\
        );

    \I__2551\ : InMux
    port map (
            O => \N__10801\,
            I => \N__10786\
        );

    \I__2550\ : Span4Mux_v
    port map (
            O => \N__10798\,
            I => \N__10781\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__10795\,
            I => \N__10781\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__10792\,
            I => \N__10778\
        );

    \I__2547\ : Sp12to4
    port map (
            O => \N__10789\,
            I => \N__10775\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__10786\,
            I => \N__10772\
        );

    \I__2545\ : Span4Mux_v
    port map (
            O => \N__10781\,
            I => \N__10769\
        );

    \I__2544\ : Span4Mux_v
    port map (
            O => \N__10778\,
            I => \N__10766\
        );

    \I__2543\ : Span12Mux_h
    port map (
            O => \N__10775\,
            I => \N__10761\
        );

    \I__2542\ : Span12Mux_v
    port map (
            O => \N__10772\,
            I => \N__10761\
        );

    \I__2541\ : Sp12to4
    port map (
            O => \N__10769\,
            I => \N__10756\
        );

    \I__2540\ : Sp12to4
    port map (
            O => \N__10766\,
            I => \N__10756\
        );

    \I__2539\ : Span12Mux_h
    port map (
            O => \N__10761\,
            I => \N__10753\
        );

    \I__2538\ : Span12Mux_h
    port map (
            O => \N__10756\,
            I => \N__10750\
        );

    \I__2537\ : Odrv12
    port map (
            O => \N__10753\,
            I => \RnW_c\
        );

    \I__2536\ : Odrv12
    port map (
            O => \N__10750\,
            I => \RnW_c\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__10745\,
            I => \N__10742\
        );

    \I__2534\ : InMux
    port map (
            O => \N__10742\,
            I => \N__10739\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__10739\,
            I => \N__10735\
        );

    \I__2532\ : InMux
    port map (
            O => \N__10738\,
            I => \N__10732\
        );

    \I__2531\ : Span12Mux_s10_v
    port map (
            O => \N__10735\,
            I => \N__10729\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__10732\,
            I => \N__10726\
        );

    \I__2529\ : Span12Mux_h
    port map (
            O => \N__10729\,
            I => \N__10717\
        );

    \I__2528\ : Span12Mux_v
    port map (
            O => \N__10726\,
            I => \N__10714\
        );

    \I__2527\ : InMux
    port map (
            O => \N__10725\,
            I => \N__10711\
        );

    \I__2526\ : InMux
    port map (
            O => \N__10724\,
            I => \N__10708\
        );

    \I__2525\ : InMux
    port map (
            O => \N__10723\,
            I => \N__10705\
        );

    \I__2524\ : InMux
    port map (
            O => \N__10722\,
            I => \N__10700\
        );

    \I__2523\ : InMux
    port map (
            O => \N__10721\,
            I => \N__10700\
        );

    \I__2522\ : InMux
    port map (
            O => \N__10720\,
            I => \N__10697\
        );

    \I__2521\ : Odrv12
    port map (
            O => \N__10717\,
            I => \WRITE_CYCLEm\
        );

    \I__2520\ : Odrv12
    port map (
            O => \N__10714\,
            I => \WRITE_CYCLEm\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__10711\,
            I => \WRITE_CYCLEm\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__10708\,
            I => \WRITE_CYCLEm\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__10705\,
            I => \WRITE_CYCLEm\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__10700\,
            I => \WRITE_CYCLEm\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__10697\,
            I => \WRITE_CYCLEm\
        );

    \I__2514\ : IoInMux
    port map (
            O => \N__10682\,
            I => \N__10679\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__10679\,
            I => \N__10676\
        );

    \I__2512\ : Span4Mux_s3_h
    port map (
            O => \N__10676\,
            I => \N__10673\
        );

    \I__2511\ : Span4Mux_v
    port map (
            O => \N__10673\,
            I => \N__10670\
        );

    \I__2510\ : Odrv4
    port map (
            O => \N__10670\,
            I => \DRDDIR_c\
        );

    \I__2509\ : InMux
    port map (
            O => \N__10667\,
            I => \N__10662\
        );

    \I__2508\ : InMux
    port map (
            O => \N__10666\,
            I => \N__10656\
        );

    \I__2507\ : InMux
    port map (
            O => \N__10665\,
            I => \N__10656\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__10662\,
            I => \N__10653\
        );

    \I__2505\ : InMux
    port map (
            O => \N__10661\,
            I => \N__10650\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__10656\,
            I => \N__10647\
        );

    \I__2503\ : Span4Mux_v
    port map (
            O => \N__10653\,
            I => \N__10644\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__10650\,
            I => \N__10641\
        );

    \I__2501\ : Span4Mux_v
    port map (
            O => \N__10647\,
            I => \N__10638\
        );

    \I__2500\ : Sp12to4
    port map (
            O => \N__10644\,
            I => \N__10633\
        );

    \I__2499\ : Sp12to4
    port map (
            O => \N__10641\,
            I => \N__10630\
        );

    \I__2498\ : Sp12to4
    port map (
            O => \N__10638\,
            I => \N__10627\
        );

    \I__2497\ : InMux
    port map (
            O => \N__10637\,
            I => \N__10622\
        );

    \I__2496\ : InMux
    port map (
            O => \N__10636\,
            I => \N__10622\
        );

    \I__2495\ : Span12Mux_h
    port map (
            O => \N__10633\,
            I => \N__10619\
        );

    \I__2494\ : Span12Mux_v
    port map (
            O => \N__10630\,
            I => \N__10616\
        );

    \I__2493\ : Span12Mux_h
    port map (
            O => \N__10627\,
            I => \N__10611\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__10622\,
            I => \N__10611\
        );

    \I__2491\ : Span12Mux_v
    port map (
            O => \N__10619\,
            I => \N__10608\
        );

    \I__2490\ : Span12Mux_h
    port map (
            O => \N__10616\,
            I => \N__10603\
        );

    \I__2489\ : Span12Mux_v
    port map (
            O => \N__10611\,
            I => \N__10603\
        );

    \I__2488\ : Odrv12
    port map (
            O => \N__10608\,
            I => \CASLn_c\
        );

    \I__2487\ : Odrv12
    port map (
            O => \N__10603\,
            I => \CASLn_c\
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__10598\,
            I => \N__10595\
        );

    \I__2485\ : InMux
    port map (
            O => \N__10595\,
            I => \N__10592\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__10592\,
            I => \N__10589\
        );

    \I__2483\ : Span4Mux_v
    port map (
            O => \N__10589\,
            I => \N__10585\
        );

    \I__2482\ : InMux
    port map (
            O => \N__10588\,
            I => \N__10581\
        );

    \I__2481\ : Span4Mux_v
    port map (
            O => \N__10585\,
            I => \N__10577\
        );

    \I__2480\ : InMux
    port map (
            O => \N__10584\,
            I => \N__10574\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__10581\,
            I => \N__10570\
        );

    \I__2478\ : InMux
    port map (
            O => \N__10580\,
            I => \N__10567\
        );

    \I__2477\ : Span4Mux_v
    port map (
            O => \N__10577\,
            I => \N__10562\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__10574\,
            I => \N__10562\
        );

    \I__2475\ : CascadeMux
    port map (
            O => \N__10573\,
            I => \N__10559\
        );

    \I__2474\ : Sp12to4
    port map (
            O => \N__10570\,
            I => \N__10555\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__10567\,
            I => \N__10552\
        );

    \I__2472\ : Span4Mux_v
    port map (
            O => \N__10562\,
            I => \N__10549\
        );

    \I__2471\ : InMux
    port map (
            O => \N__10559\,
            I => \N__10544\
        );

    \I__2470\ : InMux
    port map (
            O => \N__10558\,
            I => \N__10544\
        );

    \I__2469\ : Span12Mux_v
    port map (
            O => \N__10555\,
            I => \N__10541\
        );

    \I__2468\ : Span12Mux_h
    port map (
            O => \N__10552\,
            I => \N__10538\
        );

    \I__2467\ : Sp12to4
    port map (
            O => \N__10549\,
            I => \N__10535\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__10544\,
            I => \N__10532\
        );

    \I__2465\ : Span12Mux_h
    port map (
            O => \N__10541\,
            I => \N__10529\
        );

    \I__2464\ : Span12Mux_v
    port map (
            O => \N__10538\,
            I => \N__10524\
        );

    \I__2463\ : Span12Mux_h
    port map (
            O => \N__10535\,
            I => \N__10524\
        );

    \I__2462\ : Span4Mux_v
    port map (
            O => \N__10532\,
            I => \N__10521\
        );

    \I__2461\ : Odrv12
    port map (
            O => \N__10529\,
            I => \CASUn_c\
        );

    \I__2460\ : Odrv12
    port map (
            O => \N__10524\,
            I => \CASUn_c\
        );

    \I__2459\ : Odrv4
    port map (
            O => \N__10521\,
            I => \CASUn_c\
        );

    \I__2458\ : InMux
    port map (
            O => \N__10514\,
            I => \N__10511\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__10511\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__2456\ : IoInMux
    port map (
            O => \N__10508\,
            I => \N__10505\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__10505\,
            I => \N__10502\
        );

    \I__2454\ : Span12Mux_s4_h
    port map (
            O => \N__10502\,
            I => \N__10499\
        );

    \I__2453\ : Span12Mux_v
    port map (
            O => \N__10499\,
            I => \N__10496\
        );

    \I__2452\ : Odrv12
    port map (
            O => \N__10496\,
            I => \CMA_c_6\
        );

    \I__2451\ : InMux
    port map (
            O => \N__10493\,
            I => \N__10490\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__10490\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__2449\ : IoInMux
    port map (
            O => \N__10487\,
            I => \N__10484\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__10484\,
            I => \N__10481\
        );

    \I__2447\ : IoSpan4Mux
    port map (
            O => \N__10481\,
            I => \N__10478\
        );

    \I__2446\ : Span4Mux_s0_h
    port map (
            O => \N__10478\,
            I => \N__10475\
        );

    \I__2445\ : Sp12to4
    port map (
            O => \N__10475\,
            I => \N__10472\
        );

    \I__2444\ : Span12Mux_v
    port map (
            O => \N__10472\,
            I => \N__10469\
        );

    \I__2443\ : Odrv12
    port map (
            O => \N__10469\,
            I => \CMA_c_4\
        );

    \I__2442\ : InMux
    port map (
            O => \N__10466\,
            I => \N__10457\
        );

    \I__2441\ : InMux
    port map (
            O => \N__10465\,
            I => \N__10457\
        );

    \I__2440\ : InMux
    port map (
            O => \N__10464\,
            I => \N__10457\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__10457\,
            I => \N__10451\
        );

    \I__2438\ : InMux
    port map (
            O => \N__10456\,
            I => \N__10444\
        );

    \I__2437\ : InMux
    port map (
            O => \N__10455\,
            I => \N__10444\
        );

    \I__2436\ : InMux
    port map (
            O => \N__10454\,
            I => \N__10444\
        );

    \I__2435\ : Odrv4
    port map (
            O => \N__10451\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__10444\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\
        );

    \I__2433\ : CascadeMux
    port map (
            O => \N__10439\,
            I => \N__10432\
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__10438\,
            I => \N__10429\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__10437\,
            I => \N__10426\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__10436\,
            I => \N__10422\
        );

    \I__2429\ : CascadeMux
    port map (
            O => \N__10435\,
            I => \N__10419\
        );

    \I__2428\ : InMux
    port map (
            O => \N__10432\,
            I => \N__10412\
        );

    \I__2427\ : InMux
    port map (
            O => \N__10429\,
            I => \N__10412\
        );

    \I__2426\ : InMux
    port map (
            O => \N__10426\,
            I => \N__10412\
        );

    \I__2425\ : InMux
    port map (
            O => \N__10425\,
            I => \N__10408\
        );

    \I__2424\ : InMux
    port map (
            O => \N__10422\,
            I => \N__10403\
        );

    \I__2423\ : InMux
    port map (
            O => \N__10419\,
            I => \N__10403\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__10412\,
            I => \N__10400\
        );

    \I__2421\ : CascadeMux
    port map (
            O => \N__10411\,
            I => \N__10395\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__10408\,
            I => \N__10390\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__10403\,
            I => \N__10390\
        );

    \I__2418\ : Span4Mux_h
    port map (
            O => \N__10400\,
            I => \N__10387\
        );

    \I__2417\ : InMux
    port map (
            O => \N__10399\,
            I => \N__10384\
        );

    \I__2416\ : InMux
    port map (
            O => \N__10398\,
            I => \N__10379\
        );

    \I__2415\ : InMux
    port map (
            O => \N__10395\,
            I => \N__10379\
        );

    \I__2414\ : Odrv12
    port map (
            O => \N__10390\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2413\ : Odrv4
    port map (
            O => \N__10387\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__10384\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__10379\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2410\ : InMux
    port map (
            O => \N__10370\,
            I => \N__10367\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__10367\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__2408\ : IoInMux
    port map (
            O => \N__10364\,
            I => \N__10361\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__10361\,
            I => \N__10358\
        );

    \I__2406\ : IoSpan4Mux
    port map (
            O => \N__10358\,
            I => \N__10355\
        );

    \I__2405\ : Span4Mux_s2_h
    port map (
            O => \N__10355\,
            I => \N__10352\
        );

    \I__2404\ : Sp12to4
    port map (
            O => \N__10352\,
            I => \N__10349\
        );

    \I__2403\ : Span12Mux_v
    port map (
            O => \N__10349\,
            I => \N__10346\
        );

    \I__2402\ : Odrv12
    port map (
            O => \N__10346\,
            I => \CMA_c_7\
        );

    \I__2401\ : InMux
    port map (
            O => \N__10343\,
            I => \N__10340\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__10340\,
            I => \N__10301\
        );

    \I__2399\ : ClkMux
    port map (
            O => \N__10339\,
            I => \N__10202\
        );

    \I__2398\ : ClkMux
    port map (
            O => \N__10338\,
            I => \N__10202\
        );

    \I__2397\ : ClkMux
    port map (
            O => \N__10337\,
            I => \N__10202\
        );

    \I__2396\ : ClkMux
    port map (
            O => \N__10336\,
            I => \N__10202\
        );

    \I__2395\ : ClkMux
    port map (
            O => \N__10335\,
            I => \N__10202\
        );

    \I__2394\ : ClkMux
    port map (
            O => \N__10334\,
            I => \N__10202\
        );

    \I__2393\ : ClkMux
    port map (
            O => \N__10333\,
            I => \N__10202\
        );

    \I__2392\ : ClkMux
    port map (
            O => \N__10332\,
            I => \N__10202\
        );

    \I__2391\ : ClkMux
    port map (
            O => \N__10331\,
            I => \N__10202\
        );

    \I__2390\ : ClkMux
    port map (
            O => \N__10330\,
            I => \N__10202\
        );

    \I__2389\ : ClkMux
    port map (
            O => \N__10329\,
            I => \N__10202\
        );

    \I__2388\ : ClkMux
    port map (
            O => \N__10328\,
            I => \N__10202\
        );

    \I__2387\ : ClkMux
    port map (
            O => \N__10327\,
            I => \N__10202\
        );

    \I__2386\ : ClkMux
    port map (
            O => \N__10326\,
            I => \N__10202\
        );

    \I__2385\ : ClkMux
    port map (
            O => \N__10325\,
            I => \N__10202\
        );

    \I__2384\ : ClkMux
    port map (
            O => \N__10324\,
            I => \N__10202\
        );

    \I__2383\ : ClkMux
    port map (
            O => \N__10323\,
            I => \N__10202\
        );

    \I__2382\ : ClkMux
    port map (
            O => \N__10322\,
            I => \N__10202\
        );

    \I__2381\ : ClkMux
    port map (
            O => \N__10321\,
            I => \N__10202\
        );

    \I__2380\ : ClkMux
    port map (
            O => \N__10320\,
            I => \N__10202\
        );

    \I__2379\ : ClkMux
    port map (
            O => \N__10319\,
            I => \N__10202\
        );

    \I__2378\ : ClkMux
    port map (
            O => \N__10318\,
            I => \N__10202\
        );

    \I__2377\ : ClkMux
    port map (
            O => \N__10317\,
            I => \N__10202\
        );

    \I__2376\ : ClkMux
    port map (
            O => \N__10316\,
            I => \N__10202\
        );

    \I__2375\ : ClkMux
    port map (
            O => \N__10315\,
            I => \N__10202\
        );

    \I__2374\ : ClkMux
    port map (
            O => \N__10314\,
            I => \N__10202\
        );

    \I__2373\ : ClkMux
    port map (
            O => \N__10313\,
            I => \N__10202\
        );

    \I__2372\ : ClkMux
    port map (
            O => \N__10312\,
            I => \N__10202\
        );

    \I__2371\ : ClkMux
    port map (
            O => \N__10311\,
            I => \N__10202\
        );

    \I__2370\ : ClkMux
    port map (
            O => \N__10310\,
            I => \N__10202\
        );

    \I__2369\ : ClkMux
    port map (
            O => \N__10309\,
            I => \N__10202\
        );

    \I__2368\ : ClkMux
    port map (
            O => \N__10308\,
            I => \N__10202\
        );

    \I__2367\ : ClkMux
    port map (
            O => \N__10307\,
            I => \N__10202\
        );

    \I__2366\ : ClkMux
    port map (
            O => \N__10306\,
            I => \N__10202\
        );

    \I__2365\ : ClkMux
    port map (
            O => \N__10305\,
            I => \N__10202\
        );

    \I__2364\ : ClkMux
    port map (
            O => \N__10304\,
            I => \N__10202\
        );

    \I__2363\ : Glb2LocalMux
    port map (
            O => \N__10301\,
            I => \N__10202\
        );

    \I__2362\ : ClkMux
    port map (
            O => \N__10300\,
            I => \N__10202\
        );

    \I__2361\ : ClkMux
    port map (
            O => \N__10299\,
            I => \N__10202\
        );

    \I__2360\ : ClkMux
    port map (
            O => \N__10298\,
            I => \N__10202\
        );

    \I__2359\ : ClkMux
    port map (
            O => \N__10297\,
            I => \N__10202\
        );

    \I__2358\ : ClkMux
    port map (
            O => \N__10296\,
            I => \N__10202\
        );

    \I__2357\ : ClkMux
    port map (
            O => \N__10295\,
            I => \N__10202\
        );

    \I__2356\ : ClkMux
    port map (
            O => \N__10294\,
            I => \N__10202\
        );

    \I__2355\ : ClkMux
    port map (
            O => \N__10293\,
            I => \N__10202\
        );

    \I__2354\ : GlobalMux
    port map (
            O => \N__10202\,
            I => \CLK80_PLL\
        );

    \I__2353\ : CEMux
    port map (
            O => \N__10199\,
            I => \N__10194\
        );

    \I__2352\ : CEMux
    port map (
            O => \N__10198\,
            I => \N__10191\
        );

    \I__2351\ : CEMux
    port map (
            O => \N__10197\,
            I => \N__10187\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__10194\,
            I => \N__10182\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__10191\,
            I => \N__10182\
        );

    \I__2348\ : CEMux
    port map (
            O => \N__10190\,
            I => \N__10179\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__10187\,
            I => \N__10174\
        );

    \I__2346\ : Span4Mux_v
    port map (
            O => \N__10182\,
            I => \N__10171\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__10179\,
            I => \N__10168\
        );

    \I__2344\ : CEMux
    port map (
            O => \N__10178\,
            I => \N__10165\
        );

    \I__2343\ : CEMux
    port map (
            O => \N__10177\,
            I => \N__10162\
        );

    \I__2342\ : Span4Mux_h
    port map (
            O => \N__10174\,
            I => \N__10159\
        );

    \I__2341\ : Span4Mux_v
    port map (
            O => \N__10171\,
            I => \N__10152\
        );

    \I__2340\ : Span4Mux_h
    port map (
            O => \N__10168\,
            I => \N__10152\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__10165\,
            I => \N__10152\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__10162\,
            I => \N__10149\
        );

    \I__2337\ : Span4Mux_v
    port map (
            O => \N__10159\,
            I => \N__10146\
        );

    \I__2336\ : Span4Mux_h
    port map (
            O => \N__10152\,
            I => \N__10143\
        );

    \I__2335\ : Span4Mux_h
    port map (
            O => \N__10149\,
            I => \N__10140\
        );

    \I__2334\ : Odrv4
    port map (
            O => \N__10146\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2333\ : Odrv4
    port map (
            O => \N__10143\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2332\ : Odrv4
    port map (
            O => \N__10140\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2331\ : InMux
    port map (
            O => \N__10133\,
            I => \N__10127\
        );

    \I__2330\ : InMux
    port map (
            O => \N__10132\,
            I => \N__10124\
        );

    \I__2329\ : InMux
    port map (
            O => \N__10131\,
            I => \N__10121\
        );

    \I__2328\ : InMux
    port map (
            O => \N__10130\,
            I => \N__10118\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__10127\,
            I => \N__10111\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__10124\,
            I => \N__10111\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__10121\,
            I => \N__10111\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__10118\,
            I => \N__10108\
        );

    \I__2323\ : Span4Mux_v
    port map (
            O => \N__10111\,
            I => \N__10105\
        );

    \I__2322\ : Span4Mux_v
    port map (
            O => \N__10108\,
            I => \N__10102\
        );

    \I__2321\ : Sp12to4
    port map (
            O => \N__10105\,
            I => \N__10099\
        );

    \I__2320\ : Sp12to4
    port map (
            O => \N__10102\,
            I => \N__10096\
        );

    \I__2319\ : Span12Mux_h
    port map (
            O => \N__10099\,
            I => \N__10093\
        );

    \I__2318\ : Odrv12
    port map (
            O => \N__10096\,
            I => \DRA_c_5\
        );

    \I__2317\ : Odrv12
    port map (
            O => \N__10093\,
            I => \DRA_c_5\
        );

    \I__2316\ : InMux
    port map (
            O => \N__10088\,
            I => \N__10085\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__10085\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2314\ : InMux
    port map (
            O => \N__10082\,
            I => \N__10074\
        );

    \I__2313\ : InMux
    port map (
            O => \N__10081\,
            I => \N__10074\
        );

    \I__2312\ : InMux
    port map (
            O => \N__10080\,
            I => \N__10071\
        );

    \I__2311\ : InMux
    port map (
            O => \N__10079\,
            I => \N__10068\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__10074\,
            I => \N__10065\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__10071\,
            I => \N__10060\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__10068\,
            I => \N__10060\
        );

    \I__2307\ : Span4Mux_v
    port map (
            O => \N__10065\,
            I => \N__10057\
        );

    \I__2306\ : Span12Mux_v
    port map (
            O => \N__10060\,
            I => \N__10052\
        );

    \I__2305\ : Sp12to4
    port map (
            O => \N__10057\,
            I => \N__10052\
        );

    \I__2304\ : Span12Mux_h
    port map (
            O => \N__10052\,
            I => \N__10049\
        );

    \I__2303\ : Odrv12
    port map (
            O => \N__10049\,
            I => \DRA_c_4\
        );

    \I__2302\ : InMux
    port map (
            O => \N__10046\,
            I => \N__10038\
        );

    \I__2301\ : InMux
    port map (
            O => \N__10045\,
            I => \N__10038\
        );

    \I__2300\ : InMux
    port map (
            O => \N__10044\,
            I => \N__10035\
        );

    \I__2299\ : InMux
    port map (
            O => \N__10043\,
            I => \N__10032\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__10038\,
            I => \N__10027\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__10035\,
            I => \N__10027\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__10032\,
            I => \N__10024\
        );

    \I__2295\ : Span4Mux_v
    port map (
            O => \N__10027\,
            I => \N__10021\
        );

    \I__2294\ : Span4Mux_v
    port map (
            O => \N__10024\,
            I => \N__10018\
        );

    \I__2293\ : Sp12to4
    port map (
            O => \N__10021\,
            I => \N__10015\
        );

    \I__2292\ : Sp12to4
    port map (
            O => \N__10018\,
            I => \N__10012\
        );

    \I__2291\ : Span12Mux_h
    port map (
            O => \N__10015\,
            I => \N__10009\
        );

    \I__2290\ : Odrv12
    port map (
            O => \N__10012\,
            I => \DRA_c_3\
        );

    \I__2289\ : Odrv12
    port map (
            O => \N__10009\,
            I => \DRA_c_3\
        );

    \I__2288\ : CascadeMux
    port map (
            O => \N__10004\,
            I => \N__10001\
        );

    \I__2287\ : InMux
    port map (
            O => \N__10001\,
            I => \N__9998\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__9998\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2285\ : InMux
    port map (
            O => \N__9995\,
            I => \N__9992\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__9992\,
            I => \N__9989\
        );

    \I__2283\ : Span4Mux_h
    port map (
            O => \N__9989\,
            I => \N__9986\
        );

    \I__2282\ : Odrv4
    port map (
            O => \N__9986\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__2281\ : InMux
    port map (
            O => \N__9983\,
            I => \N__9980\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__9980\,
            I => \N__9977\
        );

    \I__2279\ : Span4Mux_v
    port map (
            O => \N__9977\,
            I => \N__9974\
        );

    \I__2278\ : Span4Mux_h
    port map (
            O => \N__9974\,
            I => \N__9971\
        );

    \I__2277\ : Odrv4
    port map (
            O => \N__9971\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2276\ : CascadeMux
    port map (
            O => \N__9968\,
            I => \N__9965\
        );

    \I__2275\ : InMux
    port map (
            O => \N__9965\,
            I => \N__9962\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__9962\,
            I => \N__9959\
        );

    \I__2273\ : Odrv12
    port map (
            O => \N__9959\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__2272\ : InMux
    port map (
            O => \N__9956\,
            I => \N__9953\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__9953\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__2270\ : IoInMux
    port map (
            O => \N__9950\,
            I => \N__9947\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__9947\,
            I => \N__9944\
        );

    \I__2268\ : IoSpan4Mux
    port map (
            O => \N__9944\,
            I => \N__9941\
        );

    \I__2267\ : Sp12to4
    port map (
            O => \N__9941\,
            I => \N__9938\
        );

    \I__2266\ : Span12Mux_s9_v
    port map (
            O => \N__9938\,
            I => \N__9935\
        );

    \I__2265\ : Odrv12
    port map (
            O => \N__9935\,
            I => \CMA_c_2\
        );

    \I__2264\ : InMux
    port map (
            O => \N__9932\,
            I => \N__9929\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__9929\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__2262\ : IoInMux
    port map (
            O => \N__9926\,
            I => \N__9923\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__9923\,
            I => \N__9920\
        );

    \I__2260\ : Span4Mux_s1_h
    port map (
            O => \N__9920\,
            I => \N__9917\
        );

    \I__2259\ : Sp12to4
    port map (
            O => \N__9917\,
            I => \N__9914\
        );

    \I__2258\ : Span12Mux_v
    port map (
            O => \N__9914\,
            I => \N__9911\
        );

    \I__2257\ : Span12Mux_h
    port map (
            O => \N__9911\,
            I => \N__9908\
        );

    \I__2256\ : Odrv12
    port map (
            O => \N__9908\,
            I => \CMA_c_3\
        );

    \I__2255\ : CascadeMux
    port map (
            O => \N__9905\,
            I => \N__9902\
        );

    \I__2254\ : InMux
    port map (
            O => \N__9902\,
            I => \N__9899\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__9899\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__2252\ : InMux
    port map (
            O => \N__9896\,
            I => \N__9893\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__9893\,
            I => \N__9890\
        );

    \I__2250\ : Span4Mux_h
    port map (
            O => \N__9890\,
            I => \N__9887\
        );

    \I__2249\ : Odrv4
    port map (
            O => \N__9887\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__2248\ : InMux
    port map (
            O => \N__9884\,
            I => \N__9881\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__9881\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__2246\ : InMux
    port map (
            O => \N__9878\,
            I => \N__9875\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__9875\,
            I => \N__9872\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__9872\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__2243\ : InMux
    port map (
            O => \N__9869\,
            I => \N__9865\
        );

    \I__2242\ : InMux
    port map (
            O => \N__9868\,
            I => \N__9860\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__9865\,
            I => \N__9857\
        );

    \I__2240\ : InMux
    port map (
            O => \N__9864\,
            I => \N__9853\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__9863\,
            I => \N__9850\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__9860\,
            I => \N__9847\
        );

    \I__2237\ : Sp12to4
    port map (
            O => \N__9857\,
            I => \N__9844\
        );

    \I__2236\ : InMux
    port map (
            O => \N__9856\,
            I => \N__9840\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__9853\,
            I => \N__9836\
        );

    \I__2234\ : InMux
    port map (
            O => \N__9850\,
            I => \N__9833\
        );

    \I__2233\ : Span12Mux_h
    port map (
            O => \N__9847\,
            I => \N__9830\
        );

    \I__2232\ : Span12Mux_v
    port map (
            O => \N__9844\,
            I => \N__9827\
        );

    \I__2231\ : InMux
    port map (
            O => \N__9843\,
            I => \N__9824\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__9840\,
            I => \N__9821\
        );

    \I__2229\ : InMux
    port map (
            O => \N__9839\,
            I => \N__9818\
        );

    \I__2228\ : Span4Mux_h
    port map (
            O => \N__9836\,
            I => \N__9815\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__9833\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2226\ : Odrv12
    port map (
            O => \N__9830\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2225\ : Odrv12
    port map (
            O => \N__9827\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__9824\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__9821\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__9818\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2221\ : Odrv4
    port map (
            O => \N__9815\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2220\ : IoInMux
    port map (
            O => \N__9800\,
            I => \N__9797\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__9797\,
            I => \N__9794\
        );

    \I__2218\ : Span4Mux_s3_h
    port map (
            O => \N__9794\,
            I => \N__9791\
        );

    \I__2217\ : Span4Mux_v
    port map (
            O => \N__9791\,
            I => \N__9788\
        );

    \I__2216\ : Span4Mux_h
    port map (
            O => \N__9788\,
            I => \N__9785\
        );

    \I__2215\ : Span4Mux_h
    port map (
            O => \N__9785\,
            I => \N__9782\
        );

    \I__2214\ : Odrv4
    port map (
            O => \N__9782\,
            I => \WEn_c\
        );

    \I__2213\ : InMux
    port map (
            O => \N__9779\,
            I => \N__9776\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__9776\,
            I => \N__9772\
        );

    \I__2211\ : InMux
    port map (
            O => \N__9775\,
            I => \N__9769\
        );

    \I__2210\ : Span4Mux_v
    port map (
            O => \N__9772\,
            I => \N__9762\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__9769\,
            I => \N__9762\
        );

    \I__2208\ : InMux
    port map (
            O => \N__9768\,
            I => \N__9759\
        );

    \I__2207\ : InMux
    port map (
            O => \N__9767\,
            I => \N__9753\
        );

    \I__2206\ : Span4Mux_h
    port map (
            O => \N__9762\,
            I => \N__9750\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__9759\,
            I => \N__9747\
        );

    \I__2204\ : InMux
    port map (
            O => \N__9758\,
            I => \N__9744\
        );

    \I__2203\ : InMux
    port map (
            O => \N__9757\,
            I => \N__9741\
        );

    \I__2202\ : InMux
    port map (
            O => \N__9756\,
            I => \N__9738\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__9753\,
            I => \N__9735\
        );

    \I__2200\ : Span4Mux_v
    port map (
            O => \N__9750\,
            I => \N__9730\
        );

    \I__2199\ : Span4Mux_h
    port map (
            O => \N__9747\,
            I => \N__9730\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__9744\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__9741\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__9738\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2195\ : Odrv4
    port map (
            O => \N__9735\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2194\ : Odrv4
    port map (
            O => \N__9730\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2193\ : IoInMux
    port map (
            O => \N__9719\,
            I => \N__9716\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__9716\,
            I => \N__9713\
        );

    \I__2191\ : Span12Mux_s9_v
    port map (
            O => \N__9713\,
            I => \N__9710\
        );

    \I__2190\ : Odrv12
    port map (
            O => \N__9710\,
            I => \RASn_c\
        );

    \I__2189\ : InMux
    port map (
            O => \N__9707\,
            I => \N__9700\
        );

    \I__2188\ : InMux
    port map (
            O => \N__9706\,
            I => \N__9695\
        );

    \I__2187\ : CascadeMux
    port map (
            O => \N__9705\,
            I => \N__9692\
        );

    \I__2186\ : CascadeMux
    port map (
            O => \N__9704\,
            I => \N__9687\
        );

    \I__2185\ : CascadeMux
    port map (
            O => \N__9703\,
            I => \N__9683\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__9700\,
            I => \N__9680\
        );

    \I__2183\ : InMux
    port map (
            O => \N__9699\,
            I => \N__9677\
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__9698\,
            I => \N__9674\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__9695\,
            I => \N__9671\
        );

    \I__2180\ : InMux
    port map (
            O => \N__9692\,
            I => \N__9664\
        );

    \I__2179\ : InMux
    port map (
            O => \N__9691\,
            I => \N__9664\
        );

    \I__2178\ : CascadeMux
    port map (
            O => \N__9690\,
            I => \N__9661\
        );

    \I__2177\ : InMux
    port map (
            O => \N__9687\,
            I => \N__9652\
        );

    \I__2176\ : InMux
    port map (
            O => \N__9686\,
            I => \N__9652\
        );

    \I__2175\ : InMux
    port map (
            O => \N__9683\,
            I => \N__9652\
        );

    \I__2174\ : Span4Mux_v
    port map (
            O => \N__9680\,
            I => \N__9647\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__9677\,
            I => \N__9647\
        );

    \I__2172\ : InMux
    port map (
            O => \N__9674\,
            I => \N__9644\
        );

    \I__2171\ : Span4Mux_v
    port map (
            O => \N__9671\,
            I => \N__9638\
        );

    \I__2170\ : InMux
    port map (
            O => \N__9670\,
            I => \N__9633\
        );

    \I__2169\ : InMux
    port map (
            O => \N__9669\,
            I => \N__9633\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__9664\,
            I => \N__9630\
        );

    \I__2167\ : InMux
    port map (
            O => \N__9661\,
            I => \N__9617\
        );

    \I__2166\ : InMux
    port map (
            O => \N__9660\,
            I => \N__9617\
        );

    \I__2165\ : InMux
    port map (
            O => \N__9659\,
            I => \N__9617\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__9652\,
            I => \N__9612\
        );

    \I__2163\ : Span4Mux_v
    port map (
            O => \N__9647\,
            I => \N__9612\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__9644\,
            I => \N__9609\
        );

    \I__2161\ : InMux
    port map (
            O => \N__9643\,
            I => \N__9602\
        );

    \I__2160\ : InMux
    port map (
            O => \N__9642\,
            I => \N__9602\
        );

    \I__2159\ : InMux
    port map (
            O => \N__9641\,
            I => \N__9602\
        );

    \I__2158\ : Span4Mux_v
    port map (
            O => \N__9638\,
            I => \N__9597\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__9633\,
            I => \N__9597\
        );

    \I__2156\ : Span4Mux_h
    port map (
            O => \N__9630\,
            I => \N__9594\
        );

    \I__2155\ : InMux
    port map (
            O => \N__9629\,
            I => \N__9589\
        );

    \I__2154\ : InMux
    port map (
            O => \N__9628\,
            I => \N__9589\
        );

    \I__2153\ : InMux
    port map (
            O => \N__9627\,
            I => \N__9582\
        );

    \I__2152\ : InMux
    port map (
            O => \N__9626\,
            I => \N__9582\
        );

    \I__2151\ : InMux
    port map (
            O => \N__9625\,
            I => \N__9582\
        );

    \I__2150\ : InMux
    port map (
            O => \N__9624\,
            I => \N__9579\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__9617\,
            I => \N__9576\
        );

    \I__2148\ : Span4Mux_h
    port map (
            O => \N__9612\,
            I => \N__9571\
        );

    \I__2147\ : Span4Mux_h
    port map (
            O => \N__9609\,
            I => \N__9571\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__9602\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2145\ : Odrv4
    port map (
            O => \N__9597\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2144\ : Odrv4
    port map (
            O => \N__9594\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__9589\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__9582\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__9579\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2140\ : Odrv12
    port map (
            O => \N__9576\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2139\ : Odrv4
    port map (
            O => \N__9571\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2138\ : IoInMux
    port map (
            O => \N__9554\,
            I => \N__9551\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__9551\,
            I => \N__9548\
        );

    \I__2136\ : Span12Mux_s10_v
    port map (
            O => \N__9548\,
            I => \N__9545\
        );

    \I__2135\ : Odrv12
    port map (
            O => \N__9545\,
            I => \CASn_c\
        );

    \I__2134\ : CascadeMux
    port map (
            O => \N__9542\,
            I => \N__9538\
        );

    \I__2133\ : InMux
    port map (
            O => \N__9541\,
            I => \N__9535\
        );

    \I__2132\ : InMux
    port map (
            O => \N__9538\,
            I => \N__9532\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__9535\,
            I => \N__9529\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__9532\,
            I => \N__9526\
        );

    \I__2129\ : Span4Mux_v
    port map (
            O => \N__9529\,
            I => \N__9523\
        );

    \I__2128\ : Odrv12
    port map (
            O => \N__9526\,
            I => \DBRn_c_i\
        );

    \I__2127\ : Odrv4
    port map (
            O => \N__9523\,
            I => \DBRn_c_i\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9518\,
            I => \N__9515\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__9515\,
            I => \N__9511\
        );

    \I__2124\ : InMux
    port map (
            O => \N__9514\,
            I => \N__9508\
        );

    \I__2123\ : Span4Mux_h
    port map (
            O => \N__9511\,
            I => \N__9505\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__9508\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__2121\ : Odrv4
    port map (
            O => \N__9505\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__2120\ : InMux
    port map (
            O => \N__9500\,
            I => \N__9496\
        );

    \I__2119\ : CascadeMux
    port map (
            O => \N__9499\,
            I => \N__9493\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__9496\,
            I => \N__9490\
        );

    \I__2117\ : InMux
    port map (
            O => \N__9493\,
            I => \N__9487\
        );

    \I__2116\ : Span4Mux_v
    port map (
            O => \N__9490\,
            I => \N__9480\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__9487\,
            I => \N__9480\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__9486\,
            I => \N__9477\
        );

    \I__2113\ : InMux
    port map (
            O => \N__9485\,
            I => \N__9474\
        );

    \I__2112\ : Span4Mux_h
    port map (
            O => \N__9480\,
            I => \N__9471\
        );

    \I__2111\ : InMux
    port map (
            O => \N__9477\,
            I => \N__9468\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__9474\,
            I => \N__9465\
        );

    \I__2109\ : Span4Mux_v
    port map (
            O => \N__9471\,
            I => \N__9458\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__9468\,
            I => \N__9458\
        );

    \I__2107\ : Span4Mux_h
    port map (
            O => \N__9465\,
            I => \N__9458\
        );

    \I__2106\ : Odrv4
    port map (
            O => \N__9458\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2105\ : IoInMux
    port map (
            O => \N__9455\,
            I => \N__9452\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__9452\,
            I => \N__9449\
        );

    \I__2103\ : Span4Mux_s3_v
    port map (
            O => \N__9449\,
            I => \N__9446\
        );

    \I__2102\ : Span4Mux_v
    port map (
            O => \N__9446\,
            I => \N__9443\
        );

    \I__2101\ : Span4Mux_h
    port map (
            O => \N__9443\,
            I => \N__9440\
        );

    \I__2100\ : Odrv4
    port map (
            O => \N__9440\,
            I => \CRCSn_c\
        );

    \I__2099\ : InMux
    port map (
            O => \N__9437\,
            I => \N__9433\
        );

    \I__2098\ : InMux
    port map (
            O => \N__9436\,
            I => \N__9430\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__9433\,
            I => \N__9424\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__9430\,
            I => \N__9424\
        );

    \I__2095\ : CascadeMux
    port map (
            O => \N__9429\,
            I => \N__9421\
        );

    \I__2094\ : Span4Mux_h
    port map (
            O => \N__9424\,
            I => \N__9417\
        );

    \I__2093\ : InMux
    port map (
            O => \N__9421\,
            I => \N__9412\
        );

    \I__2092\ : InMux
    port map (
            O => \N__9420\,
            I => \N__9412\
        );

    \I__2091\ : Span4Mux_v
    port map (
            O => \N__9417\,
            I => \N__9409\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__9412\,
            I => \N__9406\
        );

    \I__2089\ : Odrv4
    port map (
            O => \N__9409\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__2088\ : Odrv12
    port map (
            O => \N__9406\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__2087\ : InMux
    port map (
            O => \N__9401\,
            I => \N__9398\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__9398\,
            I => \N__9395\
        );

    \I__2085\ : Sp12to4
    port map (
            O => \N__9395\,
            I => \N__9392\
        );

    \I__2084\ : Span12Mux_v
    port map (
            O => \N__9392\,
            I => \N__9389\
        );

    \I__2083\ : Span12Mux_h
    port map (
            O => \N__9389\,
            I => \N__9386\
        );

    \I__2082\ : Odrv12
    port map (
            O => \N__9386\,
            I => \A_c_19\
        );

    \I__2081\ : IoInMux
    port map (
            O => \N__9383\,
            I => \N__9380\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__9380\,
            I => \N__9377\
        );

    \I__2079\ : IoSpan4Mux
    port map (
            O => \N__9377\,
            I => \N__9374\
        );

    \I__2078\ : Span4Mux_s2_h
    port map (
            O => \N__9374\,
            I => \N__9371\
        );

    \I__2077\ : Span4Mux_v
    port map (
            O => \N__9371\,
            I => \N__9368\
        );

    \I__2076\ : Sp12to4
    port map (
            O => \N__9368\,
            I => \N__9365\
        );

    \I__2075\ : Odrv12
    port map (
            O => \N__9365\,
            I => \CMA_c_9\
        );

    \I__2074\ : InMux
    port map (
            O => \N__9362\,
            I => \N__9359\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__9359\,
            I => \N__9356\
        );

    \I__2072\ : Odrv4
    port map (
            O => \N__9356\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\
        );

    \I__2071\ : InMux
    port map (
            O => \N__9353\,
            I => \N__9350\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__9350\,
            I => \N__9347\
        );

    \I__2069\ : Odrv4
    port map (
            O => \N__9347\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\
        );

    \I__2068\ : CascadeMux
    port map (
            O => \N__9344\,
            I => \N__9334\
        );

    \I__2067\ : CascadeMux
    port map (
            O => \N__9343\,
            I => \N__9328\
        );

    \I__2066\ : CascadeMux
    port map (
            O => \N__9342\,
            I => \N__9325\
        );

    \I__2065\ : CascadeMux
    port map (
            O => \N__9341\,
            I => \N__9321\
        );

    \I__2064\ : CascadeMux
    port map (
            O => \N__9340\,
            I => \N__9318\
        );

    \I__2063\ : CascadeMux
    port map (
            O => \N__9339\,
            I => \N__9315\
        );

    \I__2062\ : CascadeMux
    port map (
            O => \N__9338\,
            I => \N__9310\
        );

    \I__2061\ : InMux
    port map (
            O => \N__9337\,
            I => \N__9300\
        );

    \I__2060\ : InMux
    port map (
            O => \N__9334\,
            I => \N__9296\
        );

    \I__2059\ : InMux
    port map (
            O => \N__9333\,
            I => \N__9293\
        );

    \I__2058\ : InMux
    port map (
            O => \N__9332\,
            I => \N__9288\
        );

    \I__2057\ : InMux
    port map (
            O => \N__9331\,
            I => \N__9288\
        );

    \I__2056\ : InMux
    port map (
            O => \N__9328\,
            I => \N__9285\
        );

    \I__2055\ : InMux
    port map (
            O => \N__9325\,
            I => \N__9274\
        );

    \I__2054\ : InMux
    port map (
            O => \N__9324\,
            I => \N__9274\
        );

    \I__2053\ : InMux
    port map (
            O => \N__9321\,
            I => \N__9274\
        );

    \I__2052\ : InMux
    port map (
            O => \N__9318\,
            I => \N__9274\
        );

    \I__2051\ : InMux
    port map (
            O => \N__9315\,
            I => \N__9274\
        );

    \I__2050\ : InMux
    port map (
            O => \N__9314\,
            I => \N__9271\
        );

    \I__2049\ : InMux
    port map (
            O => \N__9313\,
            I => \N__9268\
        );

    \I__2048\ : InMux
    port map (
            O => \N__9310\,
            I => \N__9265\
        );

    \I__2047\ : InMux
    port map (
            O => \N__9309\,
            I => \N__9258\
        );

    \I__2046\ : InMux
    port map (
            O => \N__9308\,
            I => \N__9258\
        );

    \I__2045\ : InMux
    port map (
            O => \N__9307\,
            I => \N__9258\
        );

    \I__2044\ : InMux
    port map (
            O => \N__9306\,
            I => \N__9251\
        );

    \I__2043\ : InMux
    port map (
            O => \N__9305\,
            I => \N__9251\
        );

    \I__2042\ : InMux
    port map (
            O => \N__9304\,
            I => \N__9251\
        );

    \I__2041\ : InMux
    port map (
            O => \N__9303\,
            I => \N__9246\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__9300\,
            I => \N__9243\
        );

    \I__2039\ : InMux
    port map (
            O => \N__9299\,
            I => \N__9240\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__9296\,
            I => \N__9237\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__9293\,
            I => \N__9234\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__9288\,
            I => \N__9225\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__9285\,
            I => \N__9225\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__9274\,
            I => \N__9225\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__9271\,
            I => \N__9225\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__9268\,
            I => \N__9222\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__9265\,
            I => \N__9219\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__9258\,
            I => \N__9214\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__9251\,
            I => \N__9214\
        );

    \I__2028\ : InMux
    port map (
            O => \N__9250\,
            I => \N__9211\
        );

    \I__2027\ : InMux
    port map (
            O => \N__9249\,
            I => \N__9208\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__9246\,
            I => \N__9205\
        );

    \I__2025\ : Span4Mux_v
    port map (
            O => \N__9243\,
            I => \N__9194\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__9240\,
            I => \N__9194\
        );

    \I__2023\ : Span4Mux_v
    port map (
            O => \N__9237\,
            I => \N__9194\
        );

    \I__2022\ : Span4Mux_h
    port map (
            O => \N__9234\,
            I => \N__9194\
        );

    \I__2021\ : Span4Mux_v
    port map (
            O => \N__9225\,
            I => \N__9194\
        );

    \I__2020\ : Span4Mux_v
    port map (
            O => \N__9222\,
            I => \N__9187\
        );

    \I__2019\ : Span4Mux_h
    port map (
            O => \N__9219\,
            I => \N__9187\
        );

    \I__2018\ : Span4Mux_h
    port map (
            O => \N__9214\,
            I => \N__9187\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__9211\,
            I => \N__9184\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__9208\,
            I => \CPU_CYCLEm\
        );

    \I__2015\ : Odrv4
    port map (
            O => \N__9205\,
            I => \CPU_CYCLEm\
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__9194\,
            I => \CPU_CYCLEm\
        );

    \I__2013\ : Odrv4
    port map (
            O => \N__9187\,
            I => \CPU_CYCLEm\
        );

    \I__2012\ : Odrv12
    port map (
            O => \N__9184\,
            I => \CPU_CYCLEm\
        );

    \I__2011\ : InMux
    port map (
            O => \N__9173\,
            I => \N__9170\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__9170\,
            I => \N__9167\
        );

    \I__2009\ : Odrv4
    port map (
            O => \N__9167\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__2008\ : InMux
    port map (
            O => \N__9164\,
            I => \N__9161\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__9161\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__2006\ : InMux
    port map (
            O => \N__9158\,
            I => \N__9155\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__9155\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2004\ : InMux
    port map (
            O => \N__9152\,
            I => \N__9149\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__9149\,
            I => \N__9146\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__9146\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__2001\ : IoInMux
    port map (
            O => \N__9143\,
            I => \N__9140\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__9140\,
            I => \N__9137\
        );

    \I__1999\ : Span4Mux_s1_v
    port map (
            O => \N__9137\,
            I => \N__9134\
        );

    \I__1998\ : Sp12to4
    port map (
            O => \N__9134\,
            I => \N__9131\
        );

    \I__1997\ : Span12Mux_h
    port map (
            O => \N__9131\,
            I => \N__9128\
        );

    \I__1996\ : Span12Mux_v
    port map (
            O => \N__9128\,
            I => \N__9125\
        );

    \I__1995\ : Odrv12
    port map (
            O => \N__9125\,
            I => \CMA_c_0\
        );

    \I__1994\ : InMux
    port map (
            O => \N__9122\,
            I => \N__9119\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__9119\,
            I => \N__9116\
        );

    \I__1992\ : Span4Mux_v
    port map (
            O => \N__9116\,
            I => \N__9113\
        );

    \I__1991\ : Span4Mux_v
    port map (
            O => \N__9113\,
            I => \N__9110\
        );

    \I__1990\ : Sp12to4
    port map (
            O => \N__9110\,
            I => \N__9107\
        );

    \I__1989\ : Span12Mux_h
    port map (
            O => \N__9107\,
            I => \N__9104\
        );

    \I__1988\ : Odrv12
    port map (
            O => \N__9104\,
            I => \A_c_17\
        );

    \I__1987\ : IoInMux
    port map (
            O => \N__9101\,
            I => \N__9098\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__9098\,
            I => \N__9095\
        );

    \I__1985\ : IoSpan4Mux
    port map (
            O => \N__9095\,
            I => \N__9092\
        );

    \I__1984\ : IoSpan4Mux
    port map (
            O => \N__9092\,
            I => \N__9089\
        );

    \I__1983\ : Sp12to4
    port map (
            O => \N__9089\,
            I => \N__9086\
        );

    \I__1982\ : Span12Mux_s9_h
    port map (
            O => \N__9086\,
            I => \N__9083\
        );

    \I__1981\ : Odrv12
    port map (
            O => \N__9083\,
            I => \CMA_c_8\
        );

    \I__1980\ : InMux
    port map (
            O => \N__9080\,
            I => \N__9077\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__9077\,
            I => \N__9074\
        );

    \I__1978\ : Odrv4
    port map (
            O => \N__9074\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__1977\ : CascadeMux
    port map (
            O => \N__9071\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5_cascade_\
        );

    \I__1976\ : InMux
    port map (
            O => \N__9068\,
            I => \N__9065\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__9065\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\
        );

    \I__1974\ : IoInMux
    port map (
            O => \N__9062\,
            I => \N__9059\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__9059\,
            I => \N__9056\
        );

    \I__1972\ : Span12Mux_s2_h
    port map (
            O => \N__9056\,
            I => \N__9053\
        );

    \I__1971\ : Span12Mux_h
    port map (
            O => \N__9053\,
            I => \N__9050\
        );

    \I__1970\ : Span12Mux_v
    port map (
            O => \N__9050\,
            I => \N__9047\
        );

    \I__1969\ : Odrv12
    port map (
            O => \N__9047\,
            I => \CMA_c_5\
        );

    \I__1968\ : InMux
    port map (
            O => \N__9044\,
            I => \N__9038\
        );

    \I__1967\ : InMux
    port map (
            O => \N__9043\,
            I => \N__9038\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__9038\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__1965\ : InMux
    port map (
            O => \N__9035\,
            I => \N__9032\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__9032\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\
        );

    \I__1963\ : InMux
    port map (
            O => \N__9029\,
            I => \N__9026\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__9026\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\
        );

    \I__1961\ : InMux
    port map (
            O => \N__9023\,
            I => \N__9020\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__9020\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\
        );

    \I__1959\ : CascadeMux
    port map (
            O => \N__9017\,
            I => \U712_CHIP_RAM.N_11_cascade_\
        );

    \I__1958\ : InMux
    port map (
            O => \N__9014\,
            I => \N__9011\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__9011\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\
        );

    \I__1956\ : InMux
    port map (
            O => \N__9008\,
            I => \N__9005\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__9005\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5\
        );

    \I__1954\ : IoInMux
    port map (
            O => \N__9002\,
            I => \N__8999\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__8999\,
            I => \N__8996\
        );

    \I__1952\ : IoSpan4Mux
    port map (
            O => \N__8996\,
            I => \N__8993\
        );

    \I__1951\ : Span4Mux_s2_v
    port map (
            O => \N__8993\,
            I => \N__8988\
        );

    \I__1950\ : InMux
    port map (
            O => \N__8992\,
            I => \N__8983\
        );

    \I__1949\ : InMux
    port map (
            O => \N__8991\,
            I => \N__8983\
        );

    \I__1948\ : Sp12to4
    port map (
            O => \N__8988\,
            I => \N__8980\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__8983\,
            I => \N__8977\
        );

    \I__1946\ : Span12Mux_s8_v
    port map (
            O => \N__8980\,
            I => \N__8972\
        );

    \I__1945\ : Sp12to4
    port map (
            O => \N__8977\,
            I => \N__8972\
        );

    \I__1944\ : Span12Mux_v
    port map (
            O => \N__8972\,
            I => \N__8969\
        );

    \I__1943\ : Span12Mux_h
    port map (
            O => \N__8969\,
            I => \N__8966\
        );

    \I__1942\ : Odrv12
    port map (
            O => \N__8966\,
            I => \A_c_10\
        );

    \I__1941\ : InMux
    port map (
            O => \N__8963\,
            I => \N__8960\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__8960\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__1939\ : InMux
    port map (
            O => \N__8957\,
            I => \N__8954\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__8954\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__1937\ : InMux
    port map (
            O => \N__8951\,
            I => \N__8948\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__8948\,
            I => \N__8945\
        );

    \I__1935\ : Span4Mux_v
    port map (
            O => \N__8945\,
            I => \N__8942\
        );

    \I__1934\ : Sp12to4
    port map (
            O => \N__8942\,
            I => \N__8939\
        );

    \I__1933\ : Span12Mux_h
    port map (
            O => \N__8939\,
            I => \N__8936\
        );

    \I__1932\ : Odrv12
    port map (
            O => \N__8936\,
            I => \A_c_5\
        );

    \I__1931\ : InMux
    port map (
            O => \N__8933\,
            I => \N__8930\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__8930\,
            I => \N__8927\
        );

    \I__1929\ : Sp12to4
    port map (
            O => \N__8927\,
            I => \N__8924\
        );

    \I__1928\ : Span12Mux_v
    port map (
            O => \N__8924\,
            I => \N__8921\
        );

    \I__1927\ : Span12Mux_h
    port map (
            O => \N__8921\,
            I => \N__8918\
        );

    \I__1926\ : Odrv12
    port map (
            O => \N__8918\,
            I => \A_c_12\
        );

    \I__1925\ : InMux
    port map (
            O => \N__8915\,
            I => \N__8912\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__8912\,
            I => \N__8909\
        );

    \I__1923\ : Span4Mux_v
    port map (
            O => \N__8909\,
            I => \N__8906\
        );

    \I__1922\ : Sp12to4
    port map (
            O => \N__8906\,
            I => \N__8903\
        );

    \I__1921\ : Span12Mux_h
    port map (
            O => \N__8903\,
            I => \N__8900\
        );

    \I__1920\ : Odrv12
    port map (
            O => \N__8900\,
            I => \A_c_4\
        );

    \I__1919\ : IoInMux
    port map (
            O => \N__8897\,
            I => \N__8894\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__8894\,
            I => \N__8891\
        );

    \I__1917\ : IoSpan4Mux
    port map (
            O => \N__8891\,
            I => \N__8887\
        );

    \I__1916\ : InMux
    port map (
            O => \N__8890\,
            I => \N__8884\
        );

    \I__1915\ : Span4Mux_s2_v
    port map (
            O => \N__8887\,
            I => \N__8881\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__8884\,
            I => \N__8878\
        );

    \I__1913\ : Sp12to4
    port map (
            O => \N__8881\,
            I => \N__8875\
        );

    \I__1912\ : Span4Mux_v
    port map (
            O => \N__8878\,
            I => \N__8872\
        );

    \I__1911\ : Span12Mux_s8_v
    port map (
            O => \N__8875\,
            I => \N__8869\
        );

    \I__1910\ : Span4Mux_v
    port map (
            O => \N__8872\,
            I => \N__8866\
        );

    \I__1909\ : Span12Mux_h
    port map (
            O => \N__8869\,
            I => \N__8863\
        );

    \I__1908\ : Sp12to4
    port map (
            O => \N__8866\,
            I => \N__8860\
        );

    \I__1907\ : Span12Mux_v
    port map (
            O => \N__8863\,
            I => \N__8857\
        );

    \I__1906\ : Span12Mux_h
    port map (
            O => \N__8860\,
            I => \N__8854\
        );

    \I__1905\ : Odrv12
    port map (
            O => \N__8857\,
            I => \A_c_11\
        );

    \I__1904\ : Odrv12
    port map (
            O => \N__8854\,
            I => \A_c_11\
        );

    \I__1903\ : IoInMux
    port map (
            O => \N__8849\,
            I => \N__8846\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__8846\,
            I => \N__8843\
        );

    \I__1901\ : Span12Mux_s11_v
    port map (
            O => \N__8843\,
            I => \N__8840\
        );

    \I__1900\ : Odrv12
    port map (
            O => \N__8840\,
            I => \CMA_c_10\
        );

    \I__1899\ : IoInMux
    port map (
            O => \N__8837\,
            I => \N__8834\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__8834\,
            I => \N__8831\
        );

    \I__1897\ : Span4Mux_s3_v
    port map (
            O => \N__8831\,
            I => \N__8827\
        );

    \I__1896\ : InMux
    port map (
            O => \N__8830\,
            I => \N__8824\
        );

    \I__1895\ : Span4Mux_v
    port map (
            O => \N__8827\,
            I => \N__8821\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__8824\,
            I => \N__8818\
        );

    \I__1893\ : Sp12to4
    port map (
            O => \N__8821\,
            I => \N__8815\
        );

    \I__1892\ : Span4Mux_v
    port map (
            O => \N__8818\,
            I => \N__8812\
        );

    \I__1891\ : Span12Mux_h
    port map (
            O => \N__8815\,
            I => \N__8809\
        );

    \I__1890\ : Span4Mux_v
    port map (
            O => \N__8812\,
            I => \N__8806\
        );

    \I__1889\ : Odrv12
    port map (
            O => \N__8809\,
            I => \UMBEn_c\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__8806\,
            I => \UMBEn_c\
        );

    \I__1887\ : CascadeMux
    port map (
            O => \N__8801\,
            I => \U712_BYTE_ENABLE.un3_CUMBEnZ0Z_1_cascade_\
        );

    \I__1886\ : IoInMux
    port map (
            O => \N__8798\,
            I => \N__8795\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__8795\,
            I => \N__8792\
        );

    \I__1884\ : Span12Mux_s3_h
    port map (
            O => \N__8792\,
            I => \N__8789\
        );

    \I__1883\ : Span12Mux_h
    port map (
            O => \N__8789\,
            I => \N__8786\
        );

    \I__1882\ : Span12Mux_v
    port map (
            O => \N__8786\,
            I => \N__8783\
        );

    \I__1881\ : Odrv12
    port map (
            O => \N__8783\,
            I => \CUMBEn_c\
        );

    \I__1880\ : InMux
    port map (
            O => \N__8780\,
            I => \N__8776\
        );

    \I__1879\ : IoInMux
    port map (
            O => \N__8779\,
            I => \N__8773\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__8776\,
            I => \N__8770\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8773\,
            I => \N__8767\
        );

    \I__1876\ : Span4Mux_v
    port map (
            O => \N__8770\,
            I => \N__8764\
        );

    \I__1875\ : Span12Mux_s9_v
    port map (
            O => \N__8767\,
            I => \N__8761\
        );

    \I__1874\ : Span4Mux_v
    port map (
            O => \N__8764\,
            I => \N__8758\
        );

    \I__1873\ : Odrv12
    port map (
            O => \N__8761\,
            I => \UUBEn_c\
        );

    \I__1872\ : Odrv4
    port map (
            O => \N__8758\,
            I => \UUBEn_c\
        );

    \I__1871\ : CascadeMux
    port map (
            O => \N__8753\,
            I => \N__8750\
        );

    \I__1870\ : InMux
    port map (
            O => \N__8750\,
            I => \N__8747\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__8747\,
            I => \U712_BYTE_ENABLE.un3_CUMBEnZ0Z_1\
        );

    \I__1868\ : IoInMux
    port map (
            O => \N__8744\,
            I => \N__8741\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__8741\,
            I => \N__8738\
        );

    \I__1866\ : Span4Mux_s3_h
    port map (
            O => \N__8738\,
            I => \N__8735\
        );

    \I__1865\ : Sp12to4
    port map (
            O => \N__8735\,
            I => \N__8732\
        );

    \I__1864\ : Span12Mux_v
    port map (
            O => \N__8732\,
            I => \N__8729\
        );

    \I__1863\ : Span12Mux_h
    port map (
            O => \N__8729\,
            I => \N__8726\
        );

    \I__1862\ : Odrv12
    port map (
            O => \N__8726\,
            I => \CUUBEn_c\
        );

    \I__1861\ : IoInMux
    port map (
            O => \N__8723\,
            I => \N__8720\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__8720\,
            I => \N__8715\
        );

    \I__1859\ : InMux
    port map (
            O => \N__8719\,
            I => \N__8710\
        );

    \I__1858\ : InMux
    port map (
            O => \N__8718\,
            I => \N__8710\
        );

    \I__1857\ : Span12Mux_s2_v
    port map (
            O => \N__8715\,
            I => \N__8707\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__8710\,
            I => \N__8704\
        );

    \I__1855\ : Span12Mux_v
    port map (
            O => \N__8707\,
            I => \N__8700\
        );

    \I__1854\ : Span4Mux_v
    port map (
            O => \N__8704\,
            I => \N__8697\
        );

    \I__1853\ : InMux
    port map (
            O => \N__8703\,
            I => \N__8694\
        );

    \I__1852\ : Odrv12
    port map (
            O => \N__8700\,
            I => \DBENn_c\
        );

    \I__1851\ : Odrv4
    port map (
            O => \N__8697\,
            I => \DBENn_c\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__8694\,
            I => \DBENn_c\
        );

    \I__1849\ : InMux
    port map (
            O => \N__8687\,
            I => \N__8683\
        );

    \I__1848\ : InMux
    port map (
            O => \N__8686\,
            I => \N__8680\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__8683\,
            I => \N__8675\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__8680\,
            I => \N__8672\
        );

    \I__1845\ : InMux
    port map (
            O => \N__8679\,
            I => \N__8667\
        );

    \I__1844\ : InMux
    port map (
            O => \N__8678\,
            I => \N__8667\
        );

    \I__1843\ : Span4Mux_v
    port map (
            O => \N__8675\,
            I => \N__8664\
        );

    \I__1842\ : Span4Mux_h
    port map (
            O => \N__8672\,
            I => \N__8661\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__8667\,
            I => \DMA_CYCLEm\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__8664\,
            I => \DMA_CYCLEm\
        );

    \I__1839\ : Odrv4
    port map (
            O => \N__8661\,
            I => \DMA_CYCLEm\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8654\,
            I => \N__8651\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__8651\,
            I => \N__8648\
        );

    \I__1836\ : Odrv4
    port map (
            O => \N__8648\,
            I => \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_0\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8645\,
            I => \N__8642\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__8642\,
            I => \N__8639\
        );

    \I__1833\ : Span4Mux_v
    port map (
            O => \N__8639\,
            I => \N__8636\
        );

    \I__1832\ : Span4Mux_v
    port map (
            O => \N__8636\,
            I => \N__8633\
        );

    \I__1831\ : Odrv4
    port map (
            O => \N__8633\,
            I => \U712_BYTE_ENABLE.N_56\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__8630\,
            I => \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_0_cascade_\
        );

    \I__1829\ : IoInMux
    port map (
            O => \N__8627\,
            I => \N__8624\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__8624\,
            I => \N__8621\
        );

    \I__1827\ : IoSpan4Mux
    port map (
            O => \N__8621\,
            I => \N__8618\
        );

    \I__1826\ : Span4Mux_s2_v
    port map (
            O => \N__8618\,
            I => \N__8615\
        );

    \I__1825\ : Sp12to4
    port map (
            O => \N__8615\,
            I => \N__8612\
        );

    \I__1824\ : Span12Mux_v
    port map (
            O => \N__8612\,
            I => \N__8609\
        );

    \I__1823\ : Odrv12
    port map (
            O => \N__8609\,
            I => \CLLBEn_c\
        );

    \I__1822\ : IoInMux
    port map (
            O => \N__8606\,
            I => \N__8603\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__8603\,
            I => \N__8600\
        );

    \I__1820\ : IoSpan4Mux
    port map (
            O => \N__8600\,
            I => \N__8597\
        );

    \I__1819\ : Span4Mux_s2_v
    port map (
            O => \N__8597\,
            I => \N__8594\
        );

    \I__1818\ : Sp12to4
    port map (
            O => \N__8594\,
            I => \N__8591\
        );

    \I__1817\ : Span12Mux_s11_v
    port map (
            O => \N__8591\,
            I => \N__8588\
        );

    \I__1816\ : Odrv12
    port map (
            O => \N__8588\,
            I => \CMA_c_1\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8585\,
            I => \N__8582\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__8582\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8579\,
            I => \N__8576\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__8576\,
            I => \N__8573\
        );

    \I__1811\ : Span4Mux_v
    port map (
            O => \N__8573\,
            I => \N__8570\
        );

    \I__1810\ : Span4Mux_v
    port map (
            O => \N__8570\,
            I => \N__8567\
        );

    \I__1809\ : Sp12to4
    port map (
            O => \N__8567\,
            I => \N__8564\
        );

    \I__1808\ : Span12Mux_h
    port map (
            O => \N__8564\,
            I => \N__8561\
        );

    \I__1807\ : Odrv12
    port map (
            O => \N__8561\,
            I => \A_c_3\
        );

    \I__1806\ : InMux
    port map (
            O => \N__8558\,
            I => \N__8555\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__8555\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER17_1_0\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8552\,
            I => \N__8548\
        );

    \I__1803\ : InMux
    port map (
            O => \N__8551\,
            I => \N__8545\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8548\,
            I => \N__8540\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__8545\,
            I => \N__8540\
        );

    \I__1800\ : Odrv4
    port map (
            O => \N__8540\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa\
        );

    \I__1799\ : CascadeMux
    port map (
            O => \N__8537\,
            I => \U712_CHIP_RAM.N_38_cascade_\
        );

    \I__1798\ : InMux
    port map (
            O => \N__8534\,
            I => \N__8531\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__8531\,
            I => \U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8528\,
            I => \N__8525\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__8525\,
            I => \N__8522\
        );

    \I__1794\ : Span4Mux_h
    port map (
            O => \N__8522\,
            I => \N__8519\
        );

    \I__1793\ : Odrv4
    port map (
            O => \N__8519\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_i_1_1\
        );

    \I__1792\ : CascadeMux
    port map (
            O => \N__8516\,
            I => \N__8512\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8515\,
            I => \N__8509\
        );

    \I__1790\ : InMux
    port map (
            O => \N__8512\,
            I => \N__8506\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__8509\,
            I => \U712_CHIP_RAM.N_151\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__8506\,
            I => \U712_CHIP_RAM.N_151\
        );

    \I__1787\ : InMux
    port map (
            O => \N__8501\,
            I => \N__8495\
        );

    \I__1786\ : InMux
    port map (
            O => \N__8500\,
            I => \N__8495\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__8495\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER19_0\
        );

    \I__1784\ : CEMux
    port map (
            O => \N__8492\,
            I => \N__8489\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__8489\,
            I => \N__8486\
        );

    \I__1782\ : Span4Mux_v
    port map (
            O => \N__8486\,
            I => \N__8483\
        );

    \I__1781\ : Span4Mux_h
    port map (
            O => \N__8483\,
            I => \N__8480\
        );

    \I__1780\ : Odrv4
    port map (
            O => \N__8480\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_i\
        );

    \I__1779\ : InMux
    port map (
            O => \N__8477\,
            I => \N__8468\
        );

    \I__1778\ : InMux
    port map (
            O => \N__8476\,
            I => \N__8460\
        );

    \I__1777\ : InMux
    port map (
            O => \N__8475\,
            I => \N__8460\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__8474\,
            I => \N__8454\
        );

    \I__1775\ : InMux
    port map (
            O => \N__8473\,
            I => \N__8449\
        );

    \I__1774\ : InMux
    port map (
            O => \N__8472\,
            I => \N__8449\
        );

    \I__1773\ : InMux
    port map (
            O => \N__8471\,
            I => \N__8445\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__8468\,
            I => \N__8442\
        );

    \I__1771\ : InMux
    port map (
            O => \N__8467\,
            I => \N__8439\
        );

    \I__1770\ : InMux
    port map (
            O => \N__8466\,
            I => \N__8436\
        );

    \I__1769\ : InMux
    port map (
            O => \N__8465\,
            I => \N__8433\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__8460\,
            I => \N__8430\
        );

    \I__1767\ : InMux
    port map (
            O => \N__8459\,
            I => \N__8425\
        );

    \I__1766\ : InMux
    port map (
            O => \N__8458\,
            I => \N__8425\
        );

    \I__1765\ : InMux
    port map (
            O => \N__8457\,
            I => \N__8420\
        );

    \I__1764\ : InMux
    port map (
            O => \N__8454\,
            I => \N__8420\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__8449\,
            I => \N__8417\
        );

    \I__1762\ : InMux
    port map (
            O => \N__8448\,
            I => \N__8414\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__8445\,
            I => \U712_CHIP_RAM.N_331_3\
        );

    \I__1760\ : Odrv4
    port map (
            O => \N__8442\,
            I => \U712_CHIP_RAM.N_331_3\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__8439\,
            I => \U712_CHIP_RAM.N_331_3\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__8436\,
            I => \U712_CHIP_RAM.N_331_3\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__8433\,
            I => \U712_CHIP_RAM.N_331_3\
        );

    \I__1756\ : Odrv4
    port map (
            O => \N__8430\,
            I => \U712_CHIP_RAM.N_331_3\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__8425\,
            I => \U712_CHIP_RAM.N_331_3\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__8420\,
            I => \U712_CHIP_RAM.N_331_3\
        );

    \I__1753\ : Odrv4
    port map (
            O => \N__8417\,
            I => \U712_CHIP_RAM.N_331_3\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__8414\,
            I => \U712_CHIP_RAM.N_331_3\
        );

    \I__1751\ : InMux
    port map (
            O => \N__8393\,
            I => \N__8390\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__8390\,
            I => \N__8387\
        );

    \I__1749\ : Span4Mux_h
    port map (
            O => \N__8387\,
            I => \N__8384\
        );

    \I__1748\ : Odrv4
    port map (
            O => \N__8384\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_29_i_a2_i_1\
        );

    \I__1747\ : CascadeMux
    port map (
            O => \N__8381\,
            I => \U712_CHIP_RAM.N_61_cascade_\
        );

    \I__1746\ : InMux
    port map (
            O => \N__8378\,
            I => \N__8372\
        );

    \I__1745\ : InMux
    port map (
            O => \N__8377\,
            I => \N__8372\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__8372\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_1\
        );

    \I__1743\ : InMux
    port map (
            O => \N__8369\,
            I => \N__8366\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__8366\,
            I => \U712_CHIP_RAM.N_218\
        );

    \I__1741\ : InMux
    port map (
            O => \N__8363\,
            I => \N__8357\
        );

    \I__1740\ : InMux
    port map (
            O => \N__8362\,
            I => \N__8357\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__8357\,
            I => \N__8353\
        );

    \I__1738\ : InMux
    port map (
            O => \N__8356\,
            I => \N__8350\
        );

    \I__1737\ : Span4Mux_h
    port map (
            O => \N__8353\,
            I => \N__8345\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__8350\,
            I => \N__8345\
        );

    \I__1735\ : Odrv4
    port map (
            O => \N__8345\,
            I => \U712_CHIP_RAM.N_154\
        );

    \I__1734\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8339\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__8339\,
            I => \N__8334\
        );

    \I__1732\ : InMux
    port map (
            O => \N__8338\,
            I => \N__8331\
        );

    \I__1731\ : InMux
    port map (
            O => \N__8337\,
            I => \N__8323\
        );

    \I__1730\ : Span4Mux_v
    port map (
            O => \N__8334\,
            I => \N__8315\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__8331\,
            I => \N__8312\
        );

    \I__1728\ : InMux
    port map (
            O => \N__8330\,
            I => \N__8307\
        );

    \I__1727\ : InMux
    port map (
            O => \N__8329\,
            I => \N__8307\
        );

    \I__1726\ : InMux
    port map (
            O => \N__8328\,
            I => \N__8304\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__8327\,
            I => \N__8298\
        );

    \I__1724\ : InMux
    port map (
            O => \N__8326\,
            I => \N__8294\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__8323\,
            I => \N__8291\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8322\,
            I => \N__8286\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8321\,
            I => \N__8286\
        );

    \I__1720\ : InMux
    port map (
            O => \N__8320\,
            I => \N__8279\
        );

    \I__1719\ : InMux
    port map (
            O => \N__8319\,
            I => \N__8279\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8318\,
            I => \N__8279\
        );

    \I__1717\ : Span4Mux_h
    port map (
            O => \N__8315\,
            I => \N__8272\
        );

    \I__1716\ : Span4Mux_v
    port map (
            O => \N__8312\,
            I => \N__8272\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__8307\,
            I => \N__8272\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__8304\,
            I => \N__8269\
        );

    \I__1713\ : InMux
    port map (
            O => \N__8303\,
            I => \N__8266\
        );

    \I__1712\ : InMux
    port map (
            O => \N__8302\,
            I => \N__8257\
        );

    \I__1711\ : InMux
    port map (
            O => \N__8301\,
            I => \N__8257\
        );

    \I__1710\ : InMux
    port map (
            O => \N__8298\,
            I => \N__8257\
        );

    \I__1709\ : InMux
    port map (
            O => \N__8297\,
            I => \N__8257\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__8294\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1707\ : Odrv4
    port map (
            O => \N__8291\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__8286\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__8279\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1704\ : Odrv4
    port map (
            O => \N__8272\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1703\ : Odrv4
    port map (
            O => \N__8269\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__8266\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__8257\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1700\ : InMux
    port map (
            O => \N__8240\,
            I => \N__8235\
        );

    \I__1699\ : InMux
    port map (
            O => \N__8239\,
            I => \N__8231\
        );

    \I__1698\ : CascadeMux
    port map (
            O => \N__8238\,
            I => \N__8228\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__8235\,
            I => \N__8221\
        );

    \I__1696\ : CascadeMux
    port map (
            O => \N__8234\,
            I => \N__8216\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8231\,
            I => \N__8209\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8228\,
            I => \N__8204\
        );

    \I__1693\ : InMux
    port map (
            O => \N__8227\,
            I => \N__8204\
        );

    \I__1692\ : InMux
    port map (
            O => \N__8226\,
            I => \N__8201\
        );

    \I__1691\ : InMux
    port map (
            O => \N__8225\,
            I => \N__8193\
        );

    \I__1690\ : InMux
    port map (
            O => \N__8224\,
            I => \N__8190\
        );

    \I__1689\ : Span4Mux_v
    port map (
            O => \N__8221\,
            I => \N__8187\
        );

    \I__1688\ : InMux
    port map (
            O => \N__8220\,
            I => \N__8184\
        );

    \I__1687\ : InMux
    port map (
            O => \N__8219\,
            I => \N__8181\
        );

    \I__1686\ : InMux
    port map (
            O => \N__8216\,
            I => \N__8176\
        );

    \I__1685\ : InMux
    port map (
            O => \N__8215\,
            I => \N__8176\
        );

    \I__1684\ : InMux
    port map (
            O => \N__8214\,
            I => \N__8169\
        );

    \I__1683\ : InMux
    port map (
            O => \N__8213\,
            I => \N__8169\
        );

    \I__1682\ : InMux
    port map (
            O => \N__8212\,
            I => \N__8169\
        );

    \I__1681\ : Span4Mux_h
    port map (
            O => \N__8209\,
            I => \N__8162\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__8204\,
            I => \N__8162\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__8201\,
            I => \N__8162\
        );

    \I__1678\ : InMux
    port map (
            O => \N__8200\,
            I => \N__8159\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8199\,
            I => \N__8154\
        );

    \I__1676\ : InMux
    port map (
            O => \N__8198\,
            I => \N__8154\
        );

    \I__1675\ : InMux
    port map (
            O => \N__8197\,
            I => \N__8149\
        );

    \I__1674\ : InMux
    port map (
            O => \N__8196\,
            I => \N__8149\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__8193\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__8190\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1671\ : Odrv4
    port map (
            O => \N__8187\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__8184\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__8181\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__8176\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__8169\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1666\ : Odrv4
    port map (
            O => \N__8162\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__8159\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__8154\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__8149\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1662\ : CascadeMux
    port map (
            O => \N__8126\,
            I => \N__8122\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__8125\,
            I => \N__8118\
        );

    \I__1660\ : InMux
    port map (
            O => \N__8122\,
            I => \N__8114\
        );

    \I__1659\ : CascadeMux
    port map (
            O => \N__8121\,
            I => \N__8109\
        );

    \I__1658\ : InMux
    port map (
            O => \N__8118\,
            I => \N__8103\
        );

    \I__1657\ : InMux
    port map (
            O => \N__8117\,
            I => \N__8103\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__8114\,
            I => \N__8100\
        );

    \I__1655\ : InMux
    port map (
            O => \N__8113\,
            I => \N__8093\
        );

    \I__1654\ : InMux
    port map (
            O => \N__8112\,
            I => \N__8093\
        );

    \I__1653\ : InMux
    port map (
            O => \N__8109\,
            I => \N__8093\
        );

    \I__1652\ : InMux
    port map (
            O => \N__8108\,
            I => \N__8084\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__8103\,
            I => \N__8081\
        );

    \I__1650\ : Span4Mux_v
    port map (
            O => \N__8100\,
            I => \N__8076\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__8093\,
            I => \N__8076\
        );

    \I__1648\ : InMux
    port map (
            O => \N__8092\,
            I => \N__8073\
        );

    \I__1647\ : InMux
    port map (
            O => \N__8091\,
            I => \N__8070\
        );

    \I__1646\ : InMux
    port map (
            O => \N__8090\,
            I => \N__8063\
        );

    \I__1645\ : InMux
    port map (
            O => \N__8089\,
            I => \N__8063\
        );

    \I__1644\ : InMux
    port map (
            O => \N__8088\,
            I => \N__8063\
        );

    \I__1643\ : InMux
    port map (
            O => \N__8087\,
            I => \N__8060\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__8084\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1641\ : Odrv4
    port map (
            O => \N__8081\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1640\ : Odrv4
    port map (
            O => \N__8076\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__8073\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__8070\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__8063\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__8060\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1635\ : CascadeMux
    port map (
            O => \N__8045\,
            I => \N__8039\
        );

    \I__1634\ : CascadeMux
    port map (
            O => \N__8044\,
            I => \N__8036\
        );

    \I__1633\ : CascadeMux
    port map (
            O => \N__8043\,
            I => \N__8031\
        );

    \I__1632\ : InMux
    port map (
            O => \N__8042\,
            I => \N__8022\
        );

    \I__1631\ : InMux
    port map (
            O => \N__8039\,
            I => \N__8019\
        );

    \I__1630\ : InMux
    port map (
            O => \N__8036\,
            I => \N__8016\
        );

    \I__1629\ : CascadeMux
    port map (
            O => \N__8035\,
            I => \N__8012\
        );

    \I__1628\ : InMux
    port map (
            O => \N__8034\,
            I => \N__8006\
        );

    \I__1627\ : InMux
    port map (
            O => \N__8031\,
            I => \N__8001\
        );

    \I__1626\ : InMux
    port map (
            O => \N__8030\,
            I => \N__8001\
        );

    \I__1625\ : InMux
    port map (
            O => \N__8029\,
            I => \N__7998\
        );

    \I__1624\ : InMux
    port map (
            O => \N__8028\,
            I => \N__7995\
        );

    \I__1623\ : InMux
    port map (
            O => \N__8027\,
            I => \N__7988\
        );

    \I__1622\ : InMux
    port map (
            O => \N__8026\,
            I => \N__7988\
        );

    \I__1621\ : InMux
    port map (
            O => \N__8025\,
            I => \N__7988\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__8022\,
            I => \N__7981\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__8019\,
            I => \N__7981\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__8016\,
            I => \N__7981\
        );

    \I__1617\ : InMux
    port map (
            O => \N__8015\,
            I => \N__7978\
        );

    \I__1616\ : InMux
    port map (
            O => \N__8012\,
            I => \N__7974\
        );

    \I__1615\ : InMux
    port map (
            O => \N__8011\,
            I => \N__7970\
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__8010\,
            I => \N__7965\
        );

    \I__1613\ : InMux
    port map (
            O => \N__8009\,
            I => \N__7962\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__8006\,
            I => \N__7959\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__8001\,
            I => \N__7956\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__7998\,
            I => \N__7945\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__7995\,
            I => \N__7945\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__7988\,
            I => \N__7945\
        );

    \I__1607\ : Span4Mux_v
    port map (
            O => \N__7981\,
            I => \N__7945\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__7978\,
            I => \N__7945\
        );

    \I__1605\ : InMux
    port map (
            O => \N__7977\,
            I => \N__7939\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__7974\,
            I => \N__7936\
        );

    \I__1603\ : InMux
    port map (
            O => \N__7973\,
            I => \N__7933\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__7970\,
            I => \N__7930\
        );

    \I__1601\ : InMux
    port map (
            O => \N__7969\,
            I => \N__7927\
        );

    \I__1600\ : InMux
    port map (
            O => \N__7968\,
            I => \N__7922\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7965\,
            I => \N__7922\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__7962\,
            I => \N__7919\
        );

    \I__1597\ : Span4Mux_v
    port map (
            O => \N__7959\,
            I => \N__7912\
        );

    \I__1596\ : Span4Mux_h
    port map (
            O => \N__7956\,
            I => \N__7912\
        );

    \I__1595\ : Span4Mux_v
    port map (
            O => \N__7945\,
            I => \N__7912\
        );

    \I__1594\ : InMux
    port map (
            O => \N__7944\,
            I => \N__7905\
        );

    \I__1593\ : InMux
    port map (
            O => \N__7943\,
            I => \N__7905\
        );

    \I__1592\ : InMux
    port map (
            O => \N__7942\,
            I => \N__7905\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__7939\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1590\ : Odrv4
    port map (
            O => \N__7936\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__7933\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1588\ : Odrv4
    port map (
            O => \N__7930\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__7927\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__7922\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1585\ : Odrv12
    port map (
            O => \N__7919\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1584\ : Odrv4
    port map (
            O => \N__7912\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__7905\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1582\ : InMux
    port map (
            O => \N__7886\,
            I => \N__7883\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__7883\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_29_i_a2_i_1_0\
        );

    \I__1580\ : InMux
    port map (
            O => \N__7880\,
            I => \N__7873\
        );

    \I__1579\ : InMux
    port map (
            O => \N__7879\,
            I => \N__7870\
        );

    \I__1578\ : InMux
    port map (
            O => \N__7878\,
            I => \N__7863\
        );

    \I__1577\ : InMux
    port map (
            O => \N__7877\,
            I => \N__7863\
        );

    \I__1576\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7863\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__7873\,
            I => \N__7860\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__7870\,
            I => \N__7855\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__7863\,
            I => \N__7855\
        );

    \I__1572\ : Span4Mux_v
    port map (
            O => \N__7860\,
            I => \N__7840\
        );

    \I__1571\ : Span4Mux_h
    port map (
            O => \N__7855\,
            I => \N__7840\
        );

    \I__1570\ : InMux
    port map (
            O => \N__7854\,
            I => \N__7837\
        );

    \I__1569\ : InMux
    port map (
            O => \N__7853\,
            I => \N__7834\
        );

    \I__1568\ : InMux
    port map (
            O => \N__7852\,
            I => \N__7829\
        );

    \I__1567\ : InMux
    port map (
            O => \N__7851\,
            I => \N__7829\
        );

    \I__1566\ : InMux
    port map (
            O => \N__7850\,
            I => \N__7826\
        );

    \I__1565\ : InMux
    port map (
            O => \N__7849\,
            I => \N__7821\
        );

    \I__1564\ : InMux
    port map (
            O => \N__7848\,
            I => \N__7821\
        );

    \I__1563\ : InMux
    port map (
            O => \N__7847\,
            I => \N__7813\
        );

    \I__1562\ : InMux
    port map (
            O => \N__7846\,
            I => \N__7813\
        );

    \I__1561\ : InMux
    port map (
            O => \N__7845\,
            I => \N__7813\
        );

    \I__1560\ : Span4Mux_h
    port map (
            O => \N__7840\,
            I => \N__7807\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__7837\,
            I => \N__7807\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__7834\,
            I => \N__7798\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__7829\,
            I => \N__7798\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__7826\,
            I => \N__7793\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__7821\,
            I => \N__7793\
        );

    \I__1554\ : CascadeMux
    port map (
            O => \N__7820\,
            I => \N__7787\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__7813\,
            I => \N__7779\
        );

    \I__1552\ : InMux
    port map (
            O => \N__7812\,
            I => \N__7776\
        );

    \I__1551\ : Span4Mux_v
    port map (
            O => \N__7807\,
            I => \N__7773\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7806\,
            I => \N__7766\
        );

    \I__1549\ : InMux
    port map (
            O => \N__7805\,
            I => \N__7766\
        );

    \I__1548\ : InMux
    port map (
            O => \N__7804\,
            I => \N__7766\
        );

    \I__1547\ : InMux
    port map (
            O => \N__7803\,
            I => \N__7763\
        );

    \I__1546\ : Span4Mux_v
    port map (
            O => \N__7798\,
            I => \N__7756\
        );

    \I__1545\ : Span4Mux_v
    port map (
            O => \N__7793\,
            I => \N__7756\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7792\,
            I => \N__7751\
        );

    \I__1543\ : InMux
    port map (
            O => \N__7791\,
            I => \N__7751\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7790\,
            I => \N__7746\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7787\,
            I => \N__7746\
        );

    \I__1540\ : InMux
    port map (
            O => \N__7786\,
            I => \N__7739\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7785\,
            I => \N__7739\
        );

    \I__1538\ : InMux
    port map (
            O => \N__7784\,
            I => \N__7739\
        );

    \I__1537\ : InMux
    port map (
            O => \N__7783\,
            I => \N__7734\
        );

    \I__1536\ : InMux
    port map (
            O => \N__7782\,
            I => \N__7734\
        );

    \I__1535\ : Span4Mux_v
    port map (
            O => \N__7779\,
            I => \N__7731\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__7776\,
            I => \N__7722\
        );

    \I__1533\ : Sp12to4
    port map (
            O => \N__7773\,
            I => \N__7722\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__7766\,
            I => \N__7722\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__7763\,
            I => \N__7722\
        );

    \I__1530\ : InMux
    port map (
            O => \N__7762\,
            I => \N__7717\
        );

    \I__1529\ : InMux
    port map (
            O => \N__7761\,
            I => \N__7717\
        );

    \I__1528\ : Sp12to4
    port map (
            O => \N__7756\,
            I => \N__7706\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7751\,
            I => \N__7706\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__7746\,
            I => \N__7706\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__7739\,
            I => \N__7706\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__7734\,
            I => \N__7706\
        );

    \I__1523\ : Sp12to4
    port map (
            O => \N__7731\,
            I => \N__7699\
        );

    \I__1522\ : Span12Mux_v
    port map (
            O => \N__7722\,
            I => \N__7699\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__7717\,
            I => \N__7699\
        );

    \I__1520\ : Span12Mux_h
    port map (
            O => \N__7706\,
            I => \N__7696\
        );

    \I__1519\ : Span12Mux_h
    port map (
            O => \N__7699\,
            I => \N__7693\
        );

    \I__1518\ : Odrv12
    port map (
            O => \N__7696\,
            I => \RESETn_c\
        );

    \I__1517\ : Odrv12
    port map (
            O => \N__7693\,
            I => \RESETn_c\
        );

    \I__1516\ : IoInMux
    port map (
            O => \N__7688\,
            I => \N__7685\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__7685\,
            I => \N__7682\
        );

    \I__1514\ : Span12Mux_s9_v
    port map (
            O => \N__7682\,
            I => \N__7679\
        );

    \I__1513\ : Odrv12
    port map (
            O => \N__7679\,
            I => \RESETn_c_i\
        );

    \I__1512\ : InMux
    port map (
            O => \N__7676\,
            I => \N__7673\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__7673\,
            I => \N__7670\
        );

    \I__1510\ : Span4Mux_h
    port map (
            O => \N__7670\,
            I => \N__7667\
        );

    \I__1509\ : Sp12to4
    port map (
            O => \N__7667\,
            I => \N__7664\
        );

    \I__1508\ : Odrv12
    port map (
            O => \N__7664\,
            I => \U712_CHIP_RAM.un3_CPU_CYCLE_START\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__7661\,
            I => \N__7658\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7658\,
            I => \N__7653\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7657\,
            I => \N__7650\
        );

    \I__1504\ : InMux
    port map (
            O => \N__7656\,
            I => \N__7647\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7653\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__7650\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__7647\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1500\ : CascadeMux
    port map (
            O => \N__7640\,
            I => \N__7637\
        );

    \I__1499\ : InMux
    port map (
            O => \N__7637\,
            I => \N__7633\
        );

    \I__1498\ : InMux
    port map (
            O => \N__7636\,
            I => \N__7630\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__7633\,
            I => \N__7627\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__7630\,
            I => \N__7624\
        );

    \I__1495\ : Odrv4
    port map (
            O => \N__7627\,
            I => \U712_CHIP_RAM.N_177\
        );

    \I__1494\ : Odrv4
    port map (
            O => \N__7624\,
            I => \U712_CHIP_RAM.N_177\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7619\,
            I => \N__7611\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7618\,
            I => \N__7608\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7617\,
            I => \N__7605\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7616\,
            I => \N__7602\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7615\,
            I => \N__7597\
        );

    \I__1488\ : InMux
    port map (
            O => \N__7614\,
            I => \N__7597\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__7611\,
            I => \N__7594\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__7608\,
            I => \U712_CHIP_RAM.N_172\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__7605\,
            I => \U712_CHIP_RAM.N_172\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__7602\,
            I => \U712_CHIP_RAM.N_172\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7597\,
            I => \U712_CHIP_RAM.N_172\
        );

    \I__1482\ : Odrv4
    port map (
            O => \N__7594\,
            I => \U712_CHIP_RAM.N_172\
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__7583\,
            I => \N__7580\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7580\,
            I => \N__7576\
        );

    \I__1479\ : InMux
    port map (
            O => \N__7579\,
            I => \N__7573\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__7576\,
            I => \N__7570\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__7573\,
            I => \U712_CHIP_RAM.SDRAM_CMD_1_sqmuxa_1_0\
        );

    \I__1476\ : Odrv12
    port map (
            O => \N__7570\,
            I => \U712_CHIP_RAM.SDRAM_CMD_1_sqmuxa_1_0\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7565\,
            I => \N__7561\
        );

    \I__1474\ : InMux
    port map (
            O => \N__7564\,
            I => \N__7555\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__7561\,
            I => \N__7551\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7560\,
            I => \N__7548\
        );

    \I__1471\ : CascadeMux
    port map (
            O => \N__7559\,
            I => \N__7538\
        );

    \I__1470\ : InMux
    port map (
            O => \N__7558\,
            I => \N__7534\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__7555\,
            I => \N__7531\
        );

    \I__1468\ : InMux
    port map (
            O => \N__7554\,
            I => \N__7528\
        );

    \I__1467\ : Span4Mux_h
    port map (
            O => \N__7551\,
            I => \N__7525\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7548\,
            I => \N__7522\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7547\,
            I => \N__7517\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7546\,
            I => \N__7517\
        );

    \I__1463\ : InMux
    port map (
            O => \N__7545\,
            I => \N__7508\
        );

    \I__1462\ : InMux
    port map (
            O => \N__7544\,
            I => \N__7508\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7543\,
            I => \N__7508\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7542\,
            I => \N__7508\
        );

    \I__1459\ : InMux
    port map (
            O => \N__7541\,
            I => \N__7505\
        );

    \I__1458\ : InMux
    port map (
            O => \N__7538\,
            I => \N__7500\
        );

    \I__1457\ : InMux
    port map (
            O => \N__7537\,
            I => \N__7500\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__7534\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1455\ : Odrv4
    port map (
            O => \N__7531\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__7528\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1453\ : Odrv4
    port map (
            O => \N__7525\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1452\ : Odrv4
    port map (
            O => \N__7522\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__7517\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__7508\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__7505\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__7500\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7481\,
            I => \N__7475\
        );

    \I__1446\ : InMux
    port map (
            O => \N__7480\,
            I => \N__7475\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__7475\,
            I => \U712_CHIP_RAM.N_186\
        );

    \I__1444\ : CascadeMux
    port map (
            O => \N__7472\,
            I => \N__7469\
        );

    \I__1443\ : InMux
    port map (
            O => \N__7469\,
            I => \N__7466\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__7466\,
            I => \N__7463\
        );

    \I__1441\ : Odrv4
    port map (
            O => \N__7463\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER34\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__7460\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER34_cascade_\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7457\,
            I => \N__7454\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__7454\,
            I => \N__7451\
        );

    \I__1437\ : Span12Mux_v
    port map (
            O => \N__7451\,
            I => \N__7448\
        );

    \I__1436\ : Span12Mux_h
    port map (
            O => \N__7448\,
            I => \N__7445\
        );

    \I__1435\ : Odrv12
    port map (
            O => \N__7445\,
            I => \A_c_2\
        );

    \I__1434\ : IoInMux
    port map (
            O => \N__7442\,
            I => \N__7439\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__7439\,
            I => \N__7435\
        );

    \I__1432\ : InMux
    port map (
            O => \N__7438\,
            I => \N__7432\
        );

    \I__1431\ : Span12Mux_s4_v
    port map (
            O => \N__7435\,
            I => \N__7427\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__7432\,
            I => \N__7427\
        );

    \I__1429\ : Span12Mux_v
    port map (
            O => \N__7427\,
            I => \N__7424\
        );

    \I__1428\ : Span12Mux_h
    port map (
            O => \N__7424\,
            I => \N__7421\
        );

    \I__1427\ : Odrv12
    port map (
            O => \N__7421\,
            I => \A_c_9\
        );

    \I__1426\ : InMux
    port map (
            O => \N__7418\,
            I => \N__7415\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__7415\,
            I => \N__7412\
        );

    \I__1424\ : Odrv12
    port map (
            O => \N__7412\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER16_2\
        );

    \I__1423\ : InMux
    port map (
            O => \N__7409\,
            I => \N__7405\
        );

    \I__1422\ : InMux
    port map (
            O => \N__7408\,
            I => \N__7402\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__7405\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER17_0\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__7402\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER17_0\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__7397\,
            I => \N__7391\
        );

    \I__1418\ : InMux
    port map (
            O => \N__7396\,
            I => \N__7388\
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__7395\,
            I => \N__7384\
        );

    \I__1416\ : InMux
    port map (
            O => \N__7394\,
            I => \N__7381\
        );

    \I__1415\ : InMux
    port map (
            O => \N__7391\,
            I => \N__7376\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__7388\,
            I => \N__7371\
        );

    \I__1413\ : InMux
    port map (
            O => \N__7387\,
            I => \N__7368\
        );

    \I__1412\ : InMux
    port map (
            O => \N__7384\,
            I => \N__7365\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__7381\,
            I => \N__7362\
        );

    \I__1410\ : InMux
    port map (
            O => \N__7380\,
            I => \N__7359\
        );

    \I__1409\ : InMux
    port map (
            O => \N__7379\,
            I => \N__7356\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__7376\,
            I => \N__7353\
        );

    \I__1407\ : InMux
    port map (
            O => \N__7375\,
            I => \N__7348\
        );

    \I__1406\ : InMux
    port map (
            O => \N__7374\,
            I => \N__7348\
        );

    \I__1405\ : Span4Mux_v
    port map (
            O => \N__7371\,
            I => \N__7343\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__7368\,
            I => \N__7343\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__7365\,
            I => \N__7334\
        );

    \I__1402\ : Span4Mux_h
    port map (
            O => \N__7362\,
            I => \N__7334\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__7359\,
            I => \N__7334\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__7356\,
            I => \N__7334\
        );

    \I__1399\ : Odrv12
    port map (
            O => \N__7353\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__7348\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1397\ : Odrv4
    port map (
            O => \N__7343\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1396\ : Odrv4
    port map (
            O => \N__7334\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1395\ : CascadeMux
    port map (
            O => \N__7325\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER17_0_cascade_\
        );

    \I__1394\ : InMux
    port map (
            O => \N__7322\,
            I => \N__7318\
        );

    \I__1393\ : InMux
    port map (
            O => \N__7321\,
            I => \N__7315\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__7318\,
            I => \U712_CHIP_RAM.N_33\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__7315\,
            I => \U712_CHIP_RAM.N_33\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__7310\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER19_0_cascade_\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__7307\,
            I => \N__7304\
        );

    \I__1388\ : InMux
    port map (
            O => \N__7304\,
            I => \N__7301\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__7301\,
            I => \N__7296\
        );

    \I__1386\ : InMux
    port map (
            O => \N__7300\,
            I => \N__7293\
        );

    \I__1385\ : InMux
    port map (
            O => \N__7299\,
            I => \N__7290\
        );

    \I__1384\ : Odrv12
    port map (
            O => \N__7296\,
            I => \U712_CHIP_RAM.CPU_CYCLE_DISABLEZ0\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__7293\,
            I => \U712_CHIP_RAM.CPU_CYCLE_DISABLEZ0\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__7290\,
            I => \U712_CHIP_RAM.CPU_CYCLE_DISABLEZ0\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7283\,
            I => \N__7280\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7280\,
            I => \N__7277\
        );

    \I__1379\ : Span12Mux_h
    port map (
            O => \N__7277\,
            I => \N__7274\
        );

    \I__1378\ : Odrv12
    port map (
            O => \N__7274\,
            I => \U712_CHIP_RAM.N_95\
        );

    \I__1377\ : CascadeMux
    port map (
            O => \N__7271\,
            I => \N__7264\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7270\,
            I => \N__7261\
        );

    \I__1375\ : InMux
    port map (
            O => \N__7269\,
            I => \N__7258\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7268\,
            I => \N__7252\
        );

    \I__1373\ : InMux
    port map (
            O => \N__7267\,
            I => \N__7252\
        );

    \I__1372\ : InMux
    port map (
            O => \N__7264\,
            I => \N__7249\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__7261\,
            I => \N__7244\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__7258\,
            I => \N__7241\
        );

    \I__1369\ : InMux
    port map (
            O => \N__7257\,
            I => \N__7238\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__7252\,
            I => \N__7233\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__7249\,
            I => \N__7233\
        );

    \I__1366\ : InMux
    port map (
            O => \N__7248\,
            I => \N__7230\
        );

    \I__1365\ : InMux
    port map (
            O => \N__7247\,
            I => \N__7227\
        );

    \I__1364\ : Span4Mux_v
    port map (
            O => \N__7244\,
            I => \N__7220\
        );

    \I__1363\ : Span4Mux_v
    port map (
            O => \N__7241\,
            I => \N__7220\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__7238\,
            I => \N__7220\
        );

    \I__1361\ : Span4Mux_v
    port map (
            O => \N__7233\,
            I => \N__7217\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__7230\,
            I => \U712_CHIP_RAM.N_119\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__7227\,
            I => \U712_CHIP_RAM.N_119\
        );

    \I__1358\ : Odrv4
    port map (
            O => \N__7220\,
            I => \U712_CHIP_RAM.N_119\
        );

    \I__1357\ : Odrv4
    port map (
            O => \N__7217\,
            I => \U712_CHIP_RAM.N_119\
        );

    \I__1356\ : InMux
    port map (
            O => \N__7208\,
            I => \N__7205\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__7205\,
            I => \N__7201\
        );

    \I__1354\ : InMux
    port map (
            O => \N__7204\,
            I => \N__7198\
        );

    \I__1353\ : Span4Mux_h
    port map (
            O => \N__7201\,
            I => \N__7193\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__7198\,
            I => \N__7190\
        );

    \I__1351\ : InMux
    port map (
            O => \N__7197\,
            I => \N__7187\
        );

    \I__1350\ : InMux
    port map (
            O => \N__7196\,
            I => \N__7184\
        );

    \I__1349\ : Odrv4
    port map (
            O => \N__7193\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1348\ : Odrv4
    port map (
            O => \N__7190\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__7187\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__7184\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__7175\,
            I => \U712_CHIP_RAM.N_95_cascade_\
        );

    \I__1344\ : InMux
    port map (
            O => \N__7172\,
            I => \N__7169\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__7169\,
            I => \N__7166\
        );

    \I__1342\ : Span4Mux_h
    port map (
            O => \N__7166\,
            I => \N__7163\
        );

    \I__1341\ : Odrv4
    port map (
            O => \N__7163\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_3_sqmuxa_1\
        );

    \I__1340\ : CascadeMux
    port map (
            O => \N__7160\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_3_sqmuxa_1_cascade_\
        );

    \I__1339\ : CascadeMux
    port map (
            O => \N__7157\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_cascade_\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7154\,
            I => \N__7151\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__7151\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_7\
        );

    \I__1336\ : InMux
    port map (
            O => \N__7148\,
            I => \N__7142\
        );

    \I__1335\ : InMux
    port map (
            O => \N__7147\,
            I => \N__7139\
        );

    \I__1334\ : InMux
    port map (
            O => \N__7146\,
            I => \N__7136\
        );

    \I__1333\ : InMux
    port map (
            O => \N__7145\,
            I => \N__7133\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__7142\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER38_1_0\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__7139\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER38_1_0\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__7136\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER38_1_0\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__7133\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER38_1_0\
        );

    \I__1328\ : InMux
    port map (
            O => \N__7124\,
            I => \N__7121\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__7121\,
            I => \N__7115\
        );

    \I__1326\ : InMux
    port map (
            O => \N__7120\,
            I => \N__7110\
        );

    \I__1325\ : InMux
    port map (
            O => \N__7119\,
            I => \N__7110\
        );

    \I__1324\ : InMux
    port map (
            O => \N__7118\,
            I => \N__7107\
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__7115\,
            I => \U712_CHIP_RAM.N_94\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__7110\,
            I => \U712_CHIP_RAM.N_94\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__7107\,
            I => \U712_CHIP_RAM.N_94\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__7100\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_4_0_cascade_\
        );

    \I__1319\ : InMux
    port map (
            O => \N__7097\,
            I => \N__7094\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__7094\,
            I => \U712_CHIP_RAM.CPU_TACK_7_0\
        );

    \I__1317\ : InMux
    port map (
            O => \N__7091\,
            I => \N__7085\
        );

    \I__1316\ : InMux
    port map (
            O => \N__7090\,
            I => \N__7085\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__7085\,
            I => \N__7081\
        );

    \I__1314\ : InMux
    port map (
            O => \N__7084\,
            I => \N__7077\
        );

    \I__1313\ : Span4Mux_h
    port map (
            O => \N__7081\,
            I => \N__7074\
        );

    \I__1312\ : InMux
    port map (
            O => \N__7080\,
            I => \N__7071\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__7077\,
            I => \CPU_TACKm\
        );

    \I__1310\ : Odrv4
    port map (
            O => \N__7074\,
            I => \CPU_TACKm\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__7071\,
            I => \CPU_TACKm\
        );

    \I__1308\ : InMux
    port map (
            O => \N__7064\,
            I => \N__7061\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__7061\,
            I => \N__7058\
        );

    \I__1306\ : Span12Mux_h
    port map (
            O => \N__7058\,
            I => \N__7055\
        );

    \I__1305\ : Odrv12
    port map (
            O => \N__7055\,
            I => \A_c_7\
        );

    \I__1304\ : InMux
    port map (
            O => \N__7052\,
            I => \N__7049\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__7049\,
            I => \N__7046\
        );

    \I__1302\ : Span12Mux_h
    port map (
            O => \N__7046\,
            I => \N__7043\
        );

    \I__1301\ : Span12Mux_v
    port map (
            O => \N__7043\,
            I => \N__7040\
        );

    \I__1300\ : Odrv12
    port map (
            O => \N__7040\,
            I => \A_c_14\
        );

    \I__1299\ : InMux
    port map (
            O => \N__7037\,
            I => \N__7034\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__7034\,
            I => \U712_CHIP_RAM.N_173\
        );

    \I__1297\ : IoInMux
    port map (
            O => \N__7031\,
            I => \N__7028\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__7028\,
            I => \N__7025\
        );

    \I__1295\ : Span4Mux_s2_v
    port map (
            O => \N__7025\,
            I => \N__7022\
        );

    \I__1294\ : Span4Mux_h
    port map (
            O => \N__7022\,
            I => \N__7019\
        );

    \I__1293\ : Span4Mux_v
    port map (
            O => \N__7019\,
            I => \N__7016\
        );

    \I__1292\ : Odrv4
    port map (
            O => \N__7016\,
            I => \N_56_i\
        );

    \I__1291\ : InMux
    port map (
            O => \N__7013\,
            I => \N__7003\
        );

    \I__1290\ : InMux
    port map (
            O => \N__7012\,
            I => \N__7003\
        );

    \I__1289\ : InMux
    port map (
            O => \N__7011\,
            I => \N__6999\
        );

    \I__1288\ : InMux
    port map (
            O => \N__7010\,
            I => \N__6992\
        );

    \I__1287\ : InMux
    port map (
            O => \N__7009\,
            I => \N__6992\
        );

    \I__1286\ : InMux
    port map (
            O => \N__7008\,
            I => \N__6992\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__7003\,
            I => \N__6989\
        );

    \I__1284\ : CascadeMux
    port map (
            O => \N__7002\,
            I => \N__6986\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__6999\,
            I => \N__6983\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__6992\,
            I => \N__6978\
        );

    \I__1281\ : Span4Mux_v
    port map (
            O => \N__6989\,
            I => \N__6978\
        );

    \I__1280\ : InMux
    port map (
            O => \N__6986\,
            I => \N__6975\
        );

    \I__1279\ : Span4Mux_v
    port map (
            O => \N__6983\,
            I => \N__6972\
        );

    \I__1278\ : Span4Mux_h
    port map (
            O => \N__6978\,
            I => \N__6966\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6975\,
            I => \N__6966\
        );

    \I__1276\ : Span4Mux_v
    port map (
            O => \N__6972\,
            I => \N__6963\
        );

    \I__1275\ : InMux
    port map (
            O => \N__6971\,
            I => \N__6960\
        );

    \I__1274\ : Span4Mux_h
    port map (
            O => \N__6966\,
            I => \N__6957\
        );

    \I__1273\ : Span4Mux_h
    port map (
            O => \N__6963\,
            I => \N__6954\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__6960\,
            I => \N__6951\
        );

    \I__1271\ : Sp12to4
    port map (
            O => \N__6957\,
            I => \N__6948\
        );

    \I__1270\ : Sp12to4
    port map (
            O => \N__6954\,
            I => \N__6943\
        );

    \I__1269\ : Span12Mux_v
    port map (
            O => \N__6951\,
            I => \N__6943\
        );

    \I__1268\ : Span12Mux_v
    port map (
            O => \N__6948\,
            I => \N__6940\
        );

    \I__1267\ : Odrv12
    port map (
            O => \N__6943\,
            I => \SIZ_c_0\
        );

    \I__1266\ : Odrv12
    port map (
            O => \N__6940\,
            I => \SIZ_c_0\
        );

    \I__1265\ : InMux
    port map (
            O => \N__6935\,
            I => \N__6923\
        );

    \I__1264\ : InMux
    port map (
            O => \N__6934\,
            I => \N__6923\
        );

    \I__1263\ : InMux
    port map (
            O => \N__6933\,
            I => \N__6923\
        );

    \I__1262\ : InMux
    port map (
            O => \N__6932\,
            I => \N__6920\
        );

    \I__1261\ : InMux
    port map (
            O => \N__6931\,
            I => \N__6915\
        );

    \I__1260\ : InMux
    port map (
            O => \N__6930\,
            I => \N__6915\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__6923\,
            I => \N__6908\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__6920\,
            I => \N__6908\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__6915\,
            I => \N__6908\
        );

    \I__1256\ : Span4Mux_v
    port map (
            O => \N__6908\,
            I => \N__6905\
        );

    \I__1255\ : Sp12to4
    port map (
            O => \N__6905\,
            I => \N__6902\
        );

    \I__1254\ : Span12Mux_h
    port map (
            O => \N__6902\,
            I => \N__6899\
        );

    \I__1253\ : Odrv12
    port map (
            O => \N__6899\,
            I => \A_c_1\
        );

    \I__1252\ : CascadeMux
    port map (
            O => \N__6896\,
            I => \N__6891\
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__6895\,
            I => \N__6888\
        );

    \I__1250\ : CascadeMux
    port map (
            O => \N__6894\,
            I => \N__6885\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6891\,
            I => \N__6880\
        );

    \I__1248\ : InMux
    port map (
            O => \N__6888\,
            I => \N__6880\
        );

    \I__1247\ : InMux
    port map (
            O => \N__6885\,
            I => \N__6877\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__6880\,
            I => \N__6870\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__6877\,
            I => \N__6870\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__6876\,
            I => \N__6867\
        );

    \I__1243\ : CascadeMux
    port map (
            O => \N__6875\,
            I => \N__6864\
        );

    \I__1242\ : Span4Mux_v
    port map (
            O => \N__6870\,
            I => \N__6859\
        );

    \I__1241\ : InMux
    port map (
            O => \N__6867\,
            I => \N__6852\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6864\,
            I => \N__6852\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6863\,
            I => \N__6852\
        );

    \I__1238\ : InMux
    port map (
            O => \N__6862\,
            I => \N__6849\
        );

    \I__1237\ : Span4Mux_h
    port map (
            O => \N__6859\,
            I => \N__6845\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__6852\,
            I => \N__6842\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6849\,
            I => \N__6839\
        );

    \I__1234\ : InMux
    port map (
            O => \N__6848\,
            I => \N__6836\
        );

    \I__1233\ : Sp12to4
    port map (
            O => \N__6845\,
            I => \N__6827\
        );

    \I__1232\ : Span12Mux_h
    port map (
            O => \N__6842\,
            I => \N__6827\
        );

    \I__1231\ : Sp12to4
    port map (
            O => \N__6839\,
            I => \N__6827\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__6836\,
            I => \N__6827\
        );

    \I__1229\ : Odrv12
    port map (
            O => \N__6827\,
            I => \A_c_0\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__6824\,
            I => \N__6819\
        );

    \I__1227\ : InMux
    port map (
            O => \N__6823\,
            I => \N__6808\
        );

    \I__1226\ : InMux
    port map (
            O => \N__6822\,
            I => \N__6808\
        );

    \I__1225\ : InMux
    port map (
            O => \N__6819\,
            I => \N__6808\
        );

    \I__1224\ : CascadeMux
    port map (
            O => \N__6818\,
            I => \N__6805\
        );

    \I__1223\ : InMux
    port map (
            O => \N__6817\,
            I => \N__6802\
        );

    \I__1222\ : InMux
    port map (
            O => \N__6816\,
            I => \N__6797\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6815\,
            I => \N__6797\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6808\,
            I => \N__6794\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6805\,
            I => \N__6791\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__6802\,
            I => \N__6786\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__6797\,
            I => \N__6786\
        );

    \I__1216\ : Span4Mux_h
    port map (
            O => \N__6794\,
            I => \N__6781\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__6791\,
            I => \N__6781\
        );

    \I__1214\ : Span4Mux_v
    port map (
            O => \N__6786\,
            I => \N__6778\
        );

    \I__1213\ : Span4Mux_h
    port map (
            O => \N__6781\,
            I => \N__6775\
        );

    \I__1212\ : Span4Mux_v
    port map (
            O => \N__6778\,
            I => \N__6771\
        );

    \I__1211\ : Span4Mux_v
    port map (
            O => \N__6775\,
            I => \N__6768\
        );

    \I__1210\ : InMux
    port map (
            O => \N__6774\,
            I => \N__6765\
        );

    \I__1209\ : Span4Mux_h
    port map (
            O => \N__6771\,
            I => \N__6762\
        );

    \I__1208\ : Span4Mux_v
    port map (
            O => \N__6768\,
            I => \N__6759\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__6765\,
            I => \N__6756\
        );

    \I__1206\ : Sp12to4
    port map (
            O => \N__6762\,
            I => \N__6749\
        );

    \I__1205\ : Sp12to4
    port map (
            O => \N__6759\,
            I => \N__6749\
        );

    \I__1204\ : Span12Mux_v
    port map (
            O => \N__6756\,
            I => \N__6749\
        );

    \I__1203\ : Odrv12
    port map (
            O => \N__6749\,
            I => \SIZ_c_1\
        );

    \I__1202\ : IoInMux
    port map (
            O => \N__6746\,
            I => \N__6743\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__6743\,
            I => \N__6740\
        );

    \I__1200\ : Span4Mux_s1_v
    port map (
            O => \N__6740\,
            I => \N__6737\
        );

    \I__1199\ : Span4Mux_h
    port map (
            O => \N__6737\,
            I => \N__6734\
        );

    \I__1198\ : Span4Mux_v
    port map (
            O => \N__6734\,
            I => \N__6731\
        );

    \I__1197\ : Odrv4
    port map (
            O => \N__6731\,
            I => \N_58_i\
        );

    \I__1196\ : IoInMux
    port map (
            O => \N__6728\,
            I => \N__6725\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__6725\,
            I => \N__6722\
        );

    \I__1194\ : IoSpan4Mux
    port map (
            O => \N__6722\,
            I => \N__6719\
        );

    \I__1193\ : IoSpan4Mux
    port map (
            O => \N__6719\,
            I => \N__6716\
        );

    \I__1192\ : Span4Mux_s3_v
    port map (
            O => \N__6716\,
            I => \N__6713\
        );

    \I__1191\ : Odrv4
    port map (
            O => \N__6713\,
            I => \DMA_LATCH_EN_c\
        );

    \I__1190\ : CEMux
    port map (
            O => \N__6710\,
            I => \N__6707\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__6707\,
            I => \N__6704\
        );

    \I__1188\ : Odrv4
    port map (
            O => \N__6704\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_7_0_0\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6701\,
            I => \N__6698\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__6698\,
            I => \N__6695\
        );

    \I__1185\ : Span4Mux_v
    port map (
            O => \N__6695\,
            I => \N__6692\
        );

    \I__1184\ : Sp12to4
    port map (
            O => \N__6692\,
            I => \N__6689\
        );

    \I__1183\ : Span12Mux_h
    port map (
            O => \N__6689\,
            I => \N__6686\
        );

    \I__1182\ : Odrv12
    port map (
            O => \N__6686\,
            I => \A_c_8\
        );

    \I__1181\ : InMux
    port map (
            O => \N__6683\,
            I => \N__6680\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6680\,
            I => \N__6677\
        );

    \I__1179\ : Span12Mux_v
    port map (
            O => \N__6677\,
            I => \N__6674\
        );

    \I__1178\ : Span12Mux_h
    port map (
            O => \N__6674\,
            I => \N__6671\
        );

    \I__1177\ : Odrv12
    port map (
            O => \N__6671\,
            I => \A_c_15\
        );

    \I__1176\ : InMux
    port map (
            O => \N__6668\,
            I => \N__6665\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6665\,
            I => \N__6662\
        );

    \I__1174\ : Span4Mux_v
    port map (
            O => \N__6662\,
            I => \N__6659\
        );

    \I__1173\ : Sp12to4
    port map (
            O => \N__6659\,
            I => \N__6656\
        );

    \I__1172\ : Span12Mux_h
    port map (
            O => \N__6656\,
            I => \N__6653\
        );

    \I__1171\ : Span12Mux_v
    port map (
            O => \N__6653\,
            I => \N__6650\
        );

    \I__1170\ : Odrv12
    port map (
            O => \N__6650\,
            I => \A_c_16\
        );

    \I__1169\ : InMux
    port map (
            O => \N__6647\,
            I => \N__6644\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__6644\,
            I => \N__6641\
        );

    \I__1167\ : Span12Mux_h
    port map (
            O => \N__6641\,
            I => \N__6638\
        );

    \I__1166\ : Span12Mux_v
    port map (
            O => \N__6638\,
            I => \N__6635\
        );

    \I__1165\ : Odrv12
    port map (
            O => \N__6635\,
            I => \A_c_18\
        );

    \I__1164\ : InMux
    port map (
            O => \N__6632\,
            I => \N__6629\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__6629\,
            I => \N__6626\
        );

    \I__1162\ : Span12Mux_v
    port map (
            O => \N__6626\,
            I => \N__6623\
        );

    \I__1161\ : Span12Mux_h
    port map (
            O => \N__6623\,
            I => \N__6620\
        );

    \I__1160\ : Odrv12
    port map (
            O => \N__6620\,
            I => \A_c_13\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6617\,
            I => \N__6614\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__6614\,
            I => \N__6611\
        );

    \I__1157\ : Span4Mux_v
    port map (
            O => \N__6611\,
            I => \N__6608\
        );

    \I__1156\ : Sp12to4
    port map (
            O => \N__6608\,
            I => \N__6605\
        );

    \I__1155\ : Span12Mux_h
    port map (
            O => \N__6605\,
            I => \N__6602\
        );

    \I__1154\ : Odrv12
    port map (
            O => \N__6602\,
            I => \A_c_6\
        );

    \I__1153\ : InMux
    port map (
            O => \N__6599\,
            I => \N__6595\
        );

    \I__1152\ : InMux
    port map (
            O => \N__6598\,
            I => \N__6592\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__6595\,
            I => \U712_CHIP_RAM.CLK_EN_5_0\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__6592\,
            I => \U712_CHIP_RAM.CLK_EN_5_0\
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__6587\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_1_cascade_\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6584\,
            I => \N__6577\
        );

    \I__1147\ : InMux
    port map (
            O => \N__6583\,
            I => \N__6577\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6582\,
            I => \N__6574\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__6577\,
            I => \N__6571\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__6574\,
            I => \U712_CHIP_RAM.N_187\
        );

    \I__1143\ : Odrv4
    port map (
            O => \N__6571\,
            I => \U712_CHIP_RAM.N_187\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6566\,
            I => \N__6563\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__6563\,
            I => \N__6560\
        );

    \I__1140\ : Odrv12
    port map (
            O => \N__6560\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERlde_0_a3_0_0\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6557\,
            I => \N__6553\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6556\,
            I => \N__6550\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__6553\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6550\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0\
        );

    \I__1135\ : CascadeMux
    port map (
            O => \N__6545\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a3_1_1_cascade_\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6542\,
            I => \N__6539\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6539\,
            I => \U712_CHIP_RAM.N_155\
        );

    \I__1132\ : CascadeMux
    port map (
            O => \N__6536\,
            I => \N__6533\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6533\,
            I => \N__6530\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__6530\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a3_1\
        );

    \I__1129\ : CascadeMux
    port map (
            O => \N__6527\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_cascade_\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6524\,
            I => \N__6521\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__6521\,
            I => \N__6518\
        );

    \I__1126\ : Odrv12
    port map (
            O => \N__6518\,
            I => \U712_BYTE_ENABLE.N_58\
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__6515\,
            I => \N__6512\
        );

    \I__1124\ : InMux
    port map (
            O => \N__6512\,
            I => \N__6509\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6509\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_7_2\
        );

    \I__1122\ : CascadeMux
    port map (
            O => \N__6506\,
            I => \U712_CHIP_RAM.BANK0_7_0_cascade_\
        );

    \I__1121\ : IoInMux
    port map (
            O => \N__6503\,
            I => \N__6500\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__6500\,
            I => \N__6497\
        );

    \I__1119\ : IoSpan4Mux
    port map (
            O => \N__6497\,
            I => \N__6494\
        );

    \I__1118\ : Sp12to4
    port map (
            O => \N__6494\,
            I => \N__6491\
        );

    \I__1117\ : Span12Mux_s7_v
    port map (
            O => \N__6491\,
            I => \N__6487\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6490\,
            I => \N__6484\
        );

    \I__1115\ : Odrv12
    port map (
            O => \N__6487\,
            I => \BANK0_c\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__6484\,
            I => \BANK0_c\
        );

    \I__1113\ : InMux
    port map (
            O => \N__6479\,
            I => \N__6476\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__6476\,
            I => \N__6473\
        );

    \I__1111\ : Span4Mux_v
    port map (
            O => \N__6473\,
            I => \N__6470\
        );

    \I__1110\ : Sp12to4
    port map (
            O => \N__6470\,
            I => \N__6467\
        );

    \I__1109\ : Span12Mux_h
    port map (
            O => \N__6467\,
            I => \N__6464\
        );

    \I__1108\ : Odrv12
    port map (
            O => \N__6464\,
            I => \A_c_20\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6461\,
            I => \N__6458\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__6458\,
            I => \U712_CHIP_RAM.A_m_20\
        );

    \I__1105\ : CascadeMux
    port map (
            O => \N__6455\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_\
        );

    \I__1104\ : InMux
    port map (
            O => \N__6452\,
            I => \N__6449\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__6449\,
            I => \N__6445\
        );

    \I__1102\ : InMux
    port map (
            O => \N__6448\,
            I => \N__6442\
        );

    \I__1101\ : Odrv12
    port map (
            O => \N__6445\,
            I => \U712_CHIP_RAM.A_m_2_20\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__6442\,
            I => \U712_CHIP_RAM.A_m_2_20\
        );

    \I__1099\ : CascadeMux
    port map (
            O => \N__6437\,
            I => \U712_CHIP_RAM.N_94_cascade_\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__6434\,
            I => \U712_CHIP_RAM.N_108_cascade_\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__6431\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_i_0_68_i_a3_0_cascade_\
        );

    \I__1096\ : InMux
    port map (
            O => \N__6428\,
            I => \N__6425\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__6425\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_i_0_68_i_0\
        );

    \I__1094\ : CascadeMux
    port map (
            O => \N__6422\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_0_cascade_\
        );

    \I__1093\ : IoInMux
    port map (
            O => \N__6419\,
            I => \N__6416\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__6416\,
            I => \N__6413\
        );

    \I__1091\ : Span12Mux_s10_h
    port map (
            O => \N__6413\,
            I => \N__6410\
        );

    \I__1090\ : Span12Mux_v
    port map (
            O => \N__6410\,
            I => \N__6406\
        );

    \I__1089\ : InMux
    port map (
            O => \N__6409\,
            I => \N__6403\
        );

    \I__1088\ : Odrv12
    port map (
            O => \N__6406\,
            I => \CLK_EN_c\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__6403\,
            I => \CLK_EN_c\
        );

    \I__1086\ : InMux
    port map (
            O => \N__6398\,
            I => \N__6395\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__6395\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_0_0\
        );

    \I__1084\ : InMux
    port map (
            O => \N__6392\,
            I => \N__6387\
        );

    \I__1083\ : InMux
    port map (
            O => \N__6391\,
            I => \N__6384\
        );

    \I__1082\ : InMux
    port map (
            O => \N__6390\,
            I => \N__6381\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__6387\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__6384\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__6381\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1078\ : InMux
    port map (
            O => \N__6374\,
            I => \N__6369\
        );

    \I__1077\ : InMux
    port map (
            O => \N__6373\,
            I => \N__6366\
        );

    \I__1076\ : InMux
    port map (
            O => \N__6372\,
            I => \N__6363\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__6369\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__6366\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__6363\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1072\ : CascadeMux
    port map (
            O => \N__6356\,
            I => \N__6351\
        );

    \I__1071\ : CascadeMux
    port map (
            O => \N__6355\,
            I => \N__6348\
        );

    \I__1070\ : InMux
    port map (
            O => \N__6354\,
            I => \N__6345\
        );

    \I__1069\ : InMux
    port map (
            O => \N__6351\,
            I => \N__6342\
        );

    \I__1068\ : InMux
    port map (
            O => \N__6348\,
            I => \N__6339\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__6345\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__6342\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__6339\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6332\,
            I => \N__6327\
        );

    \I__1063\ : InMux
    port map (
            O => \N__6331\,
            I => \N__6324\
        );

    \I__1062\ : InMux
    port map (
            O => \N__6330\,
            I => \N__6321\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__6327\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__6324\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__6321\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1058\ : CascadeMux
    port map (
            O => \N__6314\,
            I => \U712_CHIP_RAM.N_331_3_cascade_\
        );

    \I__1057\ : CascadeMux
    port map (
            O => \N__6311\,
            I => \N__6307\
        );

    \I__1056\ : InMux
    port map (
            O => \N__6310\,
            I => \N__6301\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6307\,
            I => \N__6301\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6306\,
            I => \N__6298\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__6301\,
            I => \N__6295\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6298\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER37_0_a3_1_0\
        );

    \I__1051\ : Odrv4
    port map (
            O => \N__6295\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER37_0_a3_1_0\
        );

    \I__1050\ : CascadeMux
    port map (
            O => \N__6290\,
            I => \U712_CHIP_RAM.LATCH_CLK_0_sqmuxa_cascade_\
        );

    \I__1049\ : CascadeMux
    port map (
            O => \N__6287\,
            I => \N__6284\
        );

    \I__1048\ : InMux
    port map (
            O => \N__6284\,
            I => \N__6277\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6283\,
            I => \N__6277\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6282\,
            I => \N__6274\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__6277\,
            I => \N__6270\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__6274\,
            I => \N__6267\
        );

    \I__1043\ : InMux
    port map (
            O => \N__6273\,
            I => \N__6264\
        );

    \I__1042\ : Span4Mux_v
    port map (
            O => \N__6270\,
            I => \N__6259\
        );

    \I__1041\ : Span4Mux_h
    port map (
            O => \N__6267\,
            I => \N__6259\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__6264\,
            I => \REG_TACK\
        );

    \I__1039\ : Odrv4
    port map (
            O => \N__6259\,
            I => \REG_TACK\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6254\,
            I => \N__6251\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__6251\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1036\ : InMux
    port map (
            O => \N__6248\,
            I => \N__6245\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__6245\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_7_0\
        );

    \I__1034\ : CascadeMux
    port map (
            O => \N__6242\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_7_0_cascade_\
        );

    \I__1033\ : InMux
    port map (
            O => \N__6239\,
            I => \N__6236\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__6236\,
            I => \N__6232\
        );

    \I__1031\ : InMux
    port map (
            O => \N__6235\,
            I => \N__6229\
        );

    \I__1030\ : Span4Mux_v
    port map (
            O => \N__6232\,
            I => \N__6226\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6229\,
            I => \N__6223\
        );

    \I__1028\ : Span4Mux_h
    port map (
            O => \N__6226\,
            I => \N__6220\
        );

    \I__1027\ : Span12Mux_h
    port map (
            O => \N__6223\,
            I => \N__6215\
        );

    \I__1026\ : Sp12to4
    port map (
            O => \N__6220\,
            I => \N__6215\
        );

    \I__1025\ : Span12Mux_v
    port map (
            O => \N__6215\,
            I => \N__6212\
        );

    \I__1024\ : Odrv12
    port map (
            O => \N__6212\,
            I => \AWEn_c\
        );

    \I__1023\ : InMux
    port map (
            O => \N__6209\,
            I => \N__6206\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__6206\,
            I => \N__6202\
        );

    \I__1021\ : InMux
    port map (
            O => \N__6205\,
            I => \N__6199\
        );

    \I__1020\ : Span4Mux_h
    port map (
            O => \N__6202\,
            I => \N__6193\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__6199\,
            I => \N__6190\
        );

    \I__1018\ : InMux
    port map (
            O => \N__6198\,
            I => \N__6183\
        );

    \I__1017\ : InMux
    port map (
            O => \N__6197\,
            I => \N__6183\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6196\,
            I => \N__6183\
        );

    \I__1015\ : Span4Mux_h
    port map (
            O => \N__6193\,
            I => \N__6180\
        );

    \I__1014\ : Span4Mux_v
    port map (
            O => \N__6190\,
            I => \N__6175\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__6183\,
            I => \N__6175\
        );

    \I__1012\ : Odrv4
    port map (
            O => \N__6180\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1011\ : Odrv4
    port map (
            O => \N__6175\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6170\,
            I => \N__6167\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__6167\,
            I => \N__6164\
        );

    \I__1008\ : Odrv4
    port map (
            O => \N__6164\,
            I => \U712_CHIP_RAM.N_152\
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__6161\,
            I => \N__6158\
        );

    \I__1006\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6154\
        );

    \I__1005\ : CascadeMux
    port map (
            O => \N__6157\,
            I => \N__6148\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__6154\,
            I => \N__6145\
        );

    \I__1003\ : InMux
    port map (
            O => \N__6153\,
            I => \N__6142\
        );

    \I__1002\ : InMux
    port map (
            O => \N__6152\,
            I => \N__6139\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6151\,
            I => \N__6136\
        );

    \I__1000\ : InMux
    port map (
            O => \N__6148\,
            I => \N__6133\
        );

    \I__999\ : Span4Mux_v
    port map (
            O => \N__6145\,
            I => \N__6128\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__6142\,
            I => \N__6128\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__6139\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__6136\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__6133\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__6128\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__993\ : InMux
    port map (
            O => \N__6119\,
            I => \N__6114\
        );

    \I__992\ : InMux
    port map (
            O => \N__6118\,
            I => \N__6109\
        );

    \I__991\ : InMux
    port map (
            O => \N__6117\,
            I => \N__6109\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__6114\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__6109\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__988\ : CascadeMux
    port map (
            O => \N__6104\,
            I => \N__6101\
        );

    \I__987\ : InMux
    port map (
            O => \N__6101\,
            I => \N__6095\
        );

    \I__986\ : InMux
    port map (
            O => \N__6100\,
            I => \N__6095\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__6095\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__984\ : InMux
    port map (
            O => \N__6092\,
            I => \N__6089\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__6089\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\
        );

    \I__982\ : InMux
    port map (
            O => \N__6086\,
            I => \N__6082\
        );

    \I__981\ : InMux
    port map (
            O => \N__6085\,
            I => \N__6079\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__6082\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__6079\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__978\ : CascadeMux
    port map (
            O => \N__6074\,
            I => \N__6069\
        );

    \I__977\ : InMux
    port map (
            O => \N__6073\,
            I => \N__6066\
        );

    \I__976\ : InMux
    port map (
            O => \N__6072\,
            I => \N__6062\
        );

    \I__975\ : InMux
    port map (
            O => \N__6069\,
            I => \N__6059\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__6066\,
            I => \N__6056\
        );

    \I__973\ : InMux
    port map (
            O => \N__6065\,
            I => \N__6053\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__6062\,
            I => \N__6048\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__6059\,
            I => \N__6048\
        );

    \I__970\ : Span4Mux_h
    port map (
            O => \N__6056\,
            I => \N__6045\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__6053\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__968\ : Odrv4
    port map (
            O => \N__6048\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__967\ : Odrv4
    port map (
            O => \N__6045\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__966\ : InMux
    port map (
            O => \N__6038\,
            I => \N__6029\
        );

    \I__965\ : InMux
    port map (
            O => \N__6037\,
            I => \N__6029\
        );

    \I__964\ : InMux
    port map (
            O => \N__6036\,
            I => \N__6029\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__6029\,
            I => \N__6026\
        );

    \I__962\ : Odrv4
    port map (
            O => \N__6026\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__961\ : SRMux
    port map (
            O => \N__6023\,
            I => \N__6020\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__6020\,
            I => \N__6017\
        );

    \I__959\ : Odrv4
    port map (
            O => \N__6017\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__958\ : IoInMux
    port map (
            O => \N__6014\,
            I => \N__6011\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__6011\,
            I => \N__6008\
        );

    \I__956\ : IoSpan4Mux
    port map (
            O => \N__6008\,
            I => \N__6005\
        );

    \I__955\ : Span4Mux_s3_h
    port map (
            O => \N__6005\,
            I => \N__6002\
        );

    \I__954\ : Sp12to4
    port map (
            O => \N__6002\,
            I => \N__5999\
        );

    \I__953\ : Span12Mux_h
    port map (
            O => \N__5999\,
            I => \N__5996\
        );

    \I__952\ : Odrv12
    port map (
            O => \N__5996\,
            I => \CLMBEn_c\
        );

    \I__951\ : InMux
    port map (
            O => \N__5993\,
            I => \N__5990\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__5990\,
            I => \N__5987\
        );

    \I__949\ : Span4Mux_h
    port map (
            O => \N__5987\,
            I => \N__5984\
        );

    \I__948\ : Odrv4
    port map (
            O => \N__5984\,
            I => \U712_CHIP_RAM.LATCH_CLK_0_sqmuxa\
        );

    \I__947\ : InMux
    port map (
            O => \N__5981\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__946\ : InMux
    port map (
            O => \N__5978\,
            I => \N__5975\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__5975\,
            I => \N__5972\
        );

    \I__944\ : Odrv4
    port map (
            O => \N__5972\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__943\ : InMux
    port map (
            O => \N__5969\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__942\ : InMux
    port map (
            O => \N__5966\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__941\ : InMux
    port map (
            O => \N__5963\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__940\ : InMux
    port map (
            O => \N__5960\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__939\ : InMux
    port map (
            O => \N__5957\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__938\ : InMux
    port map (
            O => \N__5954\,
            I => \N__5941\
        );

    \I__937\ : InMux
    port map (
            O => \N__5953\,
            I => \N__5941\
        );

    \I__936\ : InMux
    port map (
            O => \N__5952\,
            I => \N__5941\
        );

    \I__935\ : InMux
    port map (
            O => \N__5951\,
            I => \N__5938\
        );

    \I__934\ : InMux
    port map (
            O => \N__5950\,
            I => \N__5931\
        );

    \I__933\ : InMux
    port map (
            O => \N__5949\,
            I => \N__5931\
        );

    \I__932\ : InMux
    port map (
            O => \N__5948\,
            I => \N__5931\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__5941\,
            I => \U712_CHIP_RAM.N_64\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__5938\,
            I => \U712_CHIP_RAM.N_64\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__5931\,
            I => \U712_CHIP_RAM.N_64\
        );

    \I__928\ : InMux
    port map (
            O => \N__5924\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__927\ : CEMux
    port map (
            O => \N__5921\,
            I => \N__5917\
        );

    \I__926\ : CEMux
    port map (
            O => \N__5920\,
            I => \N__5914\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__5917\,
            I => \N__5911\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__5914\,
            I => \N__5908\
        );

    \I__923\ : Odrv4
    port map (
            O => \N__5911\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__922\ : Odrv12
    port map (
            O => \N__5908\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__5903\,
            I => \N__5898\
        );

    \I__920\ : InMux
    port map (
            O => \N__5902\,
            I => \N__5895\
        );

    \I__919\ : InMux
    port map (
            O => \N__5901\,
            I => \N__5892\
        );

    \I__918\ : InMux
    port map (
            O => \N__5898\,
            I => \N__5889\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__5895\,
            I => \N__5885\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__5892\,
            I => \N__5880\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__5889\,
            I => \N__5880\
        );

    \I__914\ : InMux
    port map (
            O => \N__5888\,
            I => \N__5877\
        );

    \I__913\ : Span4Mux_v
    port map (
            O => \N__5885\,
            I => \N__5874\
        );

    \I__912\ : Span4Mux_v
    port map (
            O => \N__5880\,
            I => \N__5871\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__5877\,
            I => \N__5868\
        );

    \I__910\ : Span4Mux_v
    port map (
            O => \N__5874\,
            I => \N__5865\
        );

    \I__909\ : Span4Mux_v
    port map (
            O => \N__5871\,
            I => \N__5862\
        );

    \I__908\ : Span4Mux_h
    port map (
            O => \N__5868\,
            I => \N__5859\
        );

    \I__907\ : Sp12to4
    port map (
            O => \N__5865\,
            I => \N__5856\
        );

    \I__906\ : Sp12to4
    port map (
            O => \N__5862\,
            I => \N__5853\
        );

    \I__905\ : Sp12to4
    port map (
            O => \N__5859\,
            I => \N__5850\
        );

    \I__904\ : Span12Mux_h
    port map (
            O => \N__5856\,
            I => \N__5843\
        );

    \I__903\ : Span12Mux_h
    port map (
            O => \N__5853\,
            I => \N__5843\
        );

    \I__902\ : Span12Mux_v
    port map (
            O => \N__5850\,
            I => \N__5843\
        );

    \I__901\ : Odrv12
    port map (
            O => \N__5843\,
            I => \CLK40_PLL_i\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__5840\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER33_1_0_cascade_\
        );

    \I__899\ : CascadeMux
    port map (
            O => \N__5837\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_i_0_68_i_2_cascade_\
        );

    \I__898\ : CascadeMux
    port map (
            O => \N__5834\,
            I => \U712_CHIP_RAM.N_64_cascade_\
        );

    \I__897\ : IoInMux
    port map (
            O => \N__5831\,
            I => \N__5828\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__5828\,
            I => \N__5824\
        );

    \I__895\ : InMux
    port map (
            O => \N__5827\,
            I => \N__5821\
        );

    \I__894\ : Span12Mux_s7_v
    port map (
            O => \N__5824\,
            I => \N__5818\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__5821\,
            I => \N__5815\
        );

    \I__892\ : Odrv12
    port map (
            O => \N__5818\,
            I => \CONSTANT_ONE_NET\
        );

    \I__891\ : Odrv12
    port map (
            O => \N__5815\,
            I => \CONSTANT_ONE_NET\
        );

    \I__890\ : InMux
    port map (
            O => \N__5810\,
            I => \N__5807\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__5807\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0\
        );

    \I__888\ : InMux
    port map (
            O => \N__5804\,
            I => \N__5799\
        );

    \I__887\ : InMux
    port map (
            O => \N__5803\,
            I => \N__5794\
        );

    \I__886\ : InMux
    port map (
            O => \N__5802\,
            I => \N__5794\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5799\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER18\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__5794\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER18\
        );

    \I__883\ : InMux
    port map (
            O => \N__5789\,
            I => \N__5786\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__5786\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_1\
        );

    \I__881\ : InMux
    port map (
            O => \N__5783\,
            I => \N__5780\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__5780\,
            I => \U712_CHIP_RAM.LATCH_CLK_6\
        );

    \I__879\ : InMux
    port map (
            O => \N__5777\,
            I => \N__5773\
        );

    \I__878\ : InMux
    port map (
            O => \N__5776\,
            I => \N__5770\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5773\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__5770\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__875\ : InMux
    port map (
            O => \N__5765\,
            I => \N__5761\
        );

    \I__874\ : InMux
    port map (
            O => \N__5764\,
            I => \N__5758\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__5761\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__5758\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__871\ : InMux
    port map (
            O => \N__5753\,
            I => \N__5749\
        );

    \I__870\ : InMux
    port map (
            O => \N__5752\,
            I => \N__5746\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__5749\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__5746\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__867\ : InMux
    port map (
            O => \N__5741\,
            I => \N__5737\
        );

    \I__866\ : InMux
    port map (
            O => \N__5740\,
            I => \N__5734\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__5737\,
            I => \U712_CHIP_RAM.N_9\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__5734\,
            I => \U712_CHIP_RAM.N_9\
        );

    \I__863\ : InMux
    port map (
            O => \N__5729\,
            I => \N__5723\
        );

    \I__862\ : InMux
    port map (
            O => \N__5728\,
            I => \N__5720\
        );

    \I__861\ : InMux
    port map (
            O => \N__5727\,
            I => \N__5717\
        );

    \I__860\ : InMux
    port map (
            O => \N__5726\,
            I => \N__5714\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__5723\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5720\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__5717\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__5714\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__855\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5701\
        );

    \I__854\ : InMux
    port map (
            O => \N__5704\,
            I => \N__5698\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5701\,
            I => \N__5695\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__5698\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__851\ : Odrv4
    port map (
            O => \N__5695\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__850\ : InMux
    port map (
            O => \N__5690\,
            I => \N__5687\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__5687\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\
        );

    \I__848\ : InMux
    port map (
            O => \N__5684\,
            I => \N__5681\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__5681\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__5678\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER18_cascade_\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__5675\,
            I => \N__5672\
        );

    \I__844\ : InMux
    port map (
            O => \N__5672\,
            I => \N__5666\
        );

    \I__843\ : InMux
    port map (
            O => \N__5671\,
            I => \N__5661\
        );

    \I__842\ : InMux
    port map (
            O => \N__5670\,
            I => \N__5661\
        );

    \I__841\ : InMux
    port map (
            O => \N__5669\,
            I => \N__5658\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__5666\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__5661\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__5658\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__837\ : InMux
    port map (
            O => \N__5651\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__836\ : InMux
    port map (
            O => \N__5648\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__835\ : InMux
    port map (
            O => \N__5645\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__834\ : InMux
    port map (
            O => \N__5642\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__833\ : InMux
    port map (
            O => \N__5639\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__832\ : InMux
    port map (
            O => \N__5636\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__831\ : InMux
    port map (
            O => \N__5633\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__830\ : ClkMux
    port map (
            O => \N__5630\,
            I => \N__5603\
        );

    \I__829\ : ClkMux
    port map (
            O => \N__5629\,
            I => \N__5603\
        );

    \I__828\ : ClkMux
    port map (
            O => \N__5628\,
            I => \N__5603\
        );

    \I__827\ : ClkMux
    port map (
            O => \N__5627\,
            I => \N__5603\
        );

    \I__826\ : ClkMux
    port map (
            O => \N__5626\,
            I => \N__5603\
        );

    \I__825\ : ClkMux
    port map (
            O => \N__5625\,
            I => \N__5603\
        );

    \I__824\ : ClkMux
    port map (
            O => \N__5624\,
            I => \N__5603\
        );

    \I__823\ : ClkMux
    port map (
            O => \N__5623\,
            I => \N__5603\
        );

    \I__822\ : ClkMux
    port map (
            O => \N__5622\,
            I => \N__5603\
        );

    \I__821\ : GlobalMux
    port map (
            O => \N__5603\,
            I => \N__5600\
        );

    \I__820\ : gio2CtrlBuf
    port map (
            O => \N__5600\,
            I => \C1_c_g\
        );

    \I__819\ : InMux
    port map (
            O => \N__5597\,
            I => \N__5593\
        );

    \I__818\ : InMux
    port map (
            O => \N__5596\,
            I => \N__5590\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__5593\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__5590\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__815\ : InMux
    port map (
            O => \N__5585\,
            I => \N__5581\
        );

    \I__814\ : InMux
    port map (
            O => \N__5584\,
            I => \N__5578\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5581\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5578\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__811\ : CascadeMux
    port map (
            O => \N__5573\,
            I => \N__5569\
        );

    \I__810\ : InMux
    port map (
            O => \N__5572\,
            I => \N__5566\
        );

    \I__809\ : InMux
    port map (
            O => \N__5569\,
            I => \N__5563\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__5566\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__5563\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__806\ : InMux
    port map (
            O => \N__5558\,
            I => \N__5554\
        );

    \I__805\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5551\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__5554\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5551\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__802\ : InMux
    port map (
            O => \N__5546\,
            I => \N__5543\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__5543\,
            I => \U712_CHIP_RAM.DMA_CYCLE_START_2_0\
        );

    \I__800\ : InMux
    port map (
            O => \N__5540\,
            I => \N__5537\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__5537\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_3\
        );

    \I__798\ : CascadeMux
    port map (
            O => \N__5534\,
            I => \N__5527\
        );

    \I__797\ : CascadeMux
    port map (
            O => \N__5533\,
            I => \N__5518\
        );

    \I__796\ : InMux
    port map (
            O => \N__5532\,
            I => \N__5514\
        );

    \I__795\ : InMux
    port map (
            O => \N__5531\,
            I => \N__5509\
        );

    \I__794\ : InMux
    port map (
            O => \N__5530\,
            I => \N__5506\
        );

    \I__793\ : InMux
    port map (
            O => \N__5527\,
            I => \N__5501\
        );

    \I__792\ : InMux
    port map (
            O => \N__5526\,
            I => \N__5501\
        );

    \I__791\ : InMux
    port map (
            O => \N__5525\,
            I => \N__5496\
        );

    \I__790\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5496\
        );

    \I__789\ : InMux
    port map (
            O => \N__5523\,
            I => \N__5489\
        );

    \I__788\ : InMux
    port map (
            O => \N__5522\,
            I => \N__5489\
        );

    \I__787\ : InMux
    port map (
            O => \N__5521\,
            I => \N__5489\
        );

    \I__786\ : InMux
    port map (
            O => \N__5518\,
            I => \N__5485\
        );

    \I__785\ : InMux
    port map (
            O => \N__5517\,
            I => \N__5482\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__5514\,
            I => \N__5479\
        );

    \I__783\ : InMux
    port map (
            O => \N__5513\,
            I => \N__5474\
        );

    \I__782\ : InMux
    port map (
            O => \N__5512\,
            I => \N__5474\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__5509\,
            I => \N__5471\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__5506\,
            I => \N__5466\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5501\,
            I => \N__5466\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__5496\,
            I => \N__5461\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__5489\,
            I => \N__5461\
        );

    \I__776\ : InMux
    port map (
            O => \N__5488\,
            I => \N__5458\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5485\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__5482\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__773\ : Odrv4
    port map (
            O => \N__5479\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__5474\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__771\ : Odrv4
    port map (
            O => \N__5471\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__770\ : Odrv12
    port map (
            O => \N__5466\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__769\ : Odrv4
    port map (
            O => \N__5461\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__5458\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__767\ : IoInMux
    port map (
            O => \N__5441\,
            I => \N__5438\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__5438\,
            I => \N__5435\
        );

    \I__765\ : Span4Mux_s2_v
    port map (
            O => \N__5435\,
            I => \N__5432\
        );

    \I__764\ : Span4Mux_h
    port map (
            O => \N__5432\,
            I => \N__5429\
        );

    \I__763\ : Span4Mux_h
    port map (
            O => \N__5429\,
            I => \N__5426\
        );

    \I__762\ : Sp12to4
    port map (
            O => \N__5426\,
            I => \N__5423\
        );

    \I__761\ : Span12Mux_s10_v
    port map (
            O => \N__5423\,
            I => \N__5420\
        );

    \I__760\ : Odrv12
    port map (
            O => \N__5420\,
            I => \ASn_c\
        );

    \I__759\ : CEMux
    port map (
            O => \N__5417\,
            I => \N__5414\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5414\,
            I => \N__5411\
        );

    \I__757\ : Span4Mux_v
    port map (
            O => \N__5411\,
            I => \N__5408\
        );

    \I__756\ : Odrv4
    port map (
            O => \N__5408\,
            I => \U712_REG_SM.N_163_0\
        );

    \I__755\ : InMux
    port map (
            O => \N__5405\,
            I => \N__5402\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__5402\,
            I => \N__5398\
        );

    \I__753\ : InMux
    port map (
            O => \N__5401\,
            I => \N__5395\
        );

    \I__752\ : Span4Mux_v
    port map (
            O => \N__5398\,
            I => \N__5392\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__5395\,
            I => \N__5389\
        );

    \I__750\ : Span4Mux_v
    port map (
            O => \N__5392\,
            I => \N__5384\
        );

    \I__749\ : Span4Mux_h
    port map (
            O => \N__5389\,
            I => \N__5384\
        );

    \I__748\ : Span4Mux_v
    port map (
            O => \N__5384\,
            I => \N__5381\
        );

    \I__747\ : IoSpan4Mux
    port map (
            O => \N__5381\,
            I => \N__5378\
        );

    \I__746\ : Odrv4
    port map (
            O => \N__5378\,
            I => \TSn_c\
        );

    \I__745\ : InMux
    port map (
            O => \N__5375\,
            I => \N__5372\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__5372\,
            I => \N__5368\
        );

    \I__743\ : IoInMux
    port map (
            O => \N__5371\,
            I => \N__5365\
        );

    \I__742\ : Span4Mux_h
    port map (
            O => \N__5368\,
            I => \N__5362\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__5365\,
            I => \N__5359\
        );

    \I__740\ : Span4Mux_v
    port map (
            O => \N__5362\,
            I => \N__5356\
        );

    \I__739\ : IoSpan4Mux
    port map (
            O => \N__5359\,
            I => \N__5353\
        );

    \I__738\ : Odrv4
    port map (
            O => \N__5356\,
            I => \RAMENn_c\
        );

    \I__737\ : Odrv4
    port map (
            O => \N__5353\,
            I => \RAMENn_c\
        );

    \I__736\ : IoInMux
    port map (
            O => \N__5348\,
            I => \N__5345\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__5345\,
            I => \N__5342\
        );

    \I__734\ : Span4Mux_s3_v
    port map (
            O => \N__5342\,
            I => \N__5339\
        );

    \I__733\ : Span4Mux_v
    port map (
            O => \N__5339\,
            I => \N__5336\
        );

    \I__732\ : Span4Mux_v
    port map (
            O => \N__5336\,
            I => \N__5333\
        );

    \I__731\ : Odrv4
    port map (
            O => \N__5333\,
            I => \VBENn_c\
        );

    \I__730\ : InMux
    port map (
            O => \N__5330\,
            I => \N__5327\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__5327\,
            I => \U712_CYCLE_TERM.N_47_0\
        );

    \I__728\ : IoInMux
    port map (
            O => \N__5324\,
            I => \N__5320\
        );

    \I__727\ : IoInMux
    port map (
            O => \N__5323\,
            I => \N__5316\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5320\,
            I => \N__5313\
        );

    \I__725\ : IoInMux
    port map (
            O => \N__5319\,
            I => \N__5310\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__5316\,
            I => \N__5307\
        );

    \I__723\ : IoSpan4Mux
    port map (
            O => \N__5313\,
            I => \N__5304\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__5310\,
            I => \N__5301\
        );

    \I__721\ : IoSpan4Mux
    port map (
            O => \N__5307\,
            I => \N__5298\
        );

    \I__720\ : IoSpan4Mux
    port map (
            O => \N__5304\,
            I => \N__5295\
        );

    \I__719\ : IoSpan4Mux
    port map (
            O => \N__5301\,
            I => \N__5292\
        );

    \I__718\ : Sp12to4
    port map (
            O => \N__5298\,
            I => \N__5289\
        );

    \I__717\ : Span4Mux_s2_h
    port map (
            O => \N__5295\,
            I => \N__5286\
        );

    \I__716\ : IoSpan4Mux
    port map (
            O => \N__5292\,
            I => \N__5283\
        );

    \I__715\ : Span12Mux_s9_v
    port map (
            O => \N__5289\,
            I => \N__5280\
        );

    \I__714\ : Sp12to4
    port map (
            O => \N__5286\,
            I => \N__5277\
        );

    \I__713\ : Sp12to4
    port map (
            O => \N__5283\,
            I => \N__5274\
        );

    \I__712\ : Span12Mux_h
    port map (
            O => \N__5280\,
            I => \N__5266\
        );

    \I__711\ : Span12Mux_h
    port map (
            O => \N__5277\,
            I => \N__5266\
        );

    \I__710\ : Span12Mux_s9_v
    port map (
            O => \N__5274\,
            I => \N__5266\
        );

    \I__709\ : InMux
    port map (
            O => \N__5273\,
            I => \N__5263\
        );

    \I__708\ : Odrv12
    port map (
            O => \N__5266\,
            I => \TACK_EN\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__5263\,
            I => \TACK_EN\
        );

    \I__706\ : IoInMux
    port map (
            O => \N__5258\,
            I => \N__5254\
        );

    \I__705\ : IoInMux
    port map (
            O => \N__5257\,
            I => \N__5250\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__5254\,
            I => \N__5247\
        );

    \I__703\ : IoInMux
    port map (
            O => \N__5253\,
            I => \N__5244\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5250\,
            I => \N__5241\
        );

    \I__701\ : Span4Mux_s1_v
    port map (
            O => \N__5247\,
            I => \N__5238\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__5244\,
            I => \N__5235\
        );

    \I__699\ : IoSpan4Mux
    port map (
            O => \N__5241\,
            I => \N__5232\
        );

    \I__698\ : Sp12to4
    port map (
            O => \N__5238\,
            I => \N__5229\
        );

    \I__697\ : Span4Mux_s2_h
    port map (
            O => \N__5235\,
            I => \N__5226\
        );

    \I__696\ : Span4Mux_s0_v
    port map (
            O => \N__5232\,
            I => \N__5223\
        );

    \I__695\ : Span12Mux_h
    port map (
            O => \N__5229\,
            I => \N__5220\
        );

    \I__694\ : Sp12to4
    port map (
            O => \N__5226\,
            I => \N__5217\
        );

    \I__693\ : Sp12to4
    port map (
            O => \N__5223\,
            I => \N__5214\
        );

    \I__692\ : Span12Mux_v
    port map (
            O => \N__5220\,
            I => \N__5206\
        );

    \I__691\ : Span12Mux_v
    port map (
            O => \N__5217\,
            I => \N__5206\
        );

    \I__690\ : Span12Mux_v
    port map (
            O => \N__5214\,
            I => \N__5206\
        );

    \I__689\ : InMux
    port map (
            O => \N__5213\,
            I => \N__5203\
        );

    \I__688\ : Odrv12
    port map (
            O => \N__5206\,
            I => \TACK_OUTn\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__5203\,
            I => \TACK_OUTn\
        );

    \I__686\ : InMux
    port map (
            O => \N__5198\,
            I => \bfn_10_9_0_\
        );

    \I__685\ : InMux
    port map (
            O => \N__5195\,
            I => \N__5191\
        );

    \I__684\ : InMux
    port map (
            O => \N__5194\,
            I => \N__5188\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__5191\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_5\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__5188\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_5\
        );

    \I__681\ : InMux
    port map (
            O => \N__5183\,
            I => \N__5179\
        );

    \I__680\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5176\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__5179\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_6\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__5176\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_6\
        );

    \I__677\ : InMux
    port map (
            O => \N__5171\,
            I => \N__5167\
        );

    \I__676\ : InMux
    port map (
            O => \N__5170\,
            I => \N__5164\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__5167\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_7\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__5164\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_7\
        );

    \I__673\ : CascadeMux
    port map (
            O => \N__5159\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_0_cascade_\
        );

    \I__672\ : IoInMux
    port map (
            O => \N__5156\,
            I => \N__5153\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__5153\,
            I => \N__5150\
        );

    \I__670\ : IoSpan4Mux
    port map (
            O => \N__5150\,
            I => \N__5147\
        );

    \I__669\ : IoSpan4Mux
    port map (
            O => \N__5147\,
            I => \N__5144\
        );

    \I__668\ : Span4Mux_s3_v
    port map (
            O => \N__5144\,
            I => \N__5141\
        );

    \I__667\ : Sp12to4
    port map (
            O => \N__5141\,
            I => \N__5137\
        );

    \I__666\ : InMux
    port map (
            O => \N__5140\,
            I => \N__5134\
        );

    \I__665\ : Odrv12
    port map (
            O => \N__5137\,
            I => \LATCH_CLK_c\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__5134\,
            I => \LATCH_CLK_c\
        );

    \I__663\ : CascadeMux
    port map (
            O => \N__5129\,
            I => \U712_CHIP_RAM.N_144_cascade_\
        );

    \I__662\ : InMux
    port map (
            O => \N__5126\,
            I => \N__5123\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__5123\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_4\
        );

    \I__660\ : InMux
    port map (
            O => \N__5120\,
            I => \N__5115\
        );

    \I__659\ : InMux
    port map (
            O => \N__5119\,
            I => \N__5112\
        );

    \I__658\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5109\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__5115\,
            I => \U712_REG_SM.N_163\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__5112\,
            I => \U712_REG_SM.N_163\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__5109\,
            I => \U712_REG_SM.N_163\
        );

    \I__654\ : IoInMux
    port map (
            O => \N__5102\,
            I => \N__5098\
        );

    \I__653\ : IoInMux
    port map (
            O => \N__5101\,
            I => \N__5095\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__5098\,
            I => \N__5092\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__5095\,
            I => \N__5089\
        );

    \I__650\ : IoSpan4Mux
    port map (
            O => \N__5092\,
            I => \N__5085\
        );

    \I__649\ : Span4Mux_s2_v
    port map (
            O => \N__5089\,
            I => \N__5082\
        );

    \I__648\ : IoInMux
    port map (
            O => \N__5088\,
            I => \N__5079\
        );

    \I__647\ : Sp12to4
    port map (
            O => \N__5085\,
            I => \N__5076\
        );

    \I__646\ : Span4Mux_h
    port map (
            O => \N__5082\,
            I => \N__5073\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__5079\,
            I => \N__5070\
        );

    \I__644\ : Span12Mux_s7_h
    port map (
            O => \N__5076\,
            I => \N__5065\
        );

    \I__643\ : Sp12to4
    port map (
            O => \N__5073\,
            I => \N__5065\
        );

    \I__642\ : Span4Mux_s2_h
    port map (
            O => \N__5070\,
            I => \N__5062\
        );

    \I__641\ : Span12Mux_v
    port map (
            O => \N__5065\,
            I => \N__5059\
        );

    \I__640\ : Sp12to4
    port map (
            O => \N__5062\,
            I => \N__5056\
        );

    \I__639\ : Span12Mux_h
    port map (
            O => \N__5059\,
            I => \N__5053\
        );

    \I__638\ : Span12Mux_v
    port map (
            O => \N__5056\,
            I => \N__5050\
        );

    \I__637\ : Odrv12
    port map (
            O => \N__5053\,
            I => \CLK40_PLL_i_i\
        );

    \I__636\ : Odrv12
    port map (
            O => \N__5050\,
            I => \CLK40_PLL_i_i\
        );

    \I__635\ : CascadeMux
    port map (
            O => \N__5045\,
            I => \U712_CYCLE_TERM.N_51_cascade_\
        );

    \I__634\ : InMux
    port map (
            O => \N__5042\,
            I => \N__5039\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__5039\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\
        );

    \I__632\ : SRMux
    port map (
            O => \N__5036\,
            I => \N__5033\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__5033\,
            I => \N__5029\
        );

    \I__630\ : SRMux
    port map (
            O => \N__5032\,
            I => \N__5026\
        );

    \I__629\ : Span4Mux_h
    port map (
            O => \N__5029\,
            I => \N__5023\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__5026\,
            I => \N__5020\
        );

    \I__627\ : Odrv4
    port map (
            O => \N__5023\,
            I => \U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1\
        );

    \I__626\ : Odrv12
    port map (
            O => \N__5020\,
            I => \U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1\
        );

    \I__625\ : InMux
    port map (
            O => \N__5015\,
            I => \U712_CHIP_RAM.un2_DBR_COUNT_cry_5\
        );

    \I__624\ : InMux
    port map (
            O => \N__5012\,
            I => \U712_CHIP_RAM.un2_DBR_COUNT_cry_6\
        );

    \I__623\ : CascadeMux
    port map (
            O => \N__5009\,
            I => \N__5004\
        );

    \I__622\ : InMux
    port map (
            O => \N__5008\,
            I => \N__5001\
        );

    \I__621\ : InMux
    port map (
            O => \N__5007\,
            I => \N__4996\
        );

    \I__620\ : InMux
    port map (
            O => \N__5004\,
            I => \N__4996\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__5001\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_0\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__4996\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_0\
        );

    \I__617\ : InMux
    port map (
            O => \N__4991\,
            I => \N__4985\
        );

    \I__616\ : InMux
    port map (
            O => \N__4990\,
            I => \N__4985\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__4985\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_1\
        );

    \I__614\ : InMux
    port map (
            O => \N__4982\,
            I => \N__4979\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__4979\,
            I => \U712_REG_SM.N_159\
        );

    \I__612\ : InMux
    port map (
            O => \N__4976\,
            I => \N__4972\
        );

    \I__611\ : InMux
    port map (
            O => \N__4975\,
            I => \N__4969\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__4972\,
            I => \N__4966\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__4969\,
            I => \N__4962\
        );

    \I__608\ : Span4Mux_v
    port map (
            O => \N__4966\,
            I => \N__4959\
        );

    \I__607\ : InMux
    port map (
            O => \N__4965\,
            I => \N__4956\
        );

    \I__606\ : Span4Mux_h
    port map (
            O => \N__4962\,
            I => \N__4953\
        );

    \I__605\ : Odrv4
    port map (
            O => \N__4959\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__4956\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__603\ : Odrv4
    port map (
            O => \N__4953\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__602\ : InMux
    port map (
            O => \N__4946\,
            I => \N__4939\
        );

    \I__601\ : InMux
    port map (
            O => \N__4945\,
            I => \N__4939\
        );

    \I__600\ : InMux
    port map (
            O => \N__4944\,
            I => \N__4936\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__4939\,
            I => \U712_REG_SM.N_109\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__4936\,
            I => \U712_REG_SM.N_109\
        );

    \I__597\ : CascadeMux
    port map (
            O => \N__4931\,
            I => \N__4928\
        );

    \I__596\ : InMux
    port map (
            O => \N__4928\,
            I => \N__4925\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__4925\,
            I => \U712_REG_SM.N_164\
        );

    \I__594\ : InMux
    port map (
            O => \N__4922\,
            I => \N__4919\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__4919\,
            I => \U712_REG_SM.N_80\
        );

    \I__592\ : InMux
    port map (
            O => \N__4916\,
            I => \N__4908\
        );

    \I__591\ : CascadeMux
    port map (
            O => \N__4915\,
            I => \N__4904\
        );

    \I__590\ : CascadeMux
    port map (
            O => \N__4914\,
            I => \N__4899\
        );

    \I__589\ : CascadeMux
    port map (
            O => \N__4913\,
            I => \N__4895\
        );

    \I__588\ : InMux
    port map (
            O => \N__4912\,
            I => \N__4890\
        );

    \I__587\ : InMux
    port map (
            O => \N__4911\,
            I => \N__4890\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__4908\,
            I => \N__4887\
        );

    \I__585\ : CascadeMux
    port map (
            O => \N__4907\,
            I => \N__4882\
        );

    \I__584\ : InMux
    port map (
            O => \N__4904\,
            I => \N__4879\
        );

    \I__583\ : InMux
    port map (
            O => \N__4903\,
            I => \N__4872\
        );

    \I__582\ : InMux
    port map (
            O => \N__4902\,
            I => \N__4872\
        );

    \I__581\ : InMux
    port map (
            O => \N__4899\,
            I => \N__4872\
        );

    \I__580\ : InMux
    port map (
            O => \N__4898\,
            I => \N__4869\
        );

    \I__579\ : InMux
    port map (
            O => \N__4895\,
            I => \N__4866\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__4890\,
            I => \N__4863\
        );

    \I__577\ : Span4Mux_h
    port map (
            O => \N__4887\,
            I => \N__4860\
        );

    \I__576\ : InMux
    port map (
            O => \N__4886\,
            I => \N__4855\
        );

    \I__575\ : InMux
    port map (
            O => \N__4885\,
            I => \N__4855\
        );

    \I__574\ : InMux
    port map (
            O => \N__4882\,
            I => \N__4852\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__4879\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__4872\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__4869\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__4866\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__569\ : Odrv4
    port map (
            O => \N__4863\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__568\ : Odrv4
    port map (
            O => \N__4860\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__4855\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__4852\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__565\ : CascadeMux
    port map (
            O => \N__4835\,
            I => \N__4832\
        );

    \I__564\ : InMux
    port map (
            O => \N__4832\,
            I => \N__4829\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__4829\,
            I => \U712_REG_SM.N_96\
        );

    \I__562\ : CascadeMux
    port map (
            O => \N__4826\,
            I => \N__4821\
        );

    \I__561\ : InMux
    port map (
            O => \N__4825\,
            I => \N__4815\
        );

    \I__560\ : InMux
    port map (
            O => \N__4824\,
            I => \N__4812\
        );

    \I__559\ : InMux
    port map (
            O => \N__4821\,
            I => \N__4809\
        );

    \I__558\ : InMux
    port map (
            O => \N__4820\,
            I => \N__4802\
        );

    \I__557\ : InMux
    port map (
            O => \N__4819\,
            I => \N__4802\
        );

    \I__556\ : InMux
    port map (
            O => \N__4818\,
            I => \N__4802\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__4815\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__4812\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__4809\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__4802\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__551\ : CascadeMux
    port map (
            O => \N__4793\,
            I => \U712_REG_SM.N_96_cascade_\
        );

    \I__550\ : CascadeMux
    port map (
            O => \N__4790\,
            I => \N__4786\
        );

    \I__549\ : InMux
    port map (
            O => \N__4789\,
            I => \N__4780\
        );

    \I__548\ : InMux
    port map (
            O => \N__4786\,
            I => \N__4777\
        );

    \I__547\ : InMux
    port map (
            O => \N__4785\,
            I => \N__4772\
        );

    \I__546\ : InMux
    port map (
            O => \N__4784\,
            I => \N__4772\
        );

    \I__545\ : InMux
    port map (
            O => \N__4783\,
            I => \N__4769\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__4780\,
            I => \N__4766\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4777\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__4772\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__4769\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__540\ : Odrv4
    port map (
            O => \N__4766\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__539\ : IoInMux
    port map (
            O => \N__4757\,
            I => \N__4754\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__4754\,
            I => \N__4751\
        );

    \I__537\ : IoSpan4Mux
    port map (
            O => \N__4751\,
            I => \N__4748\
        );

    \I__536\ : Sp12to4
    port map (
            O => \N__4748\,
            I => \N__4745\
        );

    \I__535\ : Span12Mux_v
    port map (
            O => \N__4745\,
            I => \N__4741\
        );

    \I__534\ : CascadeMux
    port map (
            O => \N__4744\,
            I => \N__4738\
        );

    \I__533\ : Span12Mux_h
    port map (
            O => \N__4741\,
            I => \N__4735\
        );

    \I__532\ : InMux
    port map (
            O => \N__4738\,
            I => \N__4732\
        );

    \I__531\ : Odrv12
    port map (
            O => \N__4735\,
            I => \UDSn_c\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__4732\,
            I => \UDSn_c\
        );

    \I__529\ : InMux
    port map (
            O => \N__4727\,
            I => \N__4724\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__4724\,
            I => \U712_BYTE_ENABLE_UDS_0\
        );

    \I__527\ : InMux
    port map (
            O => \N__4721\,
            I => \N__4718\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__4718\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__525\ : InMux
    port map (
            O => \N__4715\,
            I => \N__4712\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__4712\,
            I => \U712_REG_SM.N_166\
        );

    \I__523\ : IoInMux
    port map (
            O => \N__4709\,
            I => \N__4706\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__4706\,
            I => \N__4703\
        );

    \I__521\ : Span4Mux_s3_v
    port map (
            O => \N__4703\,
            I => \N__4700\
        );

    \I__520\ : Span4Mux_h
    port map (
            O => \N__4700\,
            I => \N__4697\
        );

    \I__519\ : Span4Mux_h
    port map (
            O => \N__4697\,
            I => \N__4694\
        );

    \I__518\ : Sp12to4
    port map (
            O => \N__4694\,
            I => \N__4691\
        );

    \I__517\ : Span12Mux_s10_v
    port map (
            O => \N__4691\,
            I => \N__4687\
        );

    \I__516\ : InMux
    port map (
            O => \N__4690\,
            I => \N__4684\
        );

    \I__515\ : Odrv12
    port map (
            O => \N__4687\,
            I => \LDSn_c\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__4684\,
            I => \LDSn_c\
        );

    \I__513\ : IoInMux
    port map (
            O => \N__4679\,
            I => \N__4676\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__4676\,
            I => \N__4673\
        );

    \I__511\ : Span4Mux_s2_v
    port map (
            O => \N__4673\,
            I => \N__4670\
        );

    \I__510\ : Span4Mux_v
    port map (
            O => \N__4670\,
            I => \N__4667\
        );

    \I__509\ : Span4Mux_v
    port map (
            O => \N__4667\,
            I => \N__4664\
        );

    \I__508\ : Span4Mux_v
    port map (
            O => \N__4664\,
            I => \N__4660\
        );

    \I__507\ : InMux
    port map (
            O => \N__4663\,
            I => \N__4657\
        );

    \I__506\ : Odrv4
    port map (
            O => \N__4660\,
            I => \DBDIR_c\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4657\,
            I => \DBDIR_c\
        );

    \I__504\ : InMux
    port map (
            O => \N__4652\,
            I => \N__4649\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4649\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_2\
        );

    \I__502\ : InMux
    port map (
            O => \N__4646\,
            I => \U712_CHIP_RAM.un2_DBR_COUNT_cry_1\
        );

    \I__501\ : InMux
    port map (
            O => \N__4643\,
            I => \N__4640\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4640\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_3\
        );

    \I__499\ : InMux
    port map (
            O => \N__4637\,
            I => \U712_CHIP_RAM.un2_DBR_COUNT_cry_2\
        );

    \I__498\ : InMux
    port map (
            O => \N__4634\,
            I => \N__4631\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__4631\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_4\
        );

    \I__496\ : InMux
    port map (
            O => \N__4628\,
            I => \U712_CHIP_RAM.un2_DBR_COUNT_cry_3\
        );

    \I__495\ : InMux
    port map (
            O => \N__4625\,
            I => \U712_CHIP_RAM.un2_DBR_COUNT_cry_4\
        );

    \I__494\ : CascadeMux
    port map (
            O => \N__4622\,
            I => \U712_REG_SM.N_109_cascade_\
        );

    \I__493\ : CascadeMux
    port map (
            O => \N__4619\,
            I => \U712_REG_SM.STATE_COUNTc_0_0_cascade_\
        );

    \I__492\ : InMux
    port map (
            O => \N__4616\,
            I => \N__4604\
        );

    \I__491\ : InMux
    port map (
            O => \N__4615\,
            I => \N__4604\
        );

    \I__490\ : InMux
    port map (
            O => \N__4614\,
            I => \N__4604\
        );

    \I__489\ : InMux
    port map (
            O => \N__4613\,
            I => \N__4604\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__4604\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__487\ : CascadeMux
    port map (
            O => \N__4601\,
            I => \U712_REG_SM.REG_CYCLE_0_sqmuxa_cascade_\
        );

    \I__486\ : InMux
    port map (
            O => \N__4598\,
            I => \N__4594\
        );

    \I__485\ : InMux
    port map (
            O => \N__4597\,
            I => \N__4591\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4594\,
            I => \U712_REG_SM.N_185\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__4591\,
            I => \U712_REG_SM.N_185\
        );

    \I__482\ : InMux
    port map (
            O => \N__4586\,
            I => \N__4582\
        );

    \I__481\ : InMux
    port map (
            O => \N__4585\,
            I => \N__4576\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__4582\,
            I => \N__4573\
        );

    \I__479\ : InMux
    port map (
            O => \N__4581\,
            I => \N__4570\
        );

    \I__478\ : InMux
    port map (
            O => \N__4580\,
            I => \N__4565\
        );

    \I__477\ : InMux
    port map (
            O => \N__4579\,
            I => \N__4565\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__4576\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__475\ : Odrv4
    port map (
            O => \N__4573\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4570\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__4565\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__472\ : CascadeMux
    port map (
            O => \N__4556\,
            I => \N__4553\
        );

    \I__471\ : InMux
    port map (
            O => \N__4553\,
            I => \N__4550\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4550\,
            I => \U712_REG_SM.N_109_0\
        );

    \I__469\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4543\
        );

    \I__468\ : InMux
    port map (
            O => \N__4546\,
            I => \N__4540\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__4543\,
            I => \U712_REG_SM.N_105_0\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__4540\,
            I => \U712_REG_SM.N_105_0\
        );

    \I__465\ : InMux
    port map (
            O => \N__4535\,
            I => \N__4531\
        );

    \I__464\ : InMux
    port map (
            O => \N__4534\,
            I => \N__4525\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__4531\,
            I => \N__4522\
        );

    \I__462\ : InMux
    port map (
            O => \N__4530\,
            I => \N__4519\
        );

    \I__461\ : InMux
    port map (
            O => \N__4529\,
            I => \N__4516\
        );

    \I__460\ : InMux
    port map (
            O => \N__4528\,
            I => \N__4513\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__4525\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__458\ : Odrv4
    port map (
            O => \N__4522\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__4519\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__4516\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__4513\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__454\ : InMux
    port map (
            O => \N__4502\,
            I => \N__4499\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__4499\,
            I => \N__4495\
        );

    \I__452\ : IoInMux
    port map (
            O => \N__4498\,
            I => \N__4492\
        );

    \I__451\ : Span4Mux_h
    port map (
            O => \N__4495\,
            I => \N__4489\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4492\,
            I => \N__4486\
        );

    \I__449\ : Span4Mux_v
    port map (
            O => \N__4489\,
            I => \N__4483\
        );

    \I__448\ : IoSpan4Mux
    port map (
            O => \N__4486\,
            I => \N__4480\
        );

    \I__447\ : Span4Mux_v
    port map (
            O => \N__4483\,
            I => \N__4477\
        );

    \I__446\ : IoSpan4Mux
    port map (
            O => \N__4480\,
            I => \N__4474\
        );

    \I__445\ : IoSpan4Mux
    port map (
            O => \N__4477\,
            I => \N__4469\
        );

    \I__444\ : IoSpan4Mux
    port map (
            O => \N__4474\,
            I => \N__4469\
        );

    \I__443\ : Odrv4
    port map (
            O => \N__4469\,
            I => \C1_c\
        );

    \I__442\ : InMux
    port map (
            O => \N__4466\,
            I => \N__4462\
        );

    \I__441\ : InMux
    port map (
            O => \N__4465\,
            I => \N__4459\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__4462\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__4459\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__438\ : InMux
    port map (
            O => \N__4454\,
            I => \N__4450\
        );

    \I__437\ : InMux
    port map (
            O => \N__4453\,
            I => \N__4447\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__4450\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__4447\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__434\ : CascadeMux
    port map (
            O => \N__4442\,
            I => \U712_REG_SM.N_157_cascade_\
        );

    \I__433\ : InMux
    port map (
            O => \N__4439\,
            I => \N__4436\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__4436\,
            I => \N__4432\
        );

    \I__431\ : InMux
    port map (
            O => \N__4435\,
            I => \N__4429\
        );

    \I__430\ : Span4Mux_h
    port map (
            O => \N__4432\,
            I => \N__4424\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__4429\,
            I => \N__4424\
        );

    \I__428\ : Span4Mux_v
    port map (
            O => \N__4424\,
            I => \N__4421\
        );

    \I__427\ : Span4Mux_h
    port map (
            O => \N__4421\,
            I => \N__4418\
        );

    \I__426\ : Sp12to4
    port map (
            O => \N__4418\,
            I => \N__4415\
        );

    \I__425\ : Odrv12
    port map (
            O => \N__4415\,
            I => \DBRn_c\
        );

    \I__424\ : IoInMux
    port map (
            O => \N__4412\,
            I => \N__4409\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__4409\,
            I => \N__4406\
        );

    \I__422\ : IoSpan4Mux
    port map (
            O => \N__4406\,
            I => \N__4403\
        );

    \I__421\ : Span4Mux_s3_v
    port map (
            O => \N__4403\,
            I => \N__4400\
        );

    \I__420\ : Sp12to4
    port map (
            O => \N__4400\,
            I => \N__4397\
        );

    \I__419\ : Span12Mux_s11_v
    port map (
            O => \N__4397\,
            I => \N__4393\
        );

    \I__418\ : InMux
    port map (
            O => \N__4396\,
            I => \N__4390\
        );

    \I__417\ : Odrv12
    port map (
            O => \N__4393\,
            I => \REGENn_c\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__4390\,
            I => \REGENn_c\
        );

    \I__415\ : InMux
    port map (
            O => \N__4385\,
            I => \N__4381\
        );

    \I__414\ : InMux
    port map (
            O => \N__4384\,
            I => \N__4378\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__4381\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__4378\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__411\ : CascadeMux
    port map (
            O => \N__4373\,
            I => \U712_REG_SM.un6_REG_CYCLE_START_cascade_\
        );

    \I__410\ : InMux
    port map (
            O => \N__4370\,
            I => \N__4367\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__4367\,
            I => \N__4364\
        );

    \I__408\ : Span12Mux_h
    port map (
            O => \N__4364\,
            I => \N__4361\
        );

    \I__407\ : Span12Mux_v
    port map (
            O => \N__4361\,
            I => \N__4358\
        );

    \I__406\ : Odrv12
    port map (
            O => \N__4358\,
            I => \REGSPACEn_c\
        );

    \I__405\ : IoInMux
    port map (
            O => \N__4355\,
            I => \N__4352\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__4352\,
            I => \N__4349\
        );

    \I__403\ : IoSpan4Mux
    port map (
            O => \N__4349\,
            I => \N__4346\
        );

    \I__402\ : IoSpan4Mux
    port map (
            O => \N__4346\,
            I => \N__4343\
        );

    \I__401\ : Span4Mux_s3_h
    port map (
            O => \N__4343\,
            I => \N__4339\
        );

    \I__400\ : InMux
    port map (
            O => \N__4342\,
            I => \N__4336\
        );

    \I__399\ : Span4Mux_h
    port map (
            O => \N__4339\,
            I => \N__4333\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__4336\,
            I => \N__4330\
        );

    \I__397\ : Sp12to4
    port map (
            O => \N__4333\,
            I => \N__4327\
        );

    \I__396\ : Span4Mux_v
    port map (
            O => \N__4330\,
            I => \N__4324\
        );

    \I__395\ : Span12Mux_h
    port map (
            O => \N__4327\,
            I => \N__4319\
        );

    \I__394\ : Sp12to4
    port map (
            O => \N__4324\,
            I => \N__4319\
        );

    \I__393\ : Span12Mux_h
    port map (
            O => \N__4319\,
            I => \N__4316\
        );

    \I__392\ : Odrv12
    port map (
            O => \N__4316\,
            I => \C3_c\
        );

    \I__391\ : InMux
    port map (
            O => \N__4313\,
            I => \N__4310\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__4310\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__389\ : InMux
    port map (
            O => \N__4307\,
            I => \N__4304\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__4304\,
            I => \U712_REG_SM.STATE_COUNT_1_sqmuxa_1\
        );

    \I__387\ : InMux
    port map (
            O => \N__4301\,
            I => \N__4298\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__4298\,
            I => \U712_REG_SM.N_188\
        );

    \I__385\ : IoInMux
    port map (
            O => \N__4295\,
            I => \N__4292\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__4292\,
            I => \N__4289\
        );

    \I__383\ : Span4Mux_s1_h
    port map (
            O => \N__4289\,
            I => \N__4286\
        );

    \I__382\ : Span4Mux_h
    port map (
            O => \N__4286\,
            I => \N__4283\
        );

    \I__381\ : Odrv4
    port map (
            O => \N__4283\,
            I => \DBRn_c_i_0\
        );

    \I__380\ : IoInMux
    port map (
            O => \N__4280\,
            I => \N__4277\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__4277\,
            I => \N__4274\
        );

    \I__378\ : Span4Mux_s3_v
    port map (
            O => \N__4274\,
            I => \N__4271\
        );

    \I__377\ : Span4Mux_h
    port map (
            O => \N__4271\,
            I => \N__4268\
        );

    \I__376\ : Odrv4
    port map (
            O => \N__4268\,
            I => \CLK80_PLL_i_i\
        );

    \I__375\ : InMux
    port map (
            O => \N__4265\,
            I => \N__4262\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__4262\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__373\ : IoInMux
    port map (
            O => \N__4259\,
            I => \N__4256\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__4256\,
            I => \N__4253\
        );

    \I__371\ : IoSpan4Mux
    port map (
            O => \N__4253\,
            I => \N__4250\
        );

    \I__370\ : Span4Mux_s2_v
    port map (
            O => \N__4250\,
            I => \N__4247\
        );

    \I__369\ : Sp12to4
    port map (
            O => \N__4247\,
            I => \N__4244\
        );

    \I__368\ : Span12Mux_v
    port map (
            O => \N__4244\,
            I => \N__4241\
        );

    \I__367\ : Odrv12
    port map (
            O => \N__4241\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            I => \N__5628\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            I => \N__5630\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__5624\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__5625\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            I => \N__5623\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            I => \N__5627\
        );

    \INVU712_CHIP_RAM.DMA_A20C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A20C_net\,
            I => \N__5622\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__5626\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_10_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_9_0_\
        );

    \IN_MUX_bfv_10_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_13_0_\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4498\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7688\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4295\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4355\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9541\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10982\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_3_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10343\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_0_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4439\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10337\,
            ce => 'H',
            sr => \N__10953\
        );

    \DBR_SYNC_1_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4265\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10337\,
            ce => 'H',
            sr => \N__10953\
        );

    \DBRn_ibuf_RNIBAB_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4435\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101110101010"
        )
    port map (
            in0 => \N__4307\,
            in1 => \N__4301\,
            in2 => \N__4915\,
            in3 => \N__4396\,
            lcout => \REGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10339\,
            ce => 'H',
            sr => \N__10945\
        );

    \U712_REG_SM.START_RST_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__4385\,
            in1 => \N__4454\,
            in2 => \_gnd_net_\,
            in3 => \N__4535\,
            lcout => \U712_REG_SM.START_RSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10330\,
            ce => 'H',
            sr => \N__10949\
        );

    \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4384\,
            in2 => \_gnd_net_\,
            in3 => \N__4585\,
            lcout => OPEN,
            ltout => \U712_REG_SM.un6_REG_CYCLE_START_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011000100"
        )
    port map (
            in0 => \N__5405\,
            in1 => \N__7879\,
            in2 => \N__4373\,
            in3 => \N__4370\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_0_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4342\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10336\,
            ce => 'H',
            sr => \N__10938\
        );

    \U712_REG_SM.C3_SYNC_1_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4313\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10336\,
            ce => 'H',
            sr => \N__10938\
        );

    \U712_REG_SM.REGENn_RNO_1_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4586\,
            in1 => \N__5513\,
            in2 => \N__4913\,
            in3 => \N__4976\,
            lcout => \U712_REG_SM.STATE_COUNT_1_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_RNO_0_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4530\,
            in2 => \_gnd_net_\,
            in3 => \N__5512\,
            lcout => \U712_REG_SM.N_188\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_RNO_0_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6774\,
            in1 => \N__6848\,
            in2 => \N__7002\,
            in3 => \N__10805\,
            lcout => \U712_REG_SM.N_166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.WRITE_CYCLE_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__10813\,
            in1 => \N__4466\,
            in2 => \_gnd_net_\,
            in3 => \N__4453\,
            lcout => \U712_REG_SM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10326\,
            ce => 'H',
            sr => \N__10950\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__5526\,
            in1 => \N__4912\,
            in2 => \_gnd_net_\,
            in3 => \N__4818\,
            lcout => \U712_REG_SM.N_164\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__4465\,
            in1 => \N__4820\,
            in2 => \_gnd_net_\,
            in3 => \N__4597\,
            lcout => \U712_REG_SM.N_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4579\,
            in1 => \N__4911\,
            in2 => \N__5534\,
            in3 => \N__4965\,
            lcout => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4819\,
            in1 => \N__4944\,
            in2 => \N__4790\,
            in3 => \N__4580\,
            lcout => \U712_REG_SM.N_159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__4614\,
            in1 => \N__4886\,
            in2 => \N__4826\,
            in3 => \N__6196\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_157_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001010"
        )
    port map (
            in0 => \N__7878\,
            in1 => \N__5530\,
            in2 => \N__4442\,
            in3 => \N__4903\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__4783\,
            in1 => \N__4885\,
            in2 => \_gnd_net_\,
            in3 => \N__5521\,
            lcout => \U712_REG_SM.N_185\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4528\,
            in2 => \_gnd_net_\,
            in3 => \N__4613\,
            lcout => \U712_REG_SM.N_109\,
            ltout => \U712_REG_SM.N_109_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4902\,
            in1 => \N__5523\,
            in2 => \N__4622\,
            in3 => \N__6198\,
            lcout => OPEN,
            ltout => \U712_REG_SM.STATE_COUNTc_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__7877\,
            in1 => \N__4547\,
            in2 => \N__4619\,
            in3 => \N__4616\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_0_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4615\,
            in1 => \N__5522\,
            in2 => \N__4914\,
            in3 => \N__6197\,
            lcout => OPEN,
            ltout => \U712_REG_SM.REG_CYCLE_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011101100"
        )
    port map (
            in0 => \N__7876\,
            in1 => \N__11634\,
            in2 => \N__4601\,
            in3 => \N__4598\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__7880\,
            in1 => \N__4546\,
            in2 => \N__4556\,
            in3 => \N__4534\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__5524\,
            in1 => \N__4975\,
            in2 => \_gnd_net_\,
            in3 => \N__4581\,
            lcout => \U712_REG_SM.N_109_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4898\,
            in2 => \_gnd_net_\,
            in3 => \N__5525\,
            lcout => \U712_REG_SM.N_105_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIVCF31_1_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__4789\,
            in1 => \N__4529\,
            in2 => \N__4907\,
            in3 => \N__5488\,
            lcout => \U712_REG_SM.N_163\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_0_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4502\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10338\,
            ce => 'H',
            sr => \N__10922\
        );

    \U712_REG_SM.C1_SYNC_1_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4721\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10338\,
            ce => 'H',
            sr => \N__10922\
        );

    \U712_REG_SM.LDSn_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__4690\,
            in1 => \N__5120\,
            in2 => \N__5533\,
            in3 => \N__4715\,
            lcout => \LDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10338\,
            ce => 'H',
            sr => \N__10922\
        );

    \U712_CHIP_RAM.DBDIR_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__6239\,
            in1 => \N__4663\,
            in2 => \_gnd_net_\,
            in3 => \N__5042\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10312\,
            ce => 'H',
            sr => \N__10954\
        );

    \U712_CHIP_RAM.DBR_COUNT_0_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5008\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10317\,
            ce => 'H',
            sr => \N__5032\
        );

    \U712_CHIP_RAM.un2_DBR_COUNT_cry_1_c_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4990\,
            in2 => \N__5009\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \U712_CHIP_RAM.un2_DBR_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBR_COUNT_2_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4652\,
            in2 => \_gnd_net_\,
            in3 => \N__4646\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un2_DBR_COUNT_cry_1\,
            carryout => \U712_CHIP_RAM.un2_DBR_COUNT_cry_2\,
            clk => \N__10323\,
            ce => 'H',
            sr => \N__5036\
        );

    \U712_CHIP_RAM.DBR_COUNT_3_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4643\,
            in2 => \_gnd_net_\,
            in3 => \N__4637\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un2_DBR_COUNT_cry_2\,
            carryout => \U712_CHIP_RAM.un2_DBR_COUNT_cry_3\,
            clk => \N__10323\,
            ce => 'H',
            sr => \N__5036\
        );

    \U712_CHIP_RAM.DBR_COUNT_4_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4634\,
            in2 => \_gnd_net_\,
            in3 => \N__4628\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un2_DBR_COUNT_cry_3\,
            carryout => \U712_CHIP_RAM.un2_DBR_COUNT_cry_4\,
            clk => \N__10323\,
            ce => 'H',
            sr => \N__5036\
        );

    \U712_CHIP_RAM.DBR_COUNT_5_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5195\,
            in2 => \_gnd_net_\,
            in3 => \N__4625\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un2_DBR_COUNT_cry_4\,
            carryout => \U712_CHIP_RAM.un2_DBR_COUNT_cry_5\,
            clk => \N__10323\,
            ce => 'H',
            sr => \N__5036\
        );

    \U712_CHIP_RAM.DBR_COUNT_6_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5183\,
            in2 => \_gnd_net_\,
            in3 => \N__5015\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un2_DBR_COUNT_cry_5\,
            carryout => \U712_CHIP_RAM.un2_DBR_COUNT_cry_6\,
            clk => \N__10323\,
            ce => 'H',
            sr => \N__5036\
        );

    \U712_CHIP_RAM.DBR_COUNT_7_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5171\,
            in2 => \_gnd_net_\,
            in3 => \N__5012\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10323\,
            ce => 'H',
            sr => \N__5036\
        );

    \U712_CHIP_RAM.DBR_COUNT_1_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__4991\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5007\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10323\,
            ce => 'H',
            sr => \N__5036\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__4946\,
            in1 => \N__4825\,
            in2 => \N__4835\,
            in3 => \N__4982\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10327\,
            ce => 'H',
            sr => \N__10939\
        );

    \U712_REG_SM.REG_TACK_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__6273\,
            in1 => \N__4945\,
            in2 => \N__4931\,
            in3 => \N__4922\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10327\,
            ce => 'H',
            sr => \N__10939\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__4784\,
            in1 => \N__4916\,
            in2 => \_gnd_net_\,
            in3 => \N__5531\,
            lcout => \U712_REG_SM.N_96\,
            ltout => \U712_REG_SM.N_96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__7853\,
            in1 => \N__4824\,
            in2 => \N__4793\,
            in3 => \N__4785\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDSn_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__4727\,
            in1 => \N__5119\,
            in2 => \N__4744\,
            in3 => \N__5517\,
            lcout => \UDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10334\,
            ce => 'H',
            sr => \N__10923\
        );

    \U712_BYTE_ENABLE.UDS_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__6862\,
            in1 => \N__6971\,
            in2 => \N__6818\,
            in3 => \N__10806\,
            lcout => \U712_BYTE_ENABLE_UDS_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_RNO_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10980\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5118\,
            lcout => \U712_REG_SM.N_163_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_RNI8MQ3_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5901\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__6036\,
            in1 => \N__6283\,
            in2 => \_gnd_net_\,
            in3 => \N__7090\,
            lcout => \U712_CYCLE_TERM.N_47_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110111"
        )
    port map (
            in0 => \N__7091\,
            in1 => \N__6037\,
            in2 => \N__6287\,
            in3 => \N__6072\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_51_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__6038\,
            in1 => \N__7850\,
            in2 => \N__5045\,
            in3 => \N__5888\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI1KG35_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8011\,
            in1 => \N__7269\,
            in2 => \_gnd_net_\,
            in3 => \N__7394\,
            lcout => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__5729\,
            in1 => \N__5546\,
            in2 => \_gnd_net_\,
            in3 => \N__7849\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__6205\,
            in1 => \N__7848\,
            in2 => \_gnd_net_\,
            in3 => \N__6151\,
            lcout => \U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__7792\,
            in1 => \N__7977\,
            in2 => \_gnd_net_\,
            in3 => \N__5804\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_RNIGHLF1_0_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111011111111"
        )
    port map (
            in0 => \N__5727\,
            in1 => \N__5670\,
            in2 => \N__6157\,
            in3 => \N__7197\,
            lcout => \U712_CHIP_RAM.N_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7791\,
            in2 => \_gnd_net_\,
            in3 => \N__5671\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNO_0_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001000"
        )
    port map (
            in0 => \N__5194\,
            in1 => \N__5182\,
            in2 => \N__7307\,
            in3 => \N__5170\,
            lcout => \U712_CHIP_RAM.N_152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIF9JU1_2_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5740\,
            in2 => \_gnd_net_\,
            in3 => \N__8219\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_1_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5540\,
            in1 => \N__5993\,
            in2 => \N__8035\,
            in3 => \N__5126\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__7851\,
            in1 => \N__5140\,
            in2 => \N__5159\,
            in3 => \N__5783\,
            lcout => \LATCH_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_2_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__8319\,
            in1 => \N__8112\,
            in2 => \_gnd_net_\,
            in3 => \N__8213\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_144_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111101"
        )
    port map (
            in0 => \N__7852\,
            in1 => \N__8224\,
            in2 => \N__5129\,
            in3 => \N__7547\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_29_i_a2_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_3_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6391\,
            in1 => \N__6373\,
            in2 => \N__6356\,
            in3 => \N__6331\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_2_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__8320\,
            in1 => \N__8113\,
            in2 => \_gnd_net_\,
            in3 => \N__8214\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_1_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8212\,
            in1 => \N__7546\,
            in2 => \N__8121\,
            in3 => \N__8318\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER16_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5532\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10335\,
            ce => \N__5417\,
            sr => \N__10913\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5401\,
            in2 => \_gnd_net_\,
            in3 => \N__5375\,
            lcout => \U712_CHIP_RAM.un3_CPU_CYCLE_START\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_10_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__9337\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11653\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__6085\,
            in1 => \N__5273\,
            in2 => \_gnd_net_\,
            in3 => \N__5330\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10304\,
            ce => 'H',
            sr => \N__10951\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110110011101110"
        )
    port map (
            in0 => \N__5213\,
            in1 => \N__6119\,
            in2 => \N__5903\,
            in3 => \N__6065\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10304\,
            ce => 'H',
            sr => \N__10951\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5558\,
            in2 => \_gnd_net_\,
            in3 => \N__5198\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_10_9_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__5629\,
            ce => 'H',
            sr => \N__6023\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5585\,
            in2 => \_gnd_net_\,
            in3 => \N__5651\,
            lcout => \U712_CHIP_RAM.REFRESH5lto1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__5629\,
            ce => 'H',
            sr => \N__6023\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5597\,
            in2 => \_gnd_net_\,
            in3 => \N__5648\,
            lcout => \U712_CHIP_RAM.REFRESH5lto2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__5629\,
            ce => 'H',
            sr => \N__6023\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5704\,
            in2 => \_gnd_net_\,
            in3 => \N__5645\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__5629\,
            ce => 'H',
            sr => \N__6023\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5572\,
            in2 => \_gnd_net_\,
            in3 => \N__5642\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__5629\,
            ce => 'H',
            sr => \N__6023\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5753\,
            in2 => \_gnd_net_\,
            in3 => \N__5639\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__5629\,
            ce => 'H',
            sr => \N__6023\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5765\,
            in2 => \_gnd_net_\,
            in3 => \N__5636\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__5629\,
            ce => 'H',
            sr => \N__6023\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5777\,
            in2 => \_gnd_net_\,
            in3 => \N__5633\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5629\,
            ce => 'H',
            sr => \N__6023\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__5596\,
            in1 => \N__5584\,
            in2 => \N__5573\,
            in3 => \N__5557\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001101"
        )
    port map (
            in0 => \N__5728\,
            in1 => \N__8686\,
            in2 => \N__5675\,
            in3 => \N__6152\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_START_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5776\,
            in1 => \N__5764\,
            in2 => \_gnd_net_\,
            in3 => \N__5752\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011111111"
        )
    port map (
            in0 => \N__7969\,
            in1 => \N__5741\,
            in2 => \_gnd_net_\,
            in3 => \N__7380\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_i_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_RNI2NL01_0_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__6153\,
            in1 => \N__5726\,
            in2 => \_gnd_net_\,
            in3 => \N__5669\,
            lcout => \U712_CHIP_RAM.N_119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010110000"
        )
    port map (
            in0 => \N__5705\,
            in1 => \N__5690\,
            in2 => \N__7820\,
            in3 => \N__5684\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIGI6A1_2_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__7785\,
            in1 => \N__7942\,
            in2 => \_gnd_net_\,
            in3 => \N__8198\,
            lcout => \U712_CHIP_RAM.N_187\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_3_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7636\,
            in1 => \N__8328\,
            in2 => \_gnd_net_\,
            in3 => \N__8448\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER18\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7943\,
            in2 => \N__5678\,
            in3 => \N__7790\,
            lcout => \U712_CHIP_RAM.N_154\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__10580\,
            in1 => \N__7784\,
            in2 => \_gnd_net_\,
            in3 => \N__10667\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__7145\,
            in1 => \N__8199\,
            in2 => \_gnd_net_\,
            in3 => \N__7618\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER33_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100110011"
        )
    port map (
            in0 => \N__7944\,
            in1 => \N__7786\,
            in2 => \N__5840\,
            in3 => \N__5789\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4HBB7_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__7968\,
            in1 => \N__7375\,
            in2 => \_gnd_net_\,
            in3 => \N__7617\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_i_0_68_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIH3D4G_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__7973\,
            in1 => \N__5803\,
            in2 => \N__5837\,
            in3 => \N__6428\,
            lcout => \U712_CHIP_RAM.N_64\,
            ltout => \U712_CHIP_RAM.N_64_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__6582\,
            in1 => \N__5978\,
            in2 => \N__5834\,
            in3 => \N__7172\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10319\,
            ce => \N__5921\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIT7PC1_1_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__8303\,
            in1 => \N__8092\,
            in2 => \_gnd_net_\,
            in3 => \N__8197\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER37_0_a3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001011011110"
        )
    port map (
            in0 => \N__5827\,
            in1 => \N__5951\,
            in2 => \N__7559\,
            in3 => \N__5810\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10319\,
            ce => \N__5921\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_1_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8087\,
            in1 => \N__7537\,
            in2 => \_gnd_net_\,
            in3 => \N__8196\,
            lcout => \U712_CHIP_RAM.N_177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011111010"
        )
    port map (
            in0 => \N__5802\,
            in1 => \N__7579\,
            in2 => \N__8010\,
            in3 => \N__7374\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7558\,
            in2 => \_gnd_net_\,
            in3 => \N__8687\,
            lcout => \U712_CHIP_RAM.LATCH_CLK_6\,
            ltout => OPEN,
            carryin => \bfn_10_13_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5952\,
            in1 => \N__8108\,
            in2 => \_gnd_net_\,
            in3 => \N__5981\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__10324\,
            ce => \N__5920\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8225\,
            in2 => \_gnd_net_\,
            in3 => \N__5969\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5953\,
            in1 => \N__8326\,
            in2 => \_gnd_net_\,
            in3 => \N__5966\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__10324\,
            ce => \N__5920\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5948\,
            in1 => \N__6354\,
            in2 => \_gnd_net_\,
            in3 => \N__5963\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__10324\,
            ce => \N__5920\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5954\,
            in1 => \N__6374\,
            in2 => \_gnd_net_\,
            in3 => \N__5960\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__10324\,
            ce => \N__5920\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5949\,
            in1 => \N__6392\,
            in2 => \_gnd_net_\,
            in3 => \N__5957\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__10324\,
            ce => \N__5920\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__6332\,
            in1 => \N__5950\,
            in2 => \_gnd_net_\,
            in3 => \N__5924\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10324\,
            ce => \N__5920\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNIHHJP6_0_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6557\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UUBE_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010010101000"
        )
    port map (
            in0 => \N__7011\,
            in1 => \N__6932\,
            in2 => \N__6894\,
            in3 => \N__6817\,
            lcout => \UUBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7845\,
            in1 => \N__5902\,
            in2 => \_gnd_net_\,
            in3 => \N__6073\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10298\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7847\,
            in2 => \_gnd_net_\,
            in3 => \N__6118\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10298\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__7846\,
            in1 => \_gnd_net_\,
            in2 => \N__6104\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10298\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6117\,
            in2 => \_gnd_net_\,
            in3 => \N__6100\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101010001010"
        )
    port map (
            in0 => \N__9299\,
            in1 => \N__7148\,
            in2 => \N__8045\,
            in3 => \N__6452\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10305\,
            ce => 'H',
            sr => \N__10940\
        );

    \U712_CHIP_RAM.DBENn_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100111011101110"
        )
    port map (
            in0 => \N__6248\,
            in1 => \N__8703\,
            in2 => \N__7397\,
            in3 => \N__9983\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10305\,
            ce => 'H',
            sr => \N__10940\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000111000001100"
        )
    port map (
            in0 => \N__6092\,
            in1 => \N__6086\,
            in2 => \N__6074\,
            in3 => \N__6254\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10305\,
            ce => 'H',
            sr => \N__10940\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9768\,
            in1 => \N__9864\,
            in2 => \N__9698\,
            in3 => \N__9485\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000111110011"
        )
    port map (
            in0 => \N__6524\,
            in1 => \N__8654\,
            in2 => \N__10598\,
            in3 => \N__9249\,
            lcout => \CLMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNITQTQ3_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__10720\,
            in1 => \N__7560\,
            in2 => \N__6311\,
            in3 => \N__8475\,
            lcout => \U712_CHIP_RAM.LATCH_CLK_0_sqmuxa\,
            ltout => \U712_CHIP_RAM.LATCH_CLK_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI17CI7_0_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__8476\,
            in1 => \N__7565\,
            in2 => \N__6290\,
            in3 => \N__6310\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER38_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__6282\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7080\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2RSLC_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011110000"
        )
    port map (
            in0 => \N__7379\,
            in1 => \N__7247\,
            in2 => \N__8044\,
            in3 => \N__7146\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_7_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6242\,
            in3 => \N__10981\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_7_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNIQJ661_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__7656\,
            in1 => \N__7196\,
            in2 => \_gnd_net_\,
            in3 => \N__7299\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERlde_0_a3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111011101"
        )
    port map (
            in0 => \N__10801\,
            in1 => \N__7248\,
            in2 => \_gnd_net_\,
            in3 => \N__6235\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_DISABLE_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__6209\,
            in1 => \N__6170\,
            in2 => \N__6161\,
            in3 => \N__7782\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_DISABLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIDTSL_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__10722\,
            in1 => \_gnd_net_\,
            in2 => \N__8125\,
            in3 => \N__9250\,
            lcout => \U712_CHIP_RAM.CLK_EN_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10721\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7554\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_108_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIE4LR1_1_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__8220\,
            in1 => \N__8009\,
            in2 => \N__6434\,
            in3 => \N__8117\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_i_0_68_i_a3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIEL6M4_3_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010101010101"
        )
    port map (
            in0 => \N__7783\,
            in1 => \N__8337\,
            in2 => \N__6431\,
            in3 => \N__8465\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_i_0_68_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8471\,
            in1 => \N__8034\,
            in2 => \N__8238\,
            in3 => \N__6398\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000110011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6409\,
            in2 => \N__6422\,
            in3 => \N__6599\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10315\,
            ce => 'H',
            sr => \N__10924\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_1_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7545\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8302\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI7MG83_1_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__8301\,
            in1 => \N__8227\,
            in2 => \N__8474\,
            in3 => \N__8090\,
            lcout => \U712_CHIP_RAM.N_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6390\,
            in1 => \N__6372\,
            in2 => \N__6355\,
            in3 => \N__6330\,
            lcout => \U712_CHIP_RAM.N_331_3\,
            ltout => \U712_CHIP_RAM.N_331_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_1_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8297\,
            in1 => \N__8088\,
            in2 => \N__6314\,
            in3 => \N__7542\,
            lcout => \U712_CHIP_RAM.N_172\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIU95J5_0_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100111111"
        )
    port map (
            in0 => \N__7544\,
            in1 => \N__8457\,
            in2 => \N__6515\,
            in3 => \N__6306\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER17_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__8200\,
            in1 => \N__7543\,
            in2 => \N__8327\,
            in3 => \N__8089\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_0_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__6461\,
            in1 => \N__7268\,
            in2 => \N__7395\,
            in3 => \N__9518\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.BANK0_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111101001110"
        )
    port map (
            in0 => \N__8552\,
            in1 => \N__6490\,
            in2 => \N__6506\,
            in3 => \N__8515\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10320\,
            ce => 'H',
            sr => \N__10917\
        );

    \U712_CHIP_RAM.BANK0_RNO_1_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11297\,
            in1 => \N__6479\,
            in2 => \_gnd_net_\,
            in3 => \N__6448\,
            lcout => \U712_CHIP_RAM.A_m_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_3_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__8459\,
            in1 => \N__8330\,
            in2 => \N__8234\,
            in3 => \N__7118\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER15\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNI0NAU5_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7283\,
            in1 => \N__7267\,
            in2 => \N__6455\,
            in3 => \N__7208\,
            lcout => \U712_CHIP_RAM.A_m_2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8091\,
            in2 => \_gnd_net_\,
            in3 => \N__7541\,
            lcout => \U712_CHIP_RAM.N_94\,
            ltout => \U712_CHIP_RAM.N_94_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_3_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8329\,
            in1 => \N__8215\,
            in2 => \N__6437\,
            in3 => \N__8458\,
            lcout => \U712_CHIP_RAM.N_173\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRU1VF_3_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__6584\,
            in1 => \N__6556\,
            in2 => \N__6536\,
            in3 => \N__6542\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_1\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIG5PHK_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6587\,
            in3 => \N__8356\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNIHHJP6_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6583\,
            in1 => \N__6566\,
            in2 => \N__7271\,
            in3 => \N__7619\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIGELS1_2_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7854\,
            in1 => \N__7119\,
            in2 => \_gnd_net_\,
            in3 => \N__8226\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a3_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_3_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__8322\,
            in1 => \N__8015\,
            in2 => \N__6545\,
            in3 => \N__8473\,
            lcout => \U712_CHIP_RAM.N_155\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8472\,
            in1 => \N__7120\,
            in2 => \_gnd_net_\,
            in3 => \N__8321\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000000111"
        )
    port map (
            in0 => \N__9757\,
            in1 => \N__9624\,
            in2 => \N__9486\,
            in3 => \N__9839\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_CMA28_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10979\,
            in1 => \_gnd_net_\,
            in2 => \N__6527\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LMBE_i_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111001011101"
        )
    port map (
            in0 => \N__7009\,
            in1 => \N__6934\,
            in2 => \N__6875\,
            in3 => \N__6822\,
            lcout => \U712_BYTE_ENABLE.N_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_i_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010101111"
        )
    port map (
            in0 => \N__6933\,
            in1 => \N__6863\,
            in2 => \N__6824\,
            in3 => \N__7008\,
            lcout => \U712_BYTE_ENABLE.N_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UMBE_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001010"
        )
    port map (
            in0 => \N__7010\,
            in1 => \N__6935\,
            in2 => \N__6876\,
            in3 => \N__6823\,
            lcout => \UMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_56_i_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100101010"
        )
    port map (
            in0 => \N__7012\,
            in1 => \N__6930\,
            in2 => \N__6895\,
            in3 => \N__6815\,
            lcout => \N_56_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_58_i_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000110100010"
        )
    port map (
            in0 => \N__7013\,
            in1 => \N__6931\,
            in2 => \N__6896\,
            in3 => \N__6816\,
            lcout => \N_58_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DMA_LATCH_EN_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__10661\,
            in1 => \N__10584\,
            in2 => \_gnd_net_\,
            in3 => \N__10738\,
            lcout => \DMA_LATCH_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8042\,
            in1 => \N__7270\,
            in2 => \_gnd_net_\,
            in3 => \N__7396\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10297\,
            ce => \N__6710\,
            sr => \N__10930\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6701\,
            in1 => \N__6683\,
            in2 => \_gnd_net_\,
            in3 => \N__9660\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__6668\,
            in1 => \_gnd_net_\,
            in2 => \N__9690\,
            in3 => \N__6647\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6632\,
            in1 => \N__6617\,
            in2 => \_gnd_net_\,
            in3 => \N__9659\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__9313\,
            in1 => \N__6598\,
            in2 => \N__7472\,
            in3 => \N__10724\,
            lcout => \U712_CHIP_RAM.CPU_TACK_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNICP6N_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__7300\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7657\,
            lcout => \U712_CHIP_RAM.N_95\,
            ltout => \U712_CHIP_RAM.N_95_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNI1VCF5_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101100000000"
        )
    port map (
            in0 => \N__7257\,
            in1 => \N__7204\,
            in2 => \N__7175\,
            in3 => \N__7616\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_3_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_3_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIR7N96_2_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__8030\,
            in1 => \_gnd_net_\,
            in2 => \N__7160\,
            in3 => \N__8239\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__7762\,
            in1 => \N__10725\,
            in2 => \N__7157\,
            in3 => \N__7154\,
            lcout => \WRITE_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7147\,
            in1 => \N__7322\,
            in2 => \N__8043\,
            in3 => \N__7124\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100010101000"
        )
    port map (
            in0 => \N__7761\,
            in1 => \N__7084\,
            in2 => \N__7100\,
            in3 => \N__7097\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7064\,
            in1 => \N__7052\,
            in2 => \_gnd_net_\,
            in3 => \N__9629\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIGMF8A_3_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7614\,
            in1 => \N__7037\,
            in2 => \_gnd_net_\,
            in3 => \N__7480\,
            lcout => \U712_CHIP_RAM.N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000100000"
        )
    port map (
            in0 => \N__7803\,
            in1 => \N__9303\,
            in2 => \N__7661\,
            in3 => \N__7676\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_3_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8027\,
            in1 => \N__8342\,
            in2 => \N__7640\,
            in3 => \N__8467\,
            lcout => \U712_CHIP_RAM.N_151\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000001010101"
        )
    port map (
            in0 => \N__7409\,
            in1 => \N__7615\,
            in2 => \N__7583\,
            in3 => \N__8026\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER17_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7564\,
            in2 => \_gnd_net_\,
            in3 => \N__7481\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER34\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__10723\,
            in1 => \_gnd_net_\,
            in2 => \N__7460\,
            in3 => \N__8025\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9628\,
            in1 => \N__7457\,
            in2 => \_gnd_net_\,
            in3 => \N__7438\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI2MJA9_1_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__7418\,
            in1 => \N__7408\,
            in2 => \_gnd_net_\,
            in3 => \N__8466\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER17_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIH9ULN_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000010111010"
        )
    port map (
            in0 => \N__8028\,
            in1 => \N__7387\,
            in2 => \N__7325\,
            in3 => \N__7321\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER19_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER19_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI7JQ5O_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__7806\,
            in1 => \_gnd_net_\,
            in2 => \N__7310\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_38_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8558\,
            in1 => \N__8551\,
            in2 => \N__8537\,
            in3 => \N__8534\,
            lcout => \U712_CHIP_RAM.N_218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__7804\,
            in1 => \N__8528\,
            in2 => \N__8516\,
            in3 => \N__8501\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10311\,
            ce => \N__8492\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__8500\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7805\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10311\,
            ce => \N__8492\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__7886\,
            in1 => \N__8477\,
            in2 => \_gnd_net_\,
            in3 => \N__8393\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_61_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__8363\,
            in1 => \N__8378\,
            in2 => \N__8381\,
            in3 => \N__9758\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010110001"
        )
    port map (
            in0 => \N__8377\,
            in1 => \N__8369\,
            in2 => \N__9863\,
            in3 => \N__8362\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110011000000"
        )
    port map (
            in0 => \N__8338\,
            in1 => \N__8240\,
            in2 => \N__8126\,
            in3 => \N__8029\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_29_i_a2_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7812\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un3_CUMBEn_1_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8719\,
            in2 => \_gnd_net_\,
            in3 => \N__8679\,
            lcout => \U712_BYTE_ENABLE.un3_CUMBEnZ0Z_1\,
            ltout => \U712_BYTE_ENABLE.un3_CUMBEnZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001101"
        )
    port map (
            in0 => \N__9308\,
            in1 => \N__8830\,
            in2 => \N__8801\,
            in3 => \N__10666\,
            lcout => \CUMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001101"
        )
    port map (
            in0 => \N__9309\,
            in1 => \N__8780\,
            in2 => \N__8753\,
            in3 => \N__10588\,
            lcout => \CUUBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un3_CLLBEn_0_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8718\,
            in2 => \_gnd_net_\,
            in3 => \N__8678\,
            lcout => \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_0\,
            ltout => \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000111"
        )
    port map (
            in0 => \N__9307\,
            in1 => \N__8645\,
            in2 => \N__8630\,
            in3 => \N__10665\,
            lcout => \CLLBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8585\,
            in1 => \N__8963\,
            in2 => \_gnd_net_\,
            in3 => \N__9014\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10310\,
            ce => \N__10177\,
            sr => \N__10926\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110101111"
        )
    port map (
            in0 => \N__11549\,
            in1 => \N__8992\,
            in2 => \N__9429\,
            in3 => \N__9324\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__8579\,
            in1 => \_gnd_net_\,
            in2 => \N__9339\,
            in3 => \N__9896\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011111010"
        )
    port map (
            in0 => \N__10399\,
            in1 => \_gnd_net_\,
            in2 => \N__9017\,
            in3 => \N__9643\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9642\,
            in1 => \N__9008\,
            in2 => \N__9342\,
            in3 => \N__11603\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__8991\,
            in1 => \N__9420\,
            in2 => \N__9341\,
            in3 => \N__11548\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9767\,
            in2 => \_gnd_net_\,
            in3 => \N__9856\,
            lcout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9641\,
            in1 => \N__8957\,
            in2 => \N__9340\,
            in3 => \N__9995\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8951\,
            in1 => \N__8933\,
            in2 => \_gnd_net_\,
            in3 => \N__9627\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9626\,
            in1 => \N__8915\,
            in2 => \_gnd_net_\,
            in3 => \N__8890\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__9756\,
            in1 => \N__9625\,
            in2 => \_gnd_net_\,
            in3 => \N__9843\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9775\,
            in1 => \N__9706\,
            in2 => \N__9499\,
            in3 => \N__9868\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10294\,
            ce => \N__10198\,
            sr => \N__10956\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__9436\,
            in1 => \N__9122\,
            in2 => \N__9344\,
            in3 => \N__9080\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10294\,
            ce => \N__10198\,
            sr => \N__10956\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11451\,
            in1 => \N__11234\,
            in2 => \_gnd_net_\,
            in3 => \N__11132\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11066\,
            ce => \N__11025\,
            sr => \N__10946\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11131\,
            in1 => \N__11233\,
            in2 => \_gnd_net_\,
            in3 => \N__11456\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__11023\,
            sr => \N__10941\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11229\,
            in1 => \N__11366\,
            in2 => \_gnd_net_\,
            in3 => \N__10133\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11067\,
            ce => \N__11021\,
            sr => \N__10931\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100100000"
        )
    port map (
            in0 => \N__9044\,
            in1 => \N__9332\,
            in2 => \N__9705\,
            in3 => \N__10398\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9035\,
            in2 => \N__9071\,
            in3 => \N__9068\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10321\,
            ce => \N__10178\,
            sr => \N__10927\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011111111"
        )
    port map (
            in0 => \N__9331\,
            in1 => \N__9043\,
            in2 => \N__10411\,
            in3 => \N__9691\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__9314\,
            in1 => \N__9029\,
            in2 => \N__9905\,
            in3 => \N__9670\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9669\,
            in1 => \N__9023\,
            in2 => \N__9343\,
            in3 => \N__9884\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_A20_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__11124\,
            in1 => \N__11288\,
            in2 => \N__9542\,
            in3 => \N__9514\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A20C_net\,
            ce => 'H',
            sr => \N__10918\
        );

    \U712_CHIP_RAM.CRCSn_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9500\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10295\,
            ce => 'H',
            sr => \N__10962\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__9437\,
            in1 => \N__9401\,
            in2 => \N__9338\,
            in3 => \N__11081\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10299\,
            ce => \N__10199\,
            sr => \N__10958\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9333\,
            in2 => \_gnd_net_\,
            in3 => \N__9699\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__9362\,
            in1 => \N__9306\,
            in2 => \N__9968\,
            in3 => \N__9686\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9304\,
            in1 => \N__9353\,
            in2 => \N__9703\,
            in3 => \N__9158\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9305\,
            in1 => \N__9173\,
            in2 => \N__9704\,
            in3 => \N__9164\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11365\,
            in1 => \N__11275\,
            in2 => \_gnd_net_\,
            in3 => \N__10132\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__11022\,
            sr => \N__10942\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__10464\,
            in1 => \N__11468\,
            in2 => \N__10435\,
            in3 => \N__9152\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10325\,
            ce => \N__10190\,
            sr => \N__10932\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__10465\,
            in1 => \N__9878\,
            in2 => \N__10436\,
            in3 => \N__9956\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10325\,
            ce => \N__10190\,
            sr => \N__10932\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__10425\,
            in1 => \N__10466\,
            in2 => \N__10004\,
            in3 => \N__9932\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10325\,
            ce => \N__10190\,
            sr => \N__10932\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11290\,
            in1 => \N__10081\,
            in2 => \_gnd_net_\,
            in3 => \N__10046\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__11026\,
            sr => \N__10928\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10045\,
            in1 => \N__11593\,
            in2 => \_gnd_net_\,
            in3 => \N__11289\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__11026\,
            sr => \N__10928\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11291\,
            in1 => \N__10131\,
            in2 => \_gnd_net_\,
            in3 => \N__10082\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__11026\,
            sr => \N__10928\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10044\,
            in1 => \N__11287\,
            in2 => \_gnd_net_\,
            in3 => \N__11594\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11069\,
            ce => \N__11028\,
            sr => \N__10925\
        );

    \U712_CHIP_RAM.WEn_LC_16_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9869\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10293\,
            ce => 'H',
            sr => \N__10966\
        );

    \U712_CHIP_RAM.RASn_LC_16_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9779\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10296\,
            ce => 'H',
            sr => \N__10964\
        );

    \U712_CHIP_RAM.CASn_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9707\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10300\,
            ce => 'H',
            sr => \N__10963\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__10455\,
            in1 => \N__11318\,
            in2 => \N__10438\,
            in3 => \N__10514\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10322\,
            ce => \N__10197\,
            sr => \N__10952\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__10454\,
            in1 => \N__10493\,
            in2 => \N__10437\,
            in3 => \N__10088\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10322\,
            ce => \N__10197\,
            sr => \N__10952\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__10456\,
            in1 => \N__11411\,
            in2 => \N__10439\,
            in3 => \N__10370\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10322\,
            ce => \N__10197\,
            sr => \N__10952\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10080\,
            in1 => \N__11274\,
            in2 => \_gnd_net_\,
            in3 => \N__10130\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11063\,
            ce => \N__11024\,
            sr => \N__10947\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11285\,
            in1 => \N__10079\,
            in2 => \_gnd_net_\,
            in3 => \N__10043\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11064\,
            ce => \N__11027\,
            sr => \N__10943\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11589\,
            in1 => \N__11283\,
            in2 => \_gnd_net_\,
            in3 => \N__11534\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__11029\,
            sr => \N__10933\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11281\,
            in1 => \N__11523\,
            in2 => \_gnd_net_\,
            in3 => \N__11492\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__11032\,
            sr => \N__10929\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11455\,
            in1 => \N__11286\,
            in2 => \_gnd_net_\,
            in3 => \N__11395\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__11030\,
            sr => \N__10955\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11284\,
            in1 => \N__11402\,
            in2 => \_gnd_net_\,
            in3 => \N__11358\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__11031\,
            sr => \N__10948\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11579\,
            in1 => \N__11282\,
            in2 => \_gnd_net_\,
            in3 => \N__11530\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11065\,
            ce => \N__11033\,
            sr => \N__10944\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11280\,
            in1 => \N__11522\,
            in2 => \_gnd_net_\,
            in3 => \N__11491\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11068\,
            ce => \N__11035\,
            sr => \N__10934\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11293\,
            in1 => \N__11447\,
            in2 => \_gnd_net_\,
            in3 => \N__11394\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11062\,
            ce => \N__11034\,
            sr => \N__10957\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11393\,
            in1 => \N__11292\,
            in2 => \_gnd_net_\,
            in3 => \N__11352\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11062\,
            ce => \N__11034\,
            sr => \N__10957\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_22_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11309\,
            in1 => \N__11279\,
            in2 => \_gnd_net_\,
            in3 => \N__11123\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11061\,
            ce => \N__11036\,
            sr => \N__10965\
        );

    \U712_BUFFERS.DRDDIR_LC_24_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011100001111"
        )
    port map (
            in0 => \N__10814\,
            in1 => \N__10558\,
            in2 => \N__10745\,
            in3 => \N__10636\,
            lcout => \DRDDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_DRDENn_LC_24_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__10637\,
            in1 => \_gnd_net_\,
            in2 => \N__10573\,
            in3 => \N__11654\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

module U110_CYCLE_TERMINATION (

    output TACKn, TEAn

);

assign TACKn = 1'bz;
assign TEAn = 1;

endmodule

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Apr 7 2025 15:46:56

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U409_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U409_TOP
entity U409_TOP is
port (
    TM : in std_logic_vector(1 downto 0);
    TT : in std_logic_vector(1 downto 0);
    D : out std_logic_vector(7 downto 0);
    A : in std_logic_vector(31 downto 1);
    TICK60 : out std_logic;
    CIACS0n : out std_logic;
    CLK6 : in std_logic;
    CLK_CIA : out std_logic;
    BUFENn : out std_logic;
    CIACS1n : out std_logic;
    TICK50 : out std_logic;
    RAMSPACEn : out std_logic;
    CLK40_IN : in std_logic;
    CLK28_IN : in std_logic;
    REGSPACEn : out std_logic;
    TSn : in std_logic;
    RTC_ENn : out std_logic;
    RESETn : in std_logic;
    OVL : in std_logic;
    TACKn : inout std_logic;
    ROMENn : out std_logic;
    PORTSIZE : out std_logic);
end U409_TOP;

-- Architecture of U409_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U409_TOP is

signal \N__7375\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3964\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3744\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3723\ : std_logic;
signal \N__3720\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3669\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3548\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3369\ : std_logic;
signal \N__3366\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3353\ : std_logic;
signal \N__3350\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3336\ : std_logic;
signal \N__3329\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3309\ : std_logic;
signal \N__3306\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3274\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3247\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3219\ : std_logic;
signal \N__3216\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3147\ : std_logic;
signal \N__3144\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3102\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3087\ : std_logic;
signal \N__3084\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3066\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3057\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3030\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3009\ : std_logic;
signal \N__3006\ : std_logic;
signal \N__3003\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2943\ : std_logic;
signal \N__2940\ : std_logic;
signal \N__2937\ : std_logic;
signal \N__2934\ : std_logic;
signal \N__2931\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2925\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2904\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2868\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \A_c_31\ : std_logic;
signal \A_c_30\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_\ : std_logic;
signal \A_c_26\ : std_logic;
signal \A_c_24\ : std_logic;
signal \A_c_27\ : std_logic;
signal \A_c_25\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_3\ : std_logic;
signal \A_c_29\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_4_cascade_\ : std_logic;
signal \A_c_28\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RTC_ENn_i\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_1\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_1_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE_AUTOVECTOR_5_cascade_\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTOR_16\ : std_logic;
signal \TT_c_1\ : std_logic;
signal \TT_c_0\ : std_logic;
signal \U409_ADDRESS_DECODE_AUTOVECTOR_4\ : std_logic;
signal \U409_TRANSFER_ACK.N_38\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3Z0Z_2_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACE_6\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENn_2_cascade_\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U409_ADDRESS_DECODE.REGISTER_SPACEZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.RANGER_SPACEZ0Z_2_cascade_\ : std_logic;
signal \A_c_19\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_1\ : std_logic;
signal \OVL_c\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RTC_ENn\ : std_logic;
signal \PORTSIZE_0_i\ : std_logic;
signal \A_c_23\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0\ : std_logic;
signal \A_c_22\ : std_logic;
signal \A_c_21\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RAMSPACEn_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE_AUTOCONFIG_SPACE_5\ : std_logic;
signal \U409_ADDRESS_DECODE_AUTOCONFIG_SPACE_7\ : std_logic;
signal \AGNUS_SPACE_0_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE_AUTOCONFIG_SPACE_6\ : std_logic;
signal \BUFENn_c\ : std_logic;
signal \TM_c_0\ : std_logic;
signal \U409_ADDRESS_DECODE.un2_REGSPACEn_0\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0\ : std_logic;
signal \TM_c_1\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_REGSPACEn_i\ : std_logic;
signal \CIA_SPACE\ : std_logic;
signal \U409_CIA.VMA_RNOZ0Z_0_cascade_\ : std_logic;
signal \U409_CIA.un1_CIA_CLK_COUNT_3_1\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_1\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_5\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_6\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_REGSPACEn\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RAMSPACEn\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS1n_i\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS0n_i\ : std_logic;
signal \CIA_ENABLE\ : std_logic;
signal \U409_CIA.CLK_CIA6_0\ : std_logic;
signal \U409_CIA.CLK_CIA6_cascade_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_2_0\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_3\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_2\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_5\ : std_logic;
signal \CLK28_IN_c_g\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_6\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_0\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_7\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_1\ : std_logic;
signal \U409_CIA.CLK_CIA6_3\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_4\ : std_logic;
signal \U409_CIA.un1_CIA_CLK_COUNT_2_1\ : std_logic;
signal \U409_CIA.CLK_CIA6_3_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_3\ : std_logic;
signal \U409_CIA.CLK_CIA_RNOZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_6_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\ : std_logic;
signal \U409_TRANSFER_ACK.m8_ns_1_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.i6_mux_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_9\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.N_4\ : std_logic;
signal \U409_TRANSFER_ACK.N_4_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_5\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\ : std_logic;
signal \CLK_CIA_c\ : std_logic;
signal \U409_CIA.VMAZ0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_EN_e_1\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_138\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\ : std_logic;
signal \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_ENZ0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U409_TRANSFER_ACK.N_18\ : std_logic;
signal \U409_TRANSFER_ACK.N_24\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a5_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\ : std_logic;
signal \ROMENn_c\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U409_ADDRESS_DECODE_ROMEN_1\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_28_4\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.IRQ_TACK_EN_nesrC_net\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1_0\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER6\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_EN_iC_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_OUTn_0_sqmuxa_0_en\ : std_logic;
signal \U409_TICK.TICK603_8_cascade_\ : std_logic;
signal \U409_TICK.TICK603_14_cascade_\ : std_logic;
signal \U409_TICK.TICK603_9_cascade_\ : std_logic;
signal \TICK60_c\ : std_logic;
signal \U409_TICK.TICK603_10_cascade_\ : std_logic;
signal \U409_TICK.TICK603_11\ : std_logic;
signal \U409_TICK.TICK603_14\ : std_logic;
signal \U409_TICK.TICK603_9\ : std_logic;
signal \U409_TICK.TICK603_10\ : std_logic;
signal \bfn_14_1_0_\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_1\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_3\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_4\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_6\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_8\ : std_logic;
signal \bfn_14_2_0_\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_9\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_10\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_11\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_13\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_0\ : std_logic;
signal \bfn_14_4_0_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_2\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_3\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_2\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_4\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_5\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_8\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_8\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_9\ : std_logic;
signal \bfn_14_5_0_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_10\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_11\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_13\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_12\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_13\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_16\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_3\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_0\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_12\ : std_logic;
signal \U409_TICK.TICK503_8_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_10\ : std_logic;
signal \U409_TICK.TICK503_14_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_2\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_16\ : std_logic;
signal \U409_TICK.TICK503_11\ : std_logic;
signal \TICK50_c\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_6\ : std_logic;
signal \U409_TICK.TICK503_9_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_7\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_4\ : std_logic;
signal \U409_TICK.TICK503_10_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_15\ : std_logic;
signal \U409_TICK.TICK503_14\ : std_logic;
signal \U409_TICK.TICK503_10\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.TICK503_9\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_14\ : std_logic;
signal \CLK6_c_g\ : std_logic;
signal \TACK_EN_i\ : std_logic;
signal \N_475_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK28_IN_wire\ : std_logic;
signal \CLK6_wire\ : std_logic;
signal \TT_wire\ : std_logic_vector(1 downto 0);
signal \D_wire\ : std_logic_vector(7 downto 0);
signal \RTC_ENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(31 downto 1);
signal \TM_wire\ : std_logic_vector(1 downto 0);
signal \CLK_CIA_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \ROMENn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \CIACS0n_wire\ : std_logic;
signal \TICK50_wire\ : std_logic;
signal \OVL_wire\ : std_logic;
signal \TICK60_wire\ : std_logic;
signal \CIACS1n_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK28_IN_wire\ <= CLK28_IN;
    \CLK6_wire\ <= CLK6;
    \TT_wire\ <= TT;
    D <= \D_wire\;
    RTC_ENn <= \RTC_ENn_wire\;
    \A_wire\ <= A;
    \TM_wire\ <= TM;
    CLK_CIA <= \CLK_CIA_wire\;
    RAMSPACEn <= \RAMSPACEn_wire\;
    ROMENn <= \ROMENn_wire\;
    \TSn_wire\ <= TSn;
    BUFENn <= \BUFENn_wire\;
    PORTSIZE <= \PORTSIZE_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    CIACS0n <= \CIACS0n_wire\;
    TICK50 <= \TICK50_wire\;
    \OVL_wire\ <= OVL;
    TICK60 <= \TICK60_wire\;
    CIACS1n <= \CIACS1n_wire\;
    REGSPACEn <= \REGSPACEn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__5529\,
            RESETB => \N__5253\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => \CLK80_OUT\
        );

    \CLK28_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__7373\,
            GLOBALBUFFEROUTPUT => \CLK28_IN_c_g\
        );

    \CLK28_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7375\,
            DIN => \N__7374\,
            DOUT => \N__7373\,
            PACKAGEPIN => \CLK28_IN_wire\
        );

    \CLK28_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7375\,
            PADOUT => \N__7374\,
            PADIN => \N__7373\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK6_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__7363\,
            GLOBALBUFFEROUTPUT => \CLK6_c_g\
        );

    \CLK6_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7365\,
            DIN => \N__7364\,
            DOUT => \N__7363\,
            PACKAGEPIN => \CLK6_wire\
        );

    \CLK6_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7365\,
            PADOUT => \N__7364\,
            PADIN => \N__7363\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7354\,
            DIN => \N__7353\,
            DOUT => \N__7352\,
            PACKAGEPIN => \TT_wire\(0)
        );

    \TT_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7354\,
            PADOUT => \N__7353\,
            PADIN => \N__7352\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7345\,
            DIN => \N__7344\,
            DOUT => \N__7343\,
            PACKAGEPIN => \D_wire\(6)
        );

    \D_obuft_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7345\,
            PADOUT => \N__7344\,
            PADIN => \N__7343\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RTC_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7336\,
            DIN => \N__7335\,
            DOUT => \N__7334\,
            PACKAGEPIN => \RTC_ENn_wire\
        );

    \RTC_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7336\,
            PADOUT => \N__7335\,
            PADIN => \N__7334\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2934\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7327\,
            DIN => \N__7326\,
            DOUT => \N__7325\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7327\,
            PADOUT => \N__7326\,
            PADIN => \N__7325\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7318\,
            DIN => \N__7317\,
            DOUT => \N__7316\,
            PACKAGEPIN => \D_wire\(5)
        );

    \D_obuft_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7318\,
            PADOUT => \N__7317\,
            PADIN => \N__7316\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TM_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7309\,
            DIN => \N__7308\,
            DOUT => \N__7307\,
            PACKAGEPIN => \TM_wire\(1)
        );

    \TM_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7309\,
            PADOUT => \N__7308\,
            PADIN => \N__7307\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TM_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7300\,
            DIN => \N__7299\,
            DOUT => \N__7298\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7300\,
            PADOUT => \N__7299\,
            PADIN => \N__7298\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_CIA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7291\,
            DIN => \N__7290\,
            DOUT => \N__7289\,
            PACKAGEPIN => \CLK_CIA_wire\
        );

    \CLK_CIA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7291\,
            PADOUT => \N__7290\,
            PADIN => \N__7289\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4920\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7282\,
            DIN => \N__7281\,
            DOUT => \N__7280\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7282\,
            PADOUT => \N__7281\,
            PADIN => \N__7280\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7273\,
            DIN => \N__7272\,
            DOUT => \N__7271\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7273\,
            PADOUT => \N__7272\,
            PADIN => \N__7271\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4044\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7264\,
            DIN => \N__7263\,
            DOUT => \N__7262\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7264\,
            PADOUT => \N__7263\,
            PADIN => \N__7262\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6726\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__5319\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7255\,
            DIN => \N__7254\,
            DOUT => \N__7253\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7255\,
            PADOUT => \N__7254\,
            PADIN => \N__7253\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ROMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7246\,
            DIN => \N__7245\,
            DOUT => \N__7244\,
            PACKAGEPIN => \ROMENn_wire\
        );

    \ROMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7246\,
            PADOUT => \N__7245\,
            PADIN => \N__7244\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5193\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7237\,
            DIN => \N__7236\,
            DOUT => \N__7235\,
            PACKAGEPIN => \D_wire\(0)
        );

    \D_obuft_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7237\,
            PADOUT => \N__7236\,
            PADIN => \N__7235\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7228\,
            DIN => \N__7227\,
            DOUT => \N__7226\,
            PACKAGEPIN => \TT_wire\(1)
        );

    \TT_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7228\,
            PADOUT => \N__7227\,
            PADIN => \N__7226\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7219\,
            DIN => \N__7218\,
            DOUT => \N__7217\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7219\,
            PADOUT => \N__7218\,
            PADIN => \N__7217\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7210\,
            DIN => \N__7209\,
            DOUT => \N__7208\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7210\,
            PADOUT => \N__7209\,
            PADIN => \N__7208\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3717\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7201\,
            DIN => \N__7200\,
            DOUT => \N__7199\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7201\,
            PADOUT => \N__7200\,
            PADIN => \N__7199\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4002\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7192\,
            DIN => \N__7191\,
            DOUT => \N__7190\,
            PACKAGEPIN => \D_wire\(7)
        );

    \D_obuft_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7192\,
            PADOUT => \N__7191\,
            PADIN => \N__7190\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7183\,
            DIN => \N__7182\,
            DOUT => \N__7181\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7183\,
            PADOUT => \N__7182\,
            PADIN => \N__7181\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7174\,
            DIN => \N__7173\,
            DOUT => \N__7172\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7174\,
            PADOUT => \N__7173\,
            PADIN => \N__7172\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7165\,
            DIN => \N__7164\,
            DOUT => \N__7163\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7165\,
            PADOUT => \N__7164\,
            PADIN => \N__7163\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7156\,
            DIN => \N__7155\,
            DOUT => \N__7154\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7156\,
            PADOUT => \N__7155\,
            PADIN => \N__7154\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7147\,
            DIN => \N__7146\,
            DOUT => \N__7145\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7147\,
            PADOUT => \N__7146\,
            PADIN => \N__7145\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7138\,
            DIN => \N__7137\,
            DOUT => \N__7136\,
            PACKAGEPIN => \D_wire\(2)
        );

    \D_obuft_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7138\,
            PADOUT => \N__7137\,
            PADIN => \N__7136\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7129\,
            DIN => \N__7128\,
            DOUT => \N__7127\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7129\,
            PADOUT => \N__7128\,
            PADIN => \N__7127\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TM_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7120\,
            DIN => \N__7119\,
            DOUT => \N__7118\,
            PACKAGEPIN => \TM_wire\(0)
        );

    \TM_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7120\,
            PADOUT => \N__7119\,
            PADIN => \N__7118\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TM_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7111\,
            DIN => \N__7110\,
            DOUT => \N__7109\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7111\,
            PADOUT => \N__7110\,
            PADIN => \N__7109\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7102\,
            DIN => \N__7101\,
            DOUT => \N__7100\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7102\,
            PADOUT => \N__7101\,
            PADIN => \N__7100\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7093\,
            DIN => \N__7092\,
            DOUT => \N__7091\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7093\,
            PADOUT => \N__7092\,
            PADIN => \N__7091\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7084\,
            DIN => \N__7083\,
            DOUT => \N__7082\,
            PACKAGEPIN => \D_wire\(1)
        );

    \D_obuft_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7084\,
            PADOUT => \N__7083\,
            PADIN => \N__7082\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS0n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7075\,
            DIN => \N__7074\,
            DOUT => \N__7073\,
            PACKAGEPIN => \CIACS0n_wire\
        );

    \CIACS0n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7075\,
            PADOUT => \N__7074\,
            PADIN => \N__7073\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4311\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7066\,
            DIN => \N__7065\,
            DOUT => \N__7064\,
            PACKAGEPIN => \D_wire\(4)
        );

    \D_obuft_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7066\,
            PADOUT => \N__7065\,
            PADIN => \N__7064\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK50_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7057\,
            DIN => \N__7056\,
            DOUT => \N__7055\,
            PACKAGEPIN => \TICK50_wire\
        );

    \TICK50_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7057\,
            PADOUT => \N__7056\,
            PADIN => \N__7055\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6624\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7048\,
            DIN => \N__7047\,
            DOUT => \N__7046\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7048\,
            PADOUT => \N__7047\,
            PADIN => \N__7046\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7039\,
            DIN => \N__7038\,
            DOUT => \N__7037\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7039\,
            PADOUT => \N__7038\,
            PADIN => \N__7037\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7030\,
            DIN => \N__7029\,
            DOUT => \N__7028\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7030\,
            PADOUT => \N__7029\,
            PADIN => \N__7028\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \OVL_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7021\,
            DIN => \N__7020\,
            DOUT => \N__7019\,
            PACKAGEPIN => \OVL_wire\
        );

    \OVL_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7021\,
            PADOUT => \N__7020\,
            PADIN => \N__7019\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \OVL_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7012\,
            DIN => \N__7011\,
            DOUT => \N__7010\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7012\,
            PADOUT => \N__7011\,
            PADIN => \N__7010\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK60_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7003\,
            DIN => \N__7002\,
            DOUT => \N__7001\,
            PACKAGEPIN => \TICK60_wire\
        );

    \TICK60_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7003\,
            PADOUT => \N__7002\,
            PADIN => \N__7001\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6072\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6994\,
            DIN => \N__6993\,
            DOUT => \N__6992\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6994\,
            PADOUT => \N__6993\,
            PADIN => \N__6992\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6985\,
            DIN => \N__6984\,
            DOUT => \N__6983\,
            PACKAGEPIN => \D_wire\(3)
        );

    \D_obuft_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__6985\,
            PADOUT => \N__6984\,
            PADIN => \N__6983\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6976\,
            DIN => \N__6975\,
            DOUT => \N__6974\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6976\,
            PADOUT => \N__6975\,
            PADIN => \N__6974\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6967\,
            DIN => \N__6966\,
            DOUT => \N__6965\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6967\,
            PADOUT => \N__6966\,
            PADIN => \N__6965\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS1n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6958\,
            DIN => \N__6957\,
            DOUT => \N__6956\,
            PACKAGEPIN => \CIACS1n_wire\
        );

    \CIACS1n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6958\,
            PADOUT => \N__6957\,
            PADIN => \N__6956\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4149\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6949\,
            DIN => \N__6948\,
            DOUT => \N__6947\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6949\,
            PADOUT => \N__6948\,
            PADIN => \N__6947\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3489\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1603\ : InMux
    port map (
            O => \N__6930\,
            I => \N__6927\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__6927\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_15\
        );

    \I__1601\ : InMux
    port map (
            O => \N__6924\,
            I => \N__6920\
        );

    \I__1600\ : InMux
    port map (
            O => \N__6923\,
            I => \N__6917\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__6920\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__6917\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__1597\ : InMux
    port map (
            O => \N__6912\,
            I => \N__6894\
        );

    \I__1596\ : InMux
    port map (
            O => \N__6911\,
            I => \N__6894\
        );

    \I__1595\ : InMux
    port map (
            O => \N__6910\,
            I => \N__6894\
        );

    \I__1594\ : InMux
    port map (
            O => \N__6909\,
            I => \N__6894\
        );

    \I__1593\ : InMux
    port map (
            O => \N__6908\,
            I => \N__6894\
        );

    \I__1592\ : InMux
    port map (
            O => \N__6907\,
            I => \N__6887\
        );

    \I__1591\ : InMux
    port map (
            O => \N__6906\,
            I => \N__6887\
        );

    \I__1590\ : InMux
    port map (
            O => \N__6905\,
            I => \N__6887\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__6894\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__6887\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1587\ : InMux
    port map (
            O => \N__6882\,
            I => \N__6866\
        );

    \I__1586\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6866\
        );

    \I__1585\ : InMux
    port map (
            O => \N__6880\,
            I => \N__6866\
        );

    \I__1584\ : InMux
    port map (
            O => \N__6879\,
            I => \N__6866\
        );

    \I__1583\ : InMux
    port map (
            O => \N__6878\,
            I => \N__6857\
        );

    \I__1582\ : InMux
    port map (
            O => \N__6877\,
            I => \N__6857\
        );

    \I__1581\ : InMux
    port map (
            O => \N__6876\,
            I => \N__6857\
        );

    \I__1580\ : InMux
    port map (
            O => \N__6875\,
            I => \N__6857\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__6866\,
            I => \U409_TICK.TICK503_10\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__6857\,
            I => \U409_TICK.TICK503_10\
        );

    \I__1577\ : CascadeMux
    port map (
            O => \N__6852\,
            I => \N__6849\
        );

    \I__1576\ : InMux
    port map (
            O => \N__6849\,
            I => \N__6846\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__6846\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_14\
        );

    \I__1574\ : CascadeMux
    port map (
            O => \N__6843\,
            I => \N__6840\
        );

    \I__1573\ : InMux
    port map (
            O => \N__6840\,
            I => \N__6830\
        );

    \I__1572\ : InMux
    port map (
            O => \N__6839\,
            I => \N__6830\
        );

    \I__1571\ : CascadeMux
    port map (
            O => \N__6838\,
            I => \N__6827\
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__6837\,
            I => \N__6824\
        );

    \I__1569\ : CascadeMux
    port map (
            O => \N__6836\,
            I => \N__6821\
        );

    \I__1568\ : CascadeMux
    port map (
            O => \N__6835\,
            I => \N__6816\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__6830\,
            I => \N__6813\
        );

    \I__1566\ : InMux
    port map (
            O => \N__6827\,
            I => \N__6808\
        );

    \I__1565\ : InMux
    port map (
            O => \N__6824\,
            I => \N__6808\
        );

    \I__1564\ : InMux
    port map (
            O => \N__6821\,
            I => \N__6799\
        );

    \I__1563\ : InMux
    port map (
            O => \N__6820\,
            I => \N__6799\
        );

    \I__1562\ : InMux
    port map (
            O => \N__6819\,
            I => \N__6799\
        );

    \I__1561\ : InMux
    port map (
            O => \N__6816\,
            I => \N__6799\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__6813\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__6808\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__6799\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__6792\,
            I => \N__6789\
        );

    \I__1556\ : InMux
    port map (
            O => \N__6789\,
            I => \N__6785\
        );

    \I__1555\ : InMux
    port map (
            O => \N__6788\,
            I => \N__6782\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__6785\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__6782\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__1552\ : ClkMux
    port map (
            O => \N__6777\,
            I => \N__6750\
        );

    \I__1551\ : ClkMux
    port map (
            O => \N__6776\,
            I => \N__6750\
        );

    \I__1550\ : ClkMux
    port map (
            O => \N__6775\,
            I => \N__6750\
        );

    \I__1549\ : ClkMux
    port map (
            O => \N__6774\,
            I => \N__6750\
        );

    \I__1548\ : ClkMux
    port map (
            O => \N__6773\,
            I => \N__6750\
        );

    \I__1547\ : ClkMux
    port map (
            O => \N__6772\,
            I => \N__6750\
        );

    \I__1546\ : ClkMux
    port map (
            O => \N__6771\,
            I => \N__6750\
        );

    \I__1545\ : ClkMux
    port map (
            O => \N__6770\,
            I => \N__6750\
        );

    \I__1544\ : ClkMux
    port map (
            O => \N__6769\,
            I => \N__6750\
        );

    \I__1543\ : GlobalMux
    port map (
            O => \N__6750\,
            I => \N__6747\
        );

    \I__1542\ : gio2CtrlBuf
    port map (
            O => \N__6747\,
            I => \CLK6_c_g\
        );

    \I__1541\ : InMux
    port map (
            O => \N__6744\,
            I => \N__6741\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__6741\,
            I => \N__6738\
        );

    \I__1539\ : Span4Mux_v
    port map (
            O => \N__6738\,
            I => \N__6735\
        );

    \I__1538\ : Span4Mux_h
    port map (
            O => \N__6735\,
            I => \N__6732\
        );

    \I__1537\ : Span4Mux_h
    port map (
            O => \N__6732\,
            I => \N__6729\
        );

    \I__1536\ : Odrv4
    port map (
            O => \N__6729\,
            I => \TACK_EN_i\
        );

    \I__1535\ : IoInMux
    port map (
            O => \N__6726\,
            I => \N__6723\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__6723\,
            I => \N__6720\
        );

    \I__1533\ : Span4Mux_s1_v
    port map (
            O => \N__6720\,
            I => \N__6717\
        );

    \I__1532\ : Span4Mux_h
    port map (
            O => \N__6717\,
            I => \N__6714\
        );

    \I__1531\ : Span4Mux_v
    port map (
            O => \N__6714\,
            I => \N__6711\
        );

    \I__1530\ : Odrv4
    port map (
            O => \N__6711\,
            I => \N_475_i\
        );

    \I__1529\ : CascadeMux
    port map (
            O => \N__6708\,
            I => \U409_TICK.TICK503_14_cascade_\
        );

    \I__1528\ : InMux
    port map (
            O => \N__6705\,
            I => \N__6702\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__6702\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_5\
        );

    \I__1526\ : InMux
    port map (
            O => \N__6699\,
            I => \N__6695\
        );

    \I__1525\ : InMux
    port map (
            O => \N__6698\,
            I => \N__6692\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__6695\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__6692\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__1522\ : InMux
    port map (
            O => \N__6687\,
            I => \N__6683\
        );

    \I__1521\ : InMux
    port map (
            O => \N__6686\,
            I => \N__6680\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__6683\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__6680\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__1518\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6671\
        );

    \I__1517\ : InMux
    port map (
            O => \N__6674\,
            I => \N__6668\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__6671\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__6668\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__1514\ : CascadeMux
    port map (
            O => \N__6663\,
            I => \N__6659\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__6662\,
            I => \N__6656\
        );

    \I__1512\ : InMux
    port map (
            O => \N__6659\,
            I => \N__6650\
        );

    \I__1511\ : InMux
    port map (
            O => \N__6656\,
            I => \N__6650\
        );

    \I__1510\ : InMux
    port map (
            O => \N__6655\,
            I => \N__6647\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__6650\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__6647\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__1507\ : InMux
    port map (
            O => \N__6642\,
            I => \N__6638\
        );

    \I__1506\ : InMux
    port map (
            O => \N__6641\,
            I => \N__6635\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__6638\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__6635\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__1503\ : InMux
    port map (
            O => \N__6630\,
            I => \N__6627\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__6627\,
            I => \U409_TICK.TICK503_11\
        );

    \I__1501\ : IoInMux
    port map (
            O => \N__6624\,
            I => \N__6621\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__6621\,
            I => \N__6618\
        );

    \I__1499\ : Span4Mux_s3_v
    port map (
            O => \N__6618\,
            I => \N__6615\
        );

    \I__1498\ : Span4Mux_h
    port map (
            O => \N__6615\,
            I => \N__6611\
        );

    \I__1497\ : InMux
    port map (
            O => \N__6614\,
            I => \N__6608\
        );

    \I__1496\ : Odrv4
    port map (
            O => \N__6611\,
            I => \TICK50_c\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__6608\,
            I => \TICK50_c\
        );

    \I__1494\ : InMux
    port map (
            O => \N__6603\,
            I => \N__6600\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__6600\,
            I => \N__6597\
        );

    \I__1492\ : Odrv4
    port map (
            O => \N__6597\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_9\
        );

    \I__1491\ : InMux
    port map (
            O => \N__6594\,
            I => \N__6590\
        );

    \I__1490\ : InMux
    port map (
            O => \N__6593\,
            I => \N__6587\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__6590\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__6587\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__1487\ : CascadeMux
    port map (
            O => \N__6582\,
            I => \N__6579\
        );

    \I__1486\ : InMux
    port map (
            O => \N__6579\,
            I => \N__6575\
        );

    \I__1485\ : InMux
    port map (
            O => \N__6578\,
            I => \N__6572\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__6575\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__6572\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__1482\ : CascadeMux
    port map (
            O => \N__6567\,
            I => \U409_TICK.TICK503_9_cascade_\
        );

    \I__1481\ : InMux
    port map (
            O => \N__6564\,
            I => \N__6561\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__6561\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_13\
        );

    \I__1479\ : InMux
    port map (
            O => \N__6558\,
            I => \N__6554\
        );

    \I__1478\ : InMux
    port map (
            O => \N__6557\,
            I => \N__6551\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__6554\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__6551\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__1475\ : InMux
    port map (
            O => \N__6546\,
            I => \N__6542\
        );

    \I__1474\ : InMux
    port map (
            O => \N__6545\,
            I => \N__6539\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__6542\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__6539\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__1471\ : InMux
    port map (
            O => \N__6534\,
            I => \N__6530\
        );

    \I__1470\ : InMux
    port map (
            O => \N__6533\,
            I => \N__6527\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__6530\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__6527\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__1467\ : CascadeMux
    port map (
            O => \N__6522\,
            I => \U409_TICK.TICK503_10_cascade_\
        );

    \I__1466\ : InMux
    port map (
            O => \N__6519\,
            I => \N__6516\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__6516\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_11\
        );

    \I__1464\ : InMux
    port map (
            O => \N__6513\,
            I => \N__6509\
        );

    \I__1463\ : InMux
    port map (
            O => \N__6512\,
            I => \N__6506\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__6509\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__6506\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__1460\ : InMux
    port map (
            O => \N__6501\,
            I => \N__6497\
        );

    \I__1459\ : InMux
    port map (
            O => \N__6500\,
            I => \N__6494\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__6497\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__6494\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__1456\ : InMux
    port map (
            O => \N__6489\,
            I => \U409_TICK.un3_COUNTER60_1_cry_12\
        );

    \I__1455\ : InMux
    port map (
            O => \N__6486\,
            I => \N__6482\
        );

    \I__1454\ : InMux
    port map (
            O => \N__6485\,
            I => \N__6479\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__6482\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__6479\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__1451\ : InMux
    port map (
            O => \N__6474\,
            I => \N__6471\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__6471\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_14\
        );

    \I__1449\ : InMux
    port map (
            O => \N__6468\,
            I => \U409_TICK.un3_COUNTER60_1_cry_13\
        );

    \I__1448\ : InMux
    port map (
            O => \N__6465\,
            I => \N__6461\
        );

    \I__1447\ : InMux
    port map (
            O => \N__6464\,
            I => \N__6458\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__6461\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__6458\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__1444\ : InMux
    port map (
            O => \N__6453\,
            I => \N__6450\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__6450\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_15\
        );

    \I__1442\ : InMux
    port map (
            O => \N__6447\,
            I => \U409_TICK.un3_COUNTER60_1_cry_14\
        );

    \I__1441\ : InMux
    port map (
            O => \N__6444\,
            I => \U409_TICK.un3_COUNTER60_1_cry_15\
        );

    \I__1440\ : InMux
    port map (
            O => \N__6441\,
            I => \N__6437\
        );

    \I__1439\ : InMux
    port map (
            O => \N__6440\,
            I => \N__6434\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__6437\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__6434\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__1436\ : InMux
    port map (
            O => \N__6429\,
            I => \N__6426\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__6426\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_6\
        );

    \I__1434\ : InMux
    port map (
            O => \N__6423\,
            I => \N__6419\
        );

    \I__1433\ : InMux
    port map (
            O => \N__6422\,
            I => \N__6416\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__6419\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__6416\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__1430\ : CascadeMux
    port map (
            O => \N__6411\,
            I => \N__6405\
        );

    \I__1429\ : InMux
    port map (
            O => \N__6410\,
            I => \N__6398\
        );

    \I__1428\ : InMux
    port map (
            O => \N__6409\,
            I => \N__6398\
        );

    \I__1427\ : InMux
    port map (
            O => \N__6408\,
            I => \N__6398\
        );

    \I__1426\ : InMux
    port map (
            O => \N__6405\,
            I => \N__6395\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__6398\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__6395\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__1423\ : InMux
    port map (
            O => \N__6390\,
            I => \N__6386\
        );

    \I__1422\ : InMux
    port map (
            O => \N__6389\,
            I => \N__6383\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__6386\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__6383\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__6378\,
            I => \U409_TICK.TICK503_8_cascade_\
        );

    \I__1418\ : InMux
    port map (
            O => \N__6375\,
            I => \N__6371\
        );

    \I__1417\ : InMux
    port map (
            O => \N__6374\,
            I => \N__6368\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__6371\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__6368\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__1414\ : InMux
    port map (
            O => \N__6363\,
            I => \N__6359\
        );

    \I__1413\ : InMux
    port map (
            O => \N__6362\,
            I => \N__6356\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__6359\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__6356\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__1410\ : InMux
    port map (
            O => \N__6351\,
            I => \U409_TICK.un3_COUNTER60_1_cry_4\
        );

    \I__1409\ : InMux
    port map (
            O => \N__6348\,
            I => \N__6344\
        );

    \I__1408\ : InMux
    port map (
            O => \N__6347\,
            I => \N__6341\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__6344\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__6341\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__1405\ : InMux
    port map (
            O => \N__6336\,
            I => \N__6333\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__6333\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_6\
        );

    \I__1403\ : InMux
    port map (
            O => \N__6330\,
            I => \U409_TICK.un3_COUNTER60_1_cry_5\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__6327\,
            I => \N__6324\
        );

    \I__1401\ : InMux
    port map (
            O => \N__6324\,
            I => \N__6320\
        );

    \I__1400\ : InMux
    port map (
            O => \N__6323\,
            I => \N__6317\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__6320\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__6317\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__1397\ : InMux
    port map (
            O => \N__6312\,
            I => \U409_TICK.un3_COUNTER60_1_cry_6\
        );

    \I__1396\ : CascadeMux
    port map (
            O => \N__6309\,
            I => \N__6306\
        );

    \I__1395\ : InMux
    port map (
            O => \N__6306\,
            I => \N__6302\
        );

    \I__1394\ : InMux
    port map (
            O => \N__6305\,
            I => \N__6299\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__6302\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__6299\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__1391\ : InMux
    port map (
            O => \N__6294\,
            I => \N__6291\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__6291\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_8\
        );

    \I__1389\ : InMux
    port map (
            O => \N__6288\,
            I => \U409_TICK.un3_COUNTER60_1_cry_7\
        );

    \I__1388\ : InMux
    port map (
            O => \N__6285\,
            I => \N__6281\
        );

    \I__1387\ : InMux
    port map (
            O => \N__6284\,
            I => \N__6278\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__6281\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__6278\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__6273\,
            I => \N__6270\
        );

    \I__1383\ : InMux
    port map (
            O => \N__6270\,
            I => \N__6267\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__6267\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_9\
        );

    \I__1381\ : InMux
    port map (
            O => \N__6264\,
            I => \bfn_14_5_0_\
        );

    \I__1380\ : InMux
    port map (
            O => \N__6261\,
            I => \N__6257\
        );

    \I__1379\ : InMux
    port map (
            O => \N__6260\,
            I => \N__6254\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__6257\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__6254\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__1376\ : InMux
    port map (
            O => \N__6249\,
            I => \U409_TICK.un3_COUNTER60_1_cry_9\
        );

    \I__1375\ : InMux
    port map (
            O => \N__6246\,
            I => \N__6242\
        );

    \I__1374\ : InMux
    port map (
            O => \N__6245\,
            I => \N__6239\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__6242\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__6239\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__1371\ : InMux
    port map (
            O => \N__6234\,
            I => \U409_TICK.un3_COUNTER60_1_cry_10\
        );

    \I__1370\ : InMux
    port map (
            O => \N__6231\,
            I => \N__6227\
        );

    \I__1369\ : InMux
    port map (
            O => \N__6230\,
            I => \N__6224\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__6227\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__6224\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__1366\ : InMux
    port map (
            O => \N__6219\,
            I => \U409_TICK.un3_COUNTER60_1_cry_11\
        );

    \I__1365\ : InMux
    port map (
            O => \N__6216\,
            I => \U409_TICK.un2_COUNTER50_1_cry_11\
        );

    \I__1364\ : InMux
    port map (
            O => \N__6213\,
            I => \U409_TICK.un2_COUNTER50_1_cry_12\
        );

    \I__1363\ : InMux
    port map (
            O => \N__6210\,
            I => \U409_TICK.un2_COUNTER50_1_cry_13\
        );

    \I__1362\ : InMux
    port map (
            O => \N__6207\,
            I => \U409_TICK.un2_COUNTER50_1_cry_14\
        );

    \I__1361\ : InMux
    port map (
            O => \N__6204\,
            I => \U409_TICK.un2_COUNTER50_1_cry_15\
        );

    \I__1360\ : CascadeMux
    port map (
            O => \N__6201\,
            I => \N__6197\
        );

    \I__1359\ : CascadeMux
    port map (
            O => \N__6200\,
            I => \N__6194\
        );

    \I__1358\ : InMux
    port map (
            O => \N__6197\,
            I => \N__6190\
        );

    \I__1357\ : InMux
    port map (
            O => \N__6194\,
            I => \N__6187\
        );

    \I__1356\ : InMux
    port map (
            O => \N__6193\,
            I => \N__6184\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__6190\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__6187\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__6184\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__1352\ : CascadeMux
    port map (
            O => \N__6177\,
            I => \N__6171\
        );

    \I__1351\ : InMux
    port map (
            O => \N__6176\,
            I => \N__6164\
        );

    \I__1350\ : InMux
    port map (
            O => \N__6175\,
            I => \N__6164\
        );

    \I__1349\ : InMux
    port map (
            O => \N__6174\,
            I => \N__6164\
        );

    \I__1348\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6161\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__6164\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__6161\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__1345\ : InMux
    port map (
            O => \N__6156\,
            I => \N__6152\
        );

    \I__1344\ : InMux
    port map (
            O => \N__6155\,
            I => \N__6149\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__6152\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__6149\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__1341\ : InMux
    port map (
            O => \N__6144\,
            I => \U409_TICK.un3_COUNTER60_1_cry_1\
        );

    \I__1340\ : InMux
    port map (
            O => \N__6141\,
            I => \N__6137\
        );

    \I__1339\ : InMux
    port map (
            O => \N__6140\,
            I => \N__6134\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__6137\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__6134\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__1336\ : InMux
    port map (
            O => \N__6129\,
            I => \U409_TICK.un3_COUNTER60_1_cry_2\
        );

    \I__1335\ : InMux
    port map (
            O => \N__6126\,
            I => \N__6122\
        );

    \I__1334\ : InMux
    port map (
            O => \N__6125\,
            I => \N__6119\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__6122\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__6119\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__1331\ : CascadeMux
    port map (
            O => \N__6114\,
            I => \N__6111\
        );

    \I__1330\ : InMux
    port map (
            O => \N__6111\,
            I => \N__6108\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__6108\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_4\
        );

    \I__1328\ : InMux
    port map (
            O => \N__6105\,
            I => \U409_TICK.un3_COUNTER60_1_cry_3\
        );

    \I__1327\ : InMux
    port map (
            O => \N__6102\,
            I => \U409_TICK.un2_COUNTER50_1_cry_2\
        );

    \I__1326\ : InMux
    port map (
            O => \N__6099\,
            I => \U409_TICK.un2_COUNTER50_1_cry_3\
        );

    \I__1325\ : InMux
    port map (
            O => \N__6096\,
            I => \U409_TICK.un2_COUNTER50_1_cry_4\
        );

    \I__1324\ : InMux
    port map (
            O => \N__6093\,
            I => \U409_TICK.un2_COUNTER50_1_cry_5\
        );

    \I__1323\ : InMux
    port map (
            O => \N__6090\,
            I => \U409_TICK.un2_COUNTER50_1_cry_6\
        );

    \I__1322\ : InMux
    port map (
            O => \N__6087\,
            I => \U409_TICK.un2_COUNTER50_1_cry_7\
        );

    \I__1321\ : InMux
    port map (
            O => \N__6084\,
            I => \bfn_14_2_0_\
        );

    \I__1320\ : InMux
    port map (
            O => \N__6081\,
            I => \U409_TICK.un2_COUNTER50_1_cry_9\
        );

    \I__1319\ : InMux
    port map (
            O => \N__6078\,
            I => \U409_TICK.un2_COUNTER50_1_cry_10\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__6075\,
            I => \U409_TICK.TICK603_9_cascade_\
        );

    \I__1317\ : IoInMux
    port map (
            O => \N__6072\,
            I => \N__6069\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__6069\,
            I => \N__6066\
        );

    \I__1315\ : Span4Mux_s3_v
    port map (
            O => \N__6066\,
            I => \N__6063\
        );

    \I__1314\ : Span4Mux_v
    port map (
            O => \N__6063\,
            I => \N__6060\
        );

    \I__1313\ : Span4Mux_h
    port map (
            O => \N__6060\,
            I => \N__6056\
        );

    \I__1312\ : InMux
    port map (
            O => \N__6059\,
            I => \N__6053\
        );

    \I__1311\ : Odrv4
    port map (
            O => \N__6056\,
            I => \TICK60_c\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__6053\,
            I => \TICK60_c\
        );

    \I__1309\ : CascadeMux
    port map (
            O => \N__6048\,
            I => \U409_TICK.TICK603_10_cascade_\
        );

    \I__1308\ : InMux
    port map (
            O => \N__6045\,
            I => \N__6042\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__6042\,
            I => \U409_TICK.TICK603_11\
        );

    \I__1306\ : InMux
    port map (
            O => \N__6039\,
            I => \N__6030\
        );

    \I__1305\ : InMux
    port map (
            O => \N__6038\,
            I => \N__6023\
        );

    \I__1304\ : InMux
    port map (
            O => \N__6037\,
            I => \N__6023\
        );

    \I__1303\ : InMux
    port map (
            O => \N__6036\,
            I => \N__6023\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6035\,
            I => \N__6016\
        );

    \I__1301\ : InMux
    port map (
            O => \N__6034\,
            I => \N__6016\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6033\,
            I => \N__6016\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__6030\,
            I => \U409_TICK.TICK603_14\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__6023\,
            I => \U409_TICK.TICK603_14\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__6016\,
            I => \U409_TICK.TICK603_14\
        );

    \I__1296\ : CascadeMux
    port map (
            O => \N__6009\,
            I => \N__6002\
        );

    \I__1295\ : InMux
    port map (
            O => \N__6008\,
            I => \N__5997\
        );

    \I__1294\ : InMux
    port map (
            O => \N__6007\,
            I => \N__5990\
        );

    \I__1293\ : InMux
    port map (
            O => \N__6006\,
            I => \N__5990\
        );

    \I__1292\ : InMux
    port map (
            O => \N__6005\,
            I => \N__5990\
        );

    \I__1291\ : InMux
    port map (
            O => \N__6002\,
            I => \N__5983\
        );

    \I__1290\ : InMux
    port map (
            O => \N__6001\,
            I => \N__5983\
        );

    \I__1289\ : InMux
    port map (
            O => \N__6000\,
            I => \N__5983\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__5997\,
            I => \U409_TICK.TICK603_9\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__5990\,
            I => \U409_TICK.TICK603_9\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__5983\,
            I => \U409_TICK.TICK603_9\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__5976\,
            I => \N__5972\
        );

    \I__1284\ : CascadeMux
    port map (
            O => \N__5975\,
            I => \N__5969\
        );

    \I__1283\ : InMux
    port map (
            O => \N__5972\,
            I => \N__5961\
        );

    \I__1282\ : InMux
    port map (
            O => \N__5969\,
            I => \N__5956\
        );

    \I__1281\ : InMux
    port map (
            O => \N__5968\,
            I => \N__5956\
        );

    \I__1280\ : InMux
    port map (
            O => \N__5967\,
            I => \N__5947\
        );

    \I__1279\ : InMux
    port map (
            O => \N__5966\,
            I => \N__5947\
        );

    \I__1278\ : InMux
    port map (
            O => \N__5965\,
            I => \N__5947\
        );

    \I__1277\ : InMux
    port map (
            O => \N__5964\,
            I => \N__5947\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__5961\,
            I => \N__5944\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__5956\,
            I => \U409_TICK.TICK603_10\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__5947\,
            I => \U409_TICK.TICK603_10\
        );

    \I__1273\ : Odrv4
    port map (
            O => \N__5944\,
            I => \U409_TICK.TICK603_10\
        );

    \I__1272\ : InMux
    port map (
            O => \N__5937\,
            I => \U409_TICK.un2_COUNTER50_1_cry_1\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__5934\,
            I => \N__5927\
        );

    \I__1270\ : CascadeMux
    port map (
            O => \N__5933\,
            I => \N__5924\
        );

    \I__1269\ : InMux
    port map (
            O => \N__5932\,
            I => \N__5921\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5931\,
            I => \N__5912\
        );

    \I__1267\ : InMux
    port map (
            O => \N__5930\,
            I => \N__5912\
        );

    \I__1266\ : InMux
    port map (
            O => \N__5927\,
            I => \N__5912\
        );

    \I__1265\ : InMux
    port map (
            O => \N__5924\,
            I => \N__5912\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__5921\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__5912\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1262\ : InMux
    port map (
            O => \N__5907\,
            I => \N__5900\
        );

    \I__1261\ : InMux
    port map (
            O => \N__5906\,
            I => \N__5891\
        );

    \I__1260\ : InMux
    port map (
            O => \N__5905\,
            I => \N__5891\
        );

    \I__1259\ : InMux
    port map (
            O => \N__5904\,
            I => \N__5891\
        );

    \I__1258\ : InMux
    port map (
            O => \N__5903\,
            I => \N__5891\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__5900\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__5891\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1255\ : InMux
    port map (
            O => \N__5886\,
            I => \N__5882\
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__5885\,
            I => \N__5879\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__5882\,
            I => \N__5874\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5879\,
            I => \N__5871\
        );

    \I__1251\ : InMux
    port map (
            O => \N__5878\,
            I => \N__5867\
        );

    \I__1250\ : CascadeMux
    port map (
            O => \N__5877\,
            I => \N__5864\
        );

    \I__1249\ : Span4Mux_v
    port map (
            O => \N__5874\,
            I => \N__5861\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__5871\,
            I => \N__5858\
        );

    \I__1247\ : InMux
    port map (
            O => \N__5870\,
            I => \N__5855\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__5867\,
            I => \N__5852\
        );

    \I__1245\ : InMux
    port map (
            O => \N__5864\,
            I => \N__5849\
        );

    \I__1244\ : Span4Mux_h
    port map (
            O => \N__5861\,
            I => \N__5839\
        );

    \I__1243\ : Span4Mux_v
    port map (
            O => \N__5858\,
            I => \N__5839\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__5855\,
            I => \N__5839\
        );

    \I__1241\ : Span4Mux_h
    port map (
            O => \N__5852\,
            I => \N__5832\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__5849\,
            I => \N__5832\
        );

    \I__1239\ : CascadeMux
    port map (
            O => \N__5848\,
            I => \N__5829\
        );

    \I__1238\ : CascadeMux
    port map (
            O => \N__5847\,
            I => \N__5823\
        );

    \I__1237\ : CascadeMux
    port map (
            O => \N__5846\,
            I => \N__5819\
        );

    \I__1236\ : Span4Mux_v
    port map (
            O => \N__5839\,
            I => \N__5816\
        );

    \I__1235\ : InMux
    port map (
            O => \N__5838\,
            I => \N__5813\
        );

    \I__1234\ : InMux
    port map (
            O => \N__5837\,
            I => \N__5810\
        );

    \I__1233\ : Span4Mux_h
    port map (
            O => \N__5832\,
            I => \N__5807\
        );

    \I__1232\ : InMux
    port map (
            O => \N__5829\,
            I => \N__5804\
        );

    \I__1231\ : InMux
    port map (
            O => \N__5828\,
            I => \N__5801\
        );

    \I__1230\ : InMux
    port map (
            O => \N__5827\,
            I => \N__5794\
        );

    \I__1229\ : InMux
    port map (
            O => \N__5826\,
            I => \N__5794\
        );

    \I__1228\ : InMux
    port map (
            O => \N__5823\,
            I => \N__5794\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5822\,
            I => \N__5789\
        );

    \I__1226\ : InMux
    port map (
            O => \N__5819\,
            I => \N__5789\
        );

    \I__1225\ : Sp12to4
    port map (
            O => \N__5816\,
            I => \N__5785\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__5813\,
            I => \N__5780\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__5810\,
            I => \N__5780\
        );

    \I__1222\ : Sp12to4
    port map (
            O => \N__5807\,
            I => \N__5771\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__5804\,
            I => \N__5771\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__5801\,
            I => \N__5771\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__5794\,
            I => \N__5771\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__5789\,
            I => \N__5768\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5788\,
            I => \N__5765\
        );

    \I__1216\ : Span12Mux_h
    port map (
            O => \N__5785\,
            I => \N__5762\
        );

    \I__1215\ : Span4Mux_v
    port map (
            O => \N__5780\,
            I => \N__5759\
        );

    \I__1214\ : Span12Mux_v
    port map (
            O => \N__5771\,
            I => \N__5752\
        );

    \I__1213\ : Sp12to4
    port map (
            O => \N__5768\,
            I => \N__5752\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__5765\,
            I => \N__5752\
        );

    \I__1211\ : Span12Mux_v
    port map (
            O => \N__5762\,
            I => \N__5749\
        );

    \I__1210\ : Sp12to4
    port map (
            O => \N__5759\,
            I => \N__5746\
        );

    \I__1209\ : Span12Mux_v
    port map (
            O => \N__5752\,
            I => \N__5743\
        );

    \I__1208\ : Span12Mux_h
    port map (
            O => \N__5749\,
            I => \N__5740\
        );

    \I__1207\ : Span12Mux_h
    port map (
            O => \N__5746\,
            I => \N__5737\
        );

    \I__1206\ : Span12Mux_h
    port map (
            O => \N__5743\,
            I => \N__5734\
        );

    \I__1205\ : Odrv12
    port map (
            O => \N__5740\,
            I => \RESETn_c\
        );

    \I__1204\ : Odrv12
    port map (
            O => \N__5737\,
            I => \RESETn_c\
        );

    \I__1203\ : Odrv12
    port map (
            O => \N__5734\,
            I => \RESETn_c\
        );

    \I__1202\ : InMux
    port map (
            O => \N__5727\,
            I => \N__5724\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__5724\,
            I => \N__5718\
        );

    \I__1200\ : InMux
    port map (
            O => \N__5723\,
            I => \N__5711\
        );

    \I__1199\ : InMux
    port map (
            O => \N__5722\,
            I => \N__5711\
        );

    \I__1198\ : InMux
    port map (
            O => \N__5721\,
            I => \N__5711\
        );

    \I__1197\ : Odrv4
    port map (
            O => \N__5718\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__5711\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__1195\ : CEMux
    port map (
            O => \N__5706\,
            I => \N__5703\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__5703\,
            I => \N__5700\
        );

    \I__1193\ : Odrv4
    port map (
            O => \N__5700\,
            I => \U409_TRANSFER_ACK.TACK_OUTn_0_sqmuxa_0_en\
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__5697\,
            I => \U409_TICK.TICK603_8_cascade_\
        );

    \I__1191\ : CascadeMux
    port map (
            O => \N__5694\,
            I => \U409_TICK.TICK603_14_cascade_\
        );

    \I__1190\ : CascadeMux
    port map (
            O => \N__5691\,
            I => \N__5686\
        );

    \I__1189\ : CascadeMux
    port map (
            O => \N__5690\,
            I => \N__5683\
        );

    \I__1188\ : CascadeMux
    port map (
            O => \N__5689\,
            I => \N__5678\
        );

    \I__1187\ : InMux
    port map (
            O => \N__5686\,
            I => \N__5672\
        );

    \I__1186\ : InMux
    port map (
            O => \N__5683\,
            I => \N__5672\
        );

    \I__1185\ : InMux
    port map (
            O => \N__5682\,
            I => \N__5669\
        );

    \I__1184\ : InMux
    port map (
            O => \N__5681\,
            I => \N__5662\
        );

    \I__1183\ : InMux
    port map (
            O => \N__5678\,
            I => \N__5662\
        );

    \I__1182\ : InMux
    port map (
            O => \N__5677\,
            I => \N__5662\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__5672\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__5669\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__5662\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1178\ : InMux
    port map (
            O => \N__5655\,
            I => \N__5646\
        );

    \I__1177\ : InMux
    port map (
            O => \N__5654\,
            I => \N__5639\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5653\,
            I => \N__5639\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5652\,
            I => \N__5639\
        );

    \I__1174\ : InMux
    port map (
            O => \N__5651\,
            I => \N__5632\
        );

    \I__1173\ : InMux
    port map (
            O => \N__5650\,
            I => \N__5632\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5649\,
            I => \N__5632\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__5646\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__5639\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__5632\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1168\ : InMux
    port map (
            O => \N__5625\,
            I => \N__5612\
        );

    \I__1167\ : InMux
    port map (
            O => \N__5624\,
            I => \N__5612\
        );

    \I__1166\ : InMux
    port map (
            O => \N__5623\,
            I => \N__5612\
        );

    \I__1165\ : InMux
    port map (
            O => \N__5622\,
            I => \N__5609\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5621\,
            I => \N__5606\
        );

    \I__1163\ : InMux
    port map (
            O => \N__5620\,
            I => \N__5601\
        );

    \I__1162\ : InMux
    port map (
            O => \N__5619\,
            I => \N__5601\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__5612\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__5609\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__5606\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__5601\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1157\ : CascadeMux
    port map (
            O => \N__5592\,
            I => \N__5587\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__5591\,
            I => \N__5584\
        );

    \I__1155\ : InMux
    port map (
            O => \N__5590\,
            I => \N__5580\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5587\,
            I => \N__5575\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5584\,
            I => \N__5575\
        );

    \I__1152\ : InMux
    port map (
            O => \N__5583\,
            I => \N__5572\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__5580\,
            I => \N__5568\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__5575\,
            I => \N__5563\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__5572\,
            I => \N__5563\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5571\,
            I => \N__5560\
        );

    \I__1147\ : Span4Mux_v
    port map (
            O => \N__5568\,
            I => \N__5555\
        );

    \I__1146\ : Span4Mux_v
    port map (
            O => \N__5563\,
            I => \N__5555\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__5560\,
            I => \N__5550\
        );

    \I__1144\ : Sp12to4
    port map (
            O => \N__5555\,
            I => \N__5550\
        );

    \I__1143\ : Span12Mux_h
    port map (
            O => \N__5550\,
            I => \N__5547\
        );

    \I__1142\ : Span12Mux_v
    port map (
            O => \N__5547\,
            I => \N__5544\
        );

    \I__1141\ : Odrv12
    port map (
            O => \N__5544\,
            I => \TSn_c\
        );

    \I__1140\ : InMux
    port map (
            O => \N__5541\,
            I => \N__5538\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5538\,
            I => \N__5535\
        );

    \I__1138\ : Span12Mux_h
    port map (
            O => \N__5535\,
            I => \N__5532\
        );

    \I__1137\ : Odrv12
    port map (
            O => \N__5532\,
            I => \U409_ADDRESS_DECODE_ROMEN_1\
        );

    \I__1136\ : IoInMux
    port map (
            O => \N__5529\,
            I => \N__5525\
        );

    \I__1135\ : CascadeMux
    port map (
            O => \N__5528\,
            I => \N__5520\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__5525\,
            I => \N__5517\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__5524\,
            I => \N__5514\
        );

    \I__1132\ : InMux
    port map (
            O => \N__5523\,
            I => \N__5511\
        );

    \I__1131\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5508\
        );

    \I__1130\ : IoSpan4Mux
    port map (
            O => \N__5517\,
            I => \N__5504\
        );

    \I__1129\ : InMux
    port map (
            O => \N__5514\,
            I => \N__5501\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__5511\,
            I => \N__5496\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__5508\,
            I => \N__5496\
        );

    \I__1126\ : CascadeMux
    port map (
            O => \N__5507\,
            I => \N__5491\
        );

    \I__1125\ : Span4Mux_s0_v
    port map (
            O => \N__5504\,
            I => \N__5487\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__5501\,
            I => \N__5482\
        );

    \I__1123\ : Span4Mux_v
    port map (
            O => \N__5496\,
            I => \N__5482\
        );

    \I__1122\ : InMux
    port map (
            O => \N__5495\,
            I => \N__5477\
        );

    \I__1121\ : InMux
    port map (
            O => \N__5494\,
            I => \N__5477\
        );

    \I__1120\ : InMux
    port map (
            O => \N__5491\,
            I => \N__5474\
        );

    \I__1119\ : InMux
    port map (
            O => \N__5490\,
            I => \N__5471\
        );

    \I__1118\ : Sp12to4
    port map (
            O => \N__5487\,
            I => \N__5468\
        );

    \I__1117\ : Sp12to4
    port map (
            O => \N__5482\,
            I => \N__5465\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__5477\,
            I => \N__5462\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__5474\,
            I => \N__5457\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__5471\,
            I => \N__5457\
        );

    \I__1113\ : Span12Mux_v
    port map (
            O => \N__5468\,
            I => \N__5450\
        );

    \I__1112\ : Span12Mux_h
    port map (
            O => \N__5465\,
            I => \N__5450\
        );

    \I__1111\ : Sp12to4
    port map (
            O => \N__5462\,
            I => \N__5450\
        );

    \I__1110\ : Sp12to4
    port map (
            O => \N__5457\,
            I => \N__5447\
        );

    \I__1109\ : Span12Mux_v
    port map (
            O => \N__5450\,
            I => \N__5444\
        );

    \I__1108\ : Span12Mux_v
    port map (
            O => \N__5447\,
            I => \N__5441\
        );

    \I__1107\ : Odrv12
    port map (
            O => \N__5444\,
            I => \CLK40_IN_c\
        );

    \I__1106\ : Odrv12
    port map (
            O => \N__5441\,
            I => \CLK40_IN_c\
        );

    \I__1105\ : InMux
    port map (
            O => \N__5436\,
            I => \N__5427\
        );

    \I__1104\ : InMux
    port map (
            O => \N__5435\,
            I => \N__5418\
        );

    \I__1103\ : InMux
    port map (
            O => \N__5434\,
            I => \N__5418\
        );

    \I__1102\ : InMux
    port map (
            O => \N__5433\,
            I => \N__5418\
        );

    \I__1101\ : InMux
    port map (
            O => \N__5432\,
            I => \N__5418\
        );

    \I__1100\ : InMux
    port map (
            O => \N__5431\,
            I => \N__5415\
        );

    \I__1099\ : InMux
    port map (
            O => \N__5430\,
            I => \N__5412\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__5427\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__5418\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__5415\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__5412\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5403\,
            I => \N__5397\
        );

    \I__1093\ : InMux
    port map (
            O => \N__5402\,
            I => \N__5397\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__5397\,
            I => \U409_TRANSFER_ACK.N_28_4\
        );

    \I__1091\ : InMux
    port map (
            O => \N__5394\,
            I => \N__5389\
        );

    \I__1090\ : InMux
    port map (
            O => \N__5393\,
            I => \N__5384\
        );

    \I__1089\ : InMux
    port map (
            O => \N__5392\,
            I => \N__5384\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__5389\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__5384\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__1086\ : InMux
    port map (
            O => \N__5379\,
            I => \N__5376\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__5376\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__1084\ : CEMux
    port map (
            O => \N__5373\,
            I => \N__5370\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__5370\,
            I => \N__5367\
        );

    \I__1082\ : Odrv12
    port map (
            O => \N__5367\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1_0\
        );

    \I__1081\ : SRMux
    port map (
            O => \N__5364\,
            I => \N__5359\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5363\,
            I => \N__5355\
        );

    \I__1079\ : SRMux
    port map (
            O => \N__5362\,
            I => \N__5352\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__5359\,
            I => \N__5348\
        );

    \I__1077\ : SRMux
    port map (
            O => \N__5358\,
            I => \N__5345\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__5355\,
            I => \N__5340\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__5352\,
            I => \N__5340\
        );

    \I__1074\ : SRMux
    port map (
            O => \N__5351\,
            I => \N__5337\
        );

    \I__1073\ : Span4Mux_v
    port map (
            O => \N__5348\,
            I => \N__5332\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__5345\,
            I => \N__5332\
        );

    \I__1071\ : Span4Mux_v
    port map (
            O => \N__5340\,
            I => \N__5327\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__5337\,
            I => \N__5327\
        );

    \I__1069\ : Odrv4
    port map (
            O => \N__5332\,
            I => \RESETn_c_i\
        );

    \I__1068\ : Odrv4
    port map (
            O => \N__5327\,
            I => \RESETn_c_i\
        );

    \I__1067\ : CascadeMux
    port map (
            O => \N__5322\,
            I => \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\
        );

    \I__1066\ : IoInMux
    port map (
            O => \N__5319\,
            I => \N__5316\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__5316\,
            I => \N__5313\
        );

    \I__1064\ : Span12Mux_s3_v
    port map (
            O => \N__5313\,
            I => \N__5310\
        );

    \I__1063\ : Span12Mux_v
    port map (
            O => \N__5310\,
            I => \N__5305\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5309\,
            I => \N__5300\
        );

    \I__1061\ : InMux
    port map (
            O => \N__5308\,
            I => \N__5300\
        );

    \I__1060\ : Odrv12
    port map (
            O => \N__5305\,
            I => \TACK_OUTn\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__5300\,
            I => \TACK_OUTn\
        );

    \I__1058\ : CascadeMux
    port map (
            O => \N__5295\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_cascade_\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5292\,
            I => \N__5288\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5291\,
            I => \N__5285\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__5288\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__5285\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1053\ : CascadeMux
    port map (
            O => \N__5280\,
            I => \N__5276\
        );

    \I__1052\ : InMux
    port map (
            O => \N__5279\,
            I => \N__5273\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5276\,
            I => \N__5270\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__5273\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__5270\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1048\ : InMux
    port map (
            O => \N__5265\,
            I => \N__5261\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5264\,
            I => \N__5258\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__5261\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__5258\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1044\ : IoInMux
    port map (
            O => \N__5253\,
            I => \N__5250\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__5250\,
            I => \N__5247\
        );

    \I__1042\ : Span4Mux_s2_v
    port map (
            O => \N__5247\,
            I => \N__5244\
        );

    \I__1041\ : Span4Mux_v
    port map (
            O => \N__5244\,
            I => \N__5241\
        );

    \I__1040\ : Odrv4
    port map (
            O => \N__5241\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__5238\,
            I => \N__5234\
        );

    \I__1038\ : CascadeMux
    port map (
            O => \N__5237\,
            I => \N__5231\
        );

    \I__1037\ : InMux
    port map (
            O => \N__5234\,
            I => \N__5228\
        );

    \I__1036\ : InMux
    port map (
            O => \N__5231\,
            I => \N__5225\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__5228\,
            I => \N__5220\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__5225\,
            I => \N__5220\
        );

    \I__1033\ : Span4Mux_v
    port map (
            O => \N__5220\,
            I => \N__5217\
        );

    \I__1032\ : Span4Mux_h
    port map (
            O => \N__5217\,
            I => \N__5214\
        );

    \I__1031\ : Odrv4
    port map (
            O => \N__5214\,
            I => \U409_TRANSFER_ACK.N_18\
        );

    \I__1030\ : InMux
    port map (
            O => \N__5211\,
            I => \N__5208\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__5208\,
            I => \U409_TRANSFER_ACK.N_24\
        );

    \I__1028\ : InMux
    port map (
            O => \N__5205\,
            I => \N__5202\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__5202\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a5_0\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5199\,
            I => \N__5196\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__5196\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\
        );

    \I__1024\ : IoInMux
    port map (
            O => \N__5193\,
            I => \N__5190\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__5190\,
            I => \N__5187\
        );

    \I__1022\ : Span4Mux_s2_v
    port map (
            O => \N__5187\,
            I => \N__5184\
        );

    \I__1021\ : Span4Mux_h
    port map (
            O => \N__5184\,
            I => \N__5181\
        );

    \I__1020\ : Span4Mux_v
    port map (
            O => \N__5181\,
            I => \N__5177\
        );

    \I__1019\ : CascadeMux
    port map (
            O => \N__5180\,
            I => \N__5174\
        );

    \I__1018\ : Sp12to4
    port map (
            O => \N__5177\,
            I => \N__5171\
        );

    \I__1017\ : InMux
    port map (
            O => \N__5174\,
            I => \N__5168\
        );

    \I__1016\ : Odrv12
    port map (
            O => \N__5171\,
            I => \ROMENn_c\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__5168\,
            I => \ROMENn_c\
        );

    \I__1014\ : InMux
    port map (
            O => \N__5163\,
            I => \N__5160\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__5160\,
            I => \N__5157\
        );

    \I__1012\ : Span4Mux_v
    port map (
            O => \N__5157\,
            I => \N__5152\
        );

    \I__1011\ : InMux
    port map (
            O => \N__5156\,
            I => \N__5149\
        );

    \I__1010\ : InMux
    port map (
            O => \N__5155\,
            I => \N__5146\
        );

    \I__1009\ : Odrv4
    port map (
            O => \N__5152\,
            I => \U409_CIA.VMAZ0\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__5149\,
            I => \U409_CIA.VMAZ0\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__5146\,
            I => \U409_CIA.VMAZ0\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5139\,
            I => \N__5133\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5138\,
            I => \N__5126\
        );

    \I__1004\ : InMux
    port map (
            O => \N__5137\,
            I => \N__5126\
        );

    \I__1003\ : InMux
    port map (
            O => \N__5136\,
            I => \N__5126\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__5133\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__5126\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__1000\ : InMux
    port map (
            O => \N__5121\,
            I => \N__5115\
        );

    \I__999\ : InMux
    port map (
            O => \N__5120\,
            I => \N__5112\
        );

    \I__998\ : InMux
    port map (
            O => \N__5119\,
            I => \N__5107\
        );

    \I__997\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5107\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5115\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__5112\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5107\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__993\ : InMux
    port map (
            O => \N__5100\,
            I => \N__5095\
        );

    \I__992\ : InMux
    port map (
            O => \N__5099\,
            I => \N__5090\
        );

    \I__991\ : InMux
    port map (
            O => \N__5098\,
            I => \N__5090\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__5095\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__5090\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__988\ : CascadeMux
    port map (
            O => \N__5085\,
            I => \N__5082\
        );

    \I__987\ : InMux
    port map (
            O => \N__5082\,
            I => \N__5079\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__5079\,
            I => \U409_TRANSFER_ACK.ROM_TACK_EN_e_1\
        );

    \I__985\ : InMux
    port map (
            O => \N__5076\,
            I => \N__5072\
        );

    \I__984\ : InMux
    port map (
            O => \N__5075\,
            I => \N__5069\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__5072\,
            I => \N__5062\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__5069\,
            I => \N__5062\
        );

    \I__981\ : InMux
    port map (
            O => \N__5068\,
            I => \N__5057\
        );

    \I__980\ : InMux
    port map (
            O => \N__5067\,
            I => \N__5057\
        );

    \I__979\ : Odrv4
    port map (
            O => \N__5062\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__5057\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__977\ : InMux
    port map (
            O => \N__5052\,
            I => \N__5045\
        );

    \I__976\ : InMux
    port map (
            O => \N__5051\,
            I => \N__5042\
        );

    \I__975\ : InMux
    port map (
            O => \N__5050\,
            I => \N__5039\
        );

    \I__974\ : InMux
    port map (
            O => \N__5049\,
            I => \N__5034\
        );

    \I__973\ : InMux
    port map (
            O => \N__5048\,
            I => \N__5034\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__5045\,
            I => \N__5029\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__5042\,
            I => \N__5029\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__5039\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__5034\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__968\ : Odrv4
    port map (
            O => \N__5029\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__967\ : CascadeMux
    port map (
            O => \N__5022\,
            I => \N__5019\
        );

    \I__966\ : InMux
    port map (
            O => \N__5019\,
            I => \N__5016\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__5016\,
            I => \U409_TRANSFER_ACK.N_138\
        );

    \I__964\ : InMux
    port map (
            O => \N__5013\,
            I => \N__5007\
        );

    \I__963\ : InMux
    port map (
            O => \N__5012\,
            I => \N__5007\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__5007\,
            I => \N__5004\
        );

    \I__961\ : Span4Mux_v
    port map (
            O => \N__5004\,
            I => \N__5001\
        );

    \I__960\ : Sp12to4
    port map (
            O => \N__5001\,
            I => \N__4998\
        );

    \I__959\ : Odrv12
    port map (
            O => \N__4998\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_0\
        );

    \I__958\ : SRMux
    port map (
            O => \N__4995\,
            I => \N__4991\
        );

    \I__957\ : SRMux
    port map (
            O => \N__4994\,
            I => \N__4988\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__4991\,
            I => \N__4982\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4988\,
            I => \N__4982\
        );

    \I__954\ : SRMux
    port map (
            O => \N__4987\,
            I => \N__4979\
        );

    \I__953\ : Span4Mux_v
    port map (
            O => \N__4982\,
            I => \N__4976\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__4979\,
            I => \N__4973\
        );

    \I__951\ : Sp12to4
    port map (
            O => \N__4976\,
            I => \N__4970\
        );

    \I__950\ : Sp12to4
    port map (
            O => \N__4973\,
            I => \N__4967\
        );

    \I__949\ : Odrv12
    port map (
            O => \N__4970\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__948\ : Odrv12
    port map (
            O => \N__4967\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__947\ : CascadeMux
    port map (
            O => \N__4962\,
            I => \U409_TRANSFER_ACK.m8_ns_1_cascade_\
        );

    \I__946\ : CascadeMux
    port map (
            O => \N__4959\,
            I => \U409_TRANSFER_ACK.i6_mux_0_cascade_\
        );

    \I__945\ : InMux
    port map (
            O => \N__4956\,
            I => \N__4953\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4953\,
            I => \U409_TRANSFER_ACK.N_9\
        );

    \I__943\ : InMux
    port map (
            O => \N__4950\,
            I => \N__4947\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__4947\,
            I => \U409_TRANSFER_ACK.N_4\
        );

    \I__941\ : CascadeMux
    port map (
            O => \N__4944\,
            I => \U409_TRANSFER_ACK.N_4_cascade_\
        );

    \I__940\ : InMux
    port map (
            O => \N__4941\,
            I => \N__4938\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__4938\,
            I => \U409_TRANSFER_ACK.N_5\
        );

    \I__938\ : CascadeMux
    port map (
            O => \N__4935\,
            I => \N__4932\
        );

    \I__937\ : InMux
    port map (
            O => \N__4932\,
            I => \N__4923\
        );

    \I__936\ : InMux
    port map (
            O => \N__4931\,
            I => \N__4923\
        );

    \I__935\ : InMux
    port map (
            O => \N__4930\,
            I => \N__4923\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__4923\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__933\ : IoInMux
    port map (
            O => \N__4920\,
            I => \N__4917\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4917\,
            I => \N__4914\
        );

    \I__931\ : IoSpan4Mux
    port map (
            O => \N__4914\,
            I => \N__4911\
        );

    \I__930\ : Sp12to4
    port map (
            O => \N__4911\,
            I => \N__4908\
        );

    \I__929\ : Span12Mux_s6_v
    port map (
            O => \N__4908\,
            I => \N__4905\
        );

    \I__928\ : Span12Mux_v
    port map (
            O => \N__4905\,
            I => \N__4900\
        );

    \I__927\ : InMux
    port map (
            O => \N__4904\,
            I => \N__4897\
        );

    \I__926\ : InMux
    port map (
            O => \N__4903\,
            I => \N__4894\
        );

    \I__925\ : Odrv12
    port map (
            O => \N__4900\,
            I => \CLK_CIA_c\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__4897\,
            I => \CLK_CIA_c\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__4894\,
            I => \CLK_CIA_c\
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__4887\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\
        );

    \I__921\ : InMux
    port map (
            O => \N__4884\,
            I => \N__4881\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4881\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5\
        );

    \I__919\ : InMux
    port map (
            O => \N__4878\,
            I => \N__4873\
        );

    \I__918\ : InMux
    port map (
            O => \N__4877\,
            I => \N__4868\
        );

    \I__917\ : InMux
    port map (
            O => \N__4876\,
            I => \N__4868\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4873\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__4868\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__4863\,
            I => \N__4858\
        );

    \I__913\ : InMux
    port map (
            O => \N__4862\,
            I => \N__4852\
        );

    \I__912\ : InMux
    port map (
            O => \N__4861\,
            I => \N__4852\
        );

    \I__911\ : InMux
    port map (
            O => \N__4858\,
            I => \N__4847\
        );

    \I__910\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4847\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__4852\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4847\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__907\ : CascadeMux
    port map (
            O => \N__4842\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_6_cascade_\
        );

    \I__906\ : InMux
    port map (
            O => \N__4839\,
            I => \N__4836\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__4836\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1\
        );

    \I__904\ : InMux
    port map (
            O => \N__4833\,
            I => \N__4830\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4830\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\
        );

    \I__902\ : CascadeMux
    port map (
            O => \N__4827\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_\
        );

    \I__901\ : InMux
    port map (
            O => \N__4824\,
            I => \N__4817\
        );

    \I__900\ : InMux
    port map (
            O => \N__4823\,
            I => \N__4817\
        );

    \I__899\ : InMux
    port map (
            O => \N__4822\,
            I => \N__4813\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__4817\,
            I => \N__4810\
        );

    \I__897\ : InMux
    port map (
            O => \N__4816\,
            I => \N__4807\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__4813\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__895\ : Odrv4
    port map (
            O => \N__4810\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__4807\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__893\ : InMux
    port map (
            O => \N__4800\,
            I => \N__4793\
        );

    \I__892\ : InMux
    port map (
            O => \N__4799\,
            I => \N__4793\
        );

    \I__891\ : InMux
    port map (
            O => \N__4798\,
            I => \N__4790\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__4793\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__4790\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\
        );

    \I__888\ : InMux
    port map (
            O => \N__4785\,
            I => \N__4775\
        );

    \I__887\ : InMux
    port map (
            O => \N__4784\,
            I => \N__4775\
        );

    \I__886\ : InMux
    port map (
            O => \N__4783\,
            I => \N__4772\
        );

    \I__885\ : InMux
    port map (
            O => \N__4782\,
            I => \N__4765\
        );

    \I__884\ : InMux
    port map (
            O => \N__4781\,
            I => \N__4765\
        );

    \I__883\ : InMux
    port map (
            O => \N__4780\,
            I => \N__4765\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__4775\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__4772\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4765\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__4758\,
            I => \N__4753\
        );

    \I__878\ : CascadeMux
    port map (
            O => \N__4757\,
            I => \N__4750\
        );

    \I__877\ : InMux
    port map (
            O => \N__4756\,
            I => \N__4746\
        );

    \I__876\ : InMux
    port map (
            O => \N__4753\,
            I => \N__4739\
        );

    \I__875\ : InMux
    port map (
            O => \N__4750\,
            I => \N__4739\
        );

    \I__874\ : InMux
    port map (
            O => \N__4749\,
            I => \N__4739\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__4746\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4739\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__871\ : InMux
    port map (
            O => \N__4734\,
            I => \N__4729\
        );

    \I__870\ : InMux
    port map (
            O => \N__4733\,
            I => \N__4726\
        );

    \I__869\ : InMux
    port map (
            O => \N__4732\,
            I => \N__4723\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4729\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4726\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__4723\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__865\ : InMux
    port map (
            O => \N__4716\,
            I => \N__4704\
        );

    \I__864\ : InMux
    port map (
            O => \N__4715\,
            I => \N__4704\
        );

    \I__863\ : InMux
    port map (
            O => \N__4714\,
            I => \N__4704\
        );

    \I__862\ : InMux
    port map (
            O => \N__4713\,
            I => \N__4697\
        );

    \I__861\ : InMux
    port map (
            O => \N__4712\,
            I => \N__4697\
        );

    \I__860\ : InMux
    port map (
            O => \N__4711\,
            I => \N__4697\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__4704\,
            I => \N__4694\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__4697\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__857\ : Odrv4
    port map (
            O => \N__4694\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__4689\,
            I => \N__4683\
        );

    \I__855\ : CascadeMux
    port map (
            O => \N__4688\,
            I => \N__4679\
        );

    \I__854\ : CascadeMux
    port map (
            O => \N__4687\,
            I => \N__4676\
        );

    \I__853\ : InMux
    port map (
            O => \N__4686\,
            I => \N__4668\
        );

    \I__852\ : InMux
    port map (
            O => \N__4683\,
            I => \N__4668\
        );

    \I__851\ : InMux
    port map (
            O => \N__4682\,
            I => \N__4668\
        );

    \I__850\ : InMux
    port map (
            O => \N__4679\,
            I => \N__4661\
        );

    \I__849\ : InMux
    port map (
            O => \N__4676\,
            I => \N__4661\
        );

    \I__848\ : InMux
    port map (
            O => \N__4675\,
            I => \N__4661\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4668\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4661\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__845\ : InMux
    port map (
            O => \N__4656\,
            I => \N__4647\
        );

    \I__844\ : InMux
    port map (
            O => \N__4655\,
            I => \N__4647\
        );

    \I__843\ : InMux
    port map (
            O => \N__4654\,
            I => \N__4640\
        );

    \I__842\ : InMux
    port map (
            O => \N__4653\,
            I => \N__4640\
        );

    \I__841\ : InMux
    port map (
            O => \N__4652\,
            I => \N__4640\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__4647\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4640\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__838\ : InMux
    port map (
            O => \N__4635\,
            I => \N__4628\
        );

    \I__837\ : InMux
    port map (
            O => \N__4634\,
            I => \N__4621\
        );

    \I__836\ : InMux
    port map (
            O => \N__4633\,
            I => \N__4621\
        );

    \I__835\ : InMux
    port map (
            O => \N__4632\,
            I => \N__4621\
        );

    \I__834\ : InMux
    port map (
            O => \N__4631\,
            I => \N__4618\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__4628\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4621\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4618\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__830\ : CascadeMux
    port map (
            O => \N__4611\,
            I => \N__4606\
        );

    \I__829\ : InMux
    port map (
            O => \N__4610\,
            I => \N__4601\
        );

    \I__828\ : InMux
    port map (
            O => \N__4609\,
            I => \N__4594\
        );

    \I__827\ : InMux
    port map (
            O => \N__4606\,
            I => \N__4594\
        );

    \I__826\ : InMux
    port map (
            O => \N__4605\,
            I => \N__4594\
        );

    \I__825\ : InMux
    port map (
            O => \N__4604\,
            I => \N__4591\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__4601\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__4594\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__4591\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__821\ : ClkMux
    port map (
            O => \N__4584\,
            I => \N__4572\
        );

    \I__820\ : ClkMux
    port map (
            O => \N__4583\,
            I => \N__4572\
        );

    \I__819\ : ClkMux
    port map (
            O => \N__4582\,
            I => \N__4572\
        );

    \I__818\ : ClkMux
    port map (
            O => \N__4581\,
            I => \N__4572\
        );

    \I__817\ : GlobalMux
    port map (
            O => \N__4572\,
            I => \N__4569\
        );

    \I__816\ : gio2CtrlBuf
    port map (
            O => \N__4569\,
            I => \CLK28_IN_c_g\
        );

    \I__815\ : InMux
    port map (
            O => \N__4566\,
            I => \N__4560\
        );

    \I__814\ : InMux
    port map (
            O => \N__4565\,
            I => \N__4557\
        );

    \I__813\ : InMux
    port map (
            O => \N__4564\,
            I => \N__4554\
        );

    \I__812\ : InMux
    port map (
            O => \N__4563\,
            I => \N__4551\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__4560\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__4557\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__4554\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4551\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__807\ : CascadeMux
    port map (
            O => \N__4542\,
            I => \N__4534\
        );

    \I__806\ : InMux
    port map (
            O => \N__4541\,
            I => \N__4531\
        );

    \I__805\ : InMux
    port map (
            O => \N__4540\,
            I => \N__4526\
        );

    \I__804\ : InMux
    port map (
            O => \N__4539\,
            I => \N__4526\
        );

    \I__803\ : InMux
    port map (
            O => \N__4538\,
            I => \N__4523\
        );

    \I__802\ : InMux
    port map (
            O => \N__4537\,
            I => \N__4520\
        );

    \I__801\ : InMux
    port map (
            O => \N__4534\,
            I => \N__4517\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4531\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4526\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4523\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__4520\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__4517\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__4506\,
            I => \N__4500\
        );

    \I__794\ : CascadeMux
    port map (
            O => \N__4505\,
            I => \N__4497\
        );

    \I__793\ : InMux
    port map (
            O => \N__4504\,
            I => \N__4494\
        );

    \I__792\ : InMux
    port map (
            O => \N__4503\,
            I => \N__4491\
        );

    \I__791\ : InMux
    port map (
            O => \N__4500\,
            I => \N__4488\
        );

    \I__790\ : InMux
    port map (
            O => \N__4497\,
            I => \N__4485\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__4494\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__4491\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__4488\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__4485\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__785\ : InMux
    port map (
            O => \N__4476\,
            I => \N__4468\
        );

    \I__784\ : InMux
    port map (
            O => \N__4475\,
            I => \N__4468\
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__4474\,
            I => \N__4465\
        );

    \I__782\ : InMux
    port map (
            O => \N__4473\,
            I => \N__4460\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__4468\,
            I => \N__4457\
        );

    \I__780\ : InMux
    port map (
            O => \N__4465\,
            I => \N__4454\
        );

    \I__779\ : InMux
    port map (
            O => \N__4464\,
            I => \N__4451\
        );

    \I__778\ : InMux
    port map (
            O => \N__4463\,
            I => \N__4448\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__4460\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__776\ : Odrv12
    port map (
            O => \N__4457\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__4454\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__4451\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__4448\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__772\ : InMux
    port map (
            O => \N__4437\,
            I => \N__4434\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__4434\,
            I => \N__4431\
        );

    \I__770\ : Odrv4
    port map (
            O => \N__4431\,
            I => \U409_CIA.CLK_CIA6_3\
        );

    \I__769\ : CascadeMux
    port map (
            O => \N__4428\,
            I => \N__4425\
        );

    \I__768\ : InMux
    port map (
            O => \N__4425\,
            I => \N__4421\
        );

    \I__767\ : CascadeMux
    port map (
            O => \N__4424\,
            I => \N__4417\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__4421\,
            I => \N__4412\
        );

    \I__765\ : InMux
    port map (
            O => \N__4420\,
            I => \N__4407\
        );

    \I__764\ : InMux
    port map (
            O => \N__4417\,
            I => \N__4407\
        );

    \I__763\ : InMux
    port map (
            O => \N__4416\,
            I => \N__4404\
        );

    \I__762\ : InMux
    port map (
            O => \N__4415\,
            I => \N__4401\
        );

    \I__761\ : Odrv4
    port map (
            O => \N__4412\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__4407\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__4404\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__4401\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__757\ : InMux
    port map (
            O => \N__4392\,
            I => \N__4389\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__4389\,
            I => \U409_CIA.un1_CIA_CLK_COUNT_2_1\
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__4386\,
            I => \U409_CIA.CLK_CIA6_3_cascade_\
        );

    \I__754\ : InMux
    port map (
            O => \N__4383\,
            I => \N__4374\
        );

    \I__753\ : InMux
    port map (
            O => \N__4382\,
            I => \N__4374\
        );

    \I__752\ : InMux
    port map (
            O => \N__4381\,
            I => \N__4371\
        );

    \I__751\ : InMux
    port map (
            O => \N__4380\,
            I => \N__4368\
        );

    \I__750\ : InMux
    port map (
            O => \N__4379\,
            I => \N__4365\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__4374\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__4371\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__4368\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__4365\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__745\ : InMux
    port map (
            O => \N__4356\,
            I => \N__4353\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__4353\,
            I => \U409_CIA.CLK_CIA_RNOZ0Z_1\
        );

    \I__743\ : InMux
    port map (
            O => \N__4350\,
            I => \N__4345\
        );

    \I__742\ : InMux
    port map (
            O => \N__4349\,
            I => \N__4342\
        );

    \I__741\ : InMux
    port map (
            O => \N__4348\,
            I => \N__4339\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__4345\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__4342\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__4339\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__737\ : CascadeMux
    port map (
            O => \N__4332\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\
        );

    \I__736\ : InMux
    port map (
            O => \N__4329\,
            I => \N__4326\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__4326\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\
        );

    \I__734\ : InMux
    port map (
            O => \N__4323\,
            I => \N__4320\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__4320\,
            I => \N__4317\
        );

    \I__732\ : Span12Mux_h
    port map (
            O => \N__4317\,
            I => \N__4314\
        );

    \I__731\ : Odrv12
    port map (
            O => \N__4314\,
            I => \A_c_12\
        );

    \I__730\ : IoInMux
    port map (
            O => \N__4311\,
            I => \N__4308\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__4308\,
            I => \N__4305\
        );

    \I__728\ : Span4Mux_s0_h
    port map (
            O => \N__4305\,
            I => \N__4302\
        );

    \I__727\ : Sp12to4
    port map (
            O => \N__4302\,
            I => \N__4299\
        );

    \I__726\ : Span12Mux_s10_v
    port map (
            O => \N__4299\,
            I => \N__4296\
        );

    \I__725\ : Span12Mux_h
    port map (
            O => \N__4296\,
            I => \N__4293\
        );

    \I__724\ : Odrv12
    port map (
            O => \N__4293\,
            I => \U409_ADDRESS_DECODE_un1_CIACS0n_i\
        );

    \I__723\ : InMux
    port map (
            O => \N__4290\,
            I => \N__4287\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4287\,
            I => \N__4283\
        );

    \I__721\ : InMux
    port map (
            O => \N__4286\,
            I => \N__4280\
        );

    \I__720\ : Odrv4
    port map (
            O => \N__4283\,
            I => \CIA_ENABLE\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__4280\,
            I => \CIA_ENABLE\
        );

    \I__718\ : InMux
    port map (
            O => \N__4275\,
            I => \N__4271\
        );

    \I__717\ : InMux
    port map (
            O => \N__4274\,
            I => \N__4268\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__4271\,
            I => \U409_CIA.CLK_CIA6_0\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__4268\,
            I => \U409_CIA.CLK_CIA6_0\
        );

    \I__714\ : CascadeMux
    port map (
            O => \N__4263\,
            I => \U409_CIA.CLK_CIA6_cascade_\
        );

    \I__713\ : InMux
    port map (
            O => \N__4260\,
            I => \N__4257\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__4257\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\
        );

    \I__711\ : InMux
    port map (
            O => \N__4254\,
            I => \N__4251\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__4251\,
            I => \U409_CIA.CIA_CLK_COUNT11_2_0\
        );

    \I__709\ : CascadeMux
    port map (
            O => \N__4248\,
            I => \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_\
        );

    \I__708\ : InMux
    port map (
            O => \N__4245\,
            I => \N__4242\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__4242\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO\
        );

    \I__706\ : CascadeMux
    port map (
            O => \N__4239\,
            I => \N__4235\
        );

    \I__705\ : InMux
    port map (
            O => \N__4238\,
            I => \N__4230\
        );

    \I__704\ : InMux
    port map (
            O => \N__4235\,
            I => \N__4230\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__4230\,
            I => \U409_CIA.CIA_CLK_COUNT11_3\
        );

    \I__702\ : InMux
    port map (
            O => \N__4227\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\
        );

    \I__701\ : CascadeMux
    port map (
            O => \N__4224\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_cascade_\
        );

    \I__700\ : CascadeMux
    port map (
            O => \N__4221\,
            I => \N__4218\
        );

    \I__699\ : InMux
    port map (
            O => \N__4218\,
            I => \N__4212\
        );

    \I__698\ : InMux
    port map (
            O => \N__4217\,
            I => \N__4212\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__4212\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\
        );

    \I__696\ : InMux
    port map (
            O => \N__4209\,
            I => \N__4204\
        );

    \I__695\ : InMux
    port map (
            O => \N__4208\,
            I => \N__4201\
        );

    \I__694\ : InMux
    port map (
            O => \N__4207\,
            I => \N__4198\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__4204\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__4201\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__4198\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn\
        );

    \I__690\ : InMux
    port map (
            O => \N__4191\,
            I => \N__4188\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__4188\,
            I => \N__4185\
        );

    \I__688\ : Odrv4
    port map (
            O => \N__4185\,
            I => \U409_ADDRESS_DECODE_un1_RAMSPACEn\
        );

    \I__687\ : InMux
    port map (
            O => \N__4182\,
            I => \N__4179\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__4179\,
            I => \N__4176\
        );

    \I__685\ : Span12Mux_h
    port map (
            O => \N__4176\,
            I => \N__4173\
        );

    \I__684\ : Span12Mux_h
    port map (
            O => \N__4173\,
            I => \N__4170\
        );

    \I__683\ : Span12Mux_v
    port map (
            O => \N__4170\,
            I => \N__4167\
        );

    \I__682\ : Odrv12
    port map (
            O => \N__4167\,
            I => \TACKn_in\
        );

    \I__681\ : InMux
    port map (
            O => \N__4164\,
            I => \N__4161\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__4161\,
            I => \N__4158\
        );

    \I__679\ : Span12Mux_v
    port map (
            O => \N__4158\,
            I => \N__4155\
        );

    \I__678\ : Span12Mux_h
    port map (
            O => \N__4155\,
            I => \N__4152\
        );

    \I__677\ : Odrv12
    port map (
            O => \N__4152\,
            I => \A_c_13\
        );

    \I__676\ : IoInMux
    port map (
            O => \N__4149\,
            I => \N__4146\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__4146\,
            I => \N__4143\
        );

    \I__674\ : Span4Mux_s0_h
    port map (
            O => \N__4143\,
            I => \N__4140\
        );

    \I__673\ : Sp12to4
    port map (
            O => \N__4140\,
            I => \N__4137\
        );

    \I__672\ : Span12Mux_s9_v
    port map (
            O => \N__4137\,
            I => \N__4134\
        );

    \I__671\ : Span12Mux_h
    port map (
            O => \N__4134\,
            I => \N__4131\
        );

    \I__670\ : Odrv12
    port map (
            O => \N__4131\,
            I => \U409_ADDRESS_DECODE_un1_CIACS1n_i\
        );

    \I__669\ : InMux
    port map (
            O => \N__4128\,
            I => \N__4125\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__4125\,
            I => \N__4121\
        );

    \I__667\ : InMux
    port map (
            O => \N__4124\,
            I => \N__4118\
        );

    \I__666\ : Span12Mux_h
    port map (
            O => \N__4121\,
            I => \N__4115\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__4118\,
            I => \N__4112\
        );

    \I__664\ : Odrv12
    port map (
            O => \N__4115\,
            I => \CIA_SPACE\
        );

    \I__663\ : Odrv4
    port map (
            O => \N__4112\,
            I => \CIA_SPACE\
        );

    \I__662\ : CascadeMux
    port map (
            O => \N__4107\,
            I => \U409_CIA.VMA_RNOZ0Z_0_cascade_\
        );

    \I__661\ : InMux
    port map (
            O => \N__4104\,
            I => \N__4101\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__4101\,
            I => \U409_CIA.un1_CIA_CLK_COUNT_3_1\
        );

    \I__659\ : InMux
    port map (
            O => \N__4098\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\
        );

    \I__658\ : InMux
    port map (
            O => \N__4095\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\
        );

    \I__657\ : InMux
    port map (
            O => \N__4092\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\
        );

    \I__656\ : InMux
    port map (
            O => \N__4089\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\
        );

    \I__655\ : InMux
    port map (
            O => \N__4086\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\
        );

    \I__654\ : InMux
    port map (
            O => \N__4083\,
            I => \N__4080\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__4080\,
            I => \N__4076\
        );

    \I__652\ : InMux
    port map (
            O => \N__4079\,
            I => \N__4073\
        );

    \I__651\ : Span4Mux_v
    port map (
            O => \N__4076\,
            I => \N__4070\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__4073\,
            I => \N__4067\
        );

    \I__649\ : Sp12to4
    port map (
            O => \N__4070\,
            I => \N__4064\
        );

    \I__648\ : Sp12to4
    port map (
            O => \N__4067\,
            I => \N__4061\
        );

    \I__647\ : Span12Mux_h
    port map (
            O => \N__4064\,
            I => \N__4058\
        );

    \I__646\ : Span12Mux_v
    port map (
            O => \N__4061\,
            I => \N__4055\
        );

    \I__645\ : Span12Mux_v
    port map (
            O => \N__4058\,
            I => \N__4050\
        );

    \I__644\ : Span12Mux_h
    port map (
            O => \N__4055\,
            I => \N__4050\
        );

    \I__643\ : Odrv12
    port map (
            O => \N__4050\,
            I => \OVL_c\
        );

    \I__642\ : CascadeMux
    port map (
            O => \N__4047\,
            I => \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0_cascade_\
        );

    \I__641\ : IoInMux
    port map (
            O => \N__4044\,
            I => \N__4041\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__4041\,
            I => \N__4038\
        );

    \I__639\ : Span4Mux_s3_v
    port map (
            O => \N__4038\,
            I => \N__4035\
        );

    \I__638\ : Sp12to4
    port map (
            O => \N__4035\,
            I => \N__4032\
        );

    \I__637\ : Span12Mux_h
    port map (
            O => \N__4032\,
            I => \N__4029\
        );

    \I__636\ : Span12Mux_v
    port map (
            O => \N__4029\,
            I => \N__4026\
        );

    \I__635\ : Odrv12
    port map (
            O => \N__4026\,
            I => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\
        );

    \I__634\ : InMux
    port map (
            O => \N__4023\,
            I => \N__4020\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__4020\,
            I => \N__4016\
        );

    \I__632\ : InMux
    port map (
            O => \N__4019\,
            I => \N__4013\
        );

    \I__631\ : Span4Mux_v
    port map (
            O => \N__4016\,
            I => \N__4010\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4013\,
            I => \N__4007\
        );

    \I__629\ : Odrv4
    port map (
            O => \N__4010\,
            I => \U409_ADDRESS_DECODE_un1_RTC_ENn\
        );

    \I__628\ : Odrv4
    port map (
            O => \N__4007\,
            I => \U409_ADDRESS_DECODE_un1_RTC_ENn\
        );

    \I__627\ : IoInMux
    port map (
            O => \N__4002\,
            I => \N__3999\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__3999\,
            I => \N__3996\
        );

    \I__625\ : Span4Mux_s2_v
    port map (
            O => \N__3996\,
            I => \N__3993\
        );

    \I__624\ : Sp12to4
    port map (
            O => \N__3993\,
            I => \N__3990\
        );

    \I__623\ : Span12Mux_h
    port map (
            O => \N__3990\,
            I => \N__3987\
        );

    \I__622\ : Span12Mux_v
    port map (
            O => \N__3987\,
            I => \N__3984\
        );

    \I__621\ : Odrv12
    port map (
            O => \N__3984\,
            I => \PORTSIZE_0_i\
        );

    \I__620\ : InMux
    port map (
            O => \N__3981\,
            I => \N__3972\
        );

    \I__619\ : InMux
    port map (
            O => \N__3980\,
            I => \N__3965\
        );

    \I__618\ : InMux
    port map (
            O => \N__3979\,
            I => \N__3965\
        );

    \I__617\ : InMux
    port map (
            O => \N__3978\,
            I => \N__3965\
        );

    \I__616\ : InMux
    port map (
            O => \N__3977\,
            I => \N__3960\
        );

    \I__615\ : InMux
    port map (
            O => \N__3976\,
            I => \N__3955\
        );

    \I__614\ : InMux
    port map (
            O => \N__3975\,
            I => \N__3955\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__3972\,
            I => \N__3950\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__3965\,
            I => \N__3950\
        );

    \I__611\ : InMux
    port map (
            O => \N__3964\,
            I => \N__3947\
        );

    \I__610\ : InMux
    port map (
            O => \N__3963\,
            I => \N__3944\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__3960\,
            I => \N__3939\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__3955\,
            I => \N__3939\
        );

    \I__607\ : Span4Mux_h
    port map (
            O => \N__3950\,
            I => \N__3932\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3947\,
            I => \N__3932\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__3944\,
            I => \N__3932\
        );

    \I__604\ : Span4Mux_v
    port map (
            O => \N__3939\,
            I => \N__3929\
        );

    \I__603\ : Span4Mux_v
    port map (
            O => \N__3932\,
            I => \N__3926\
        );

    \I__602\ : Sp12to4
    port map (
            O => \N__3929\,
            I => \N__3921\
        );

    \I__601\ : Sp12to4
    port map (
            O => \N__3926\,
            I => \N__3921\
        );

    \I__600\ : Odrv12
    port map (
            O => \N__3921\,
            I => \A_c_23\
        );

    \I__599\ : InMux
    port map (
            O => \N__3918\,
            I => \N__3915\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3915\,
            I => \N__3912\
        );

    \I__597\ : Odrv4
    port map (
            O => \N__3912\,
            I => \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0\
        );

    \I__596\ : CascadeMux
    port map (
            O => \N__3909\,
            I => \N__3906\
        );

    \I__595\ : InMux
    port map (
            O => \N__3906\,
            I => \N__3903\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__3903\,
            I => \N__3895\
        );

    \I__593\ : InMux
    port map (
            O => \N__3902\,
            I => \N__3889\
        );

    \I__592\ : InMux
    port map (
            O => \N__3901\,
            I => \N__3889\
        );

    \I__591\ : InMux
    port map (
            O => \N__3900\,
            I => \N__3884\
        );

    \I__590\ : InMux
    port map (
            O => \N__3899\,
            I => \N__3884\
        );

    \I__589\ : InMux
    port map (
            O => \N__3898\,
            I => \N__3881\
        );

    \I__588\ : Span4Mux_v
    port map (
            O => \N__3895\,
            I => \N__3878\
        );

    \I__587\ : InMux
    port map (
            O => \N__3894\,
            I => \N__3872\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__3889\,
            I => \N__3865\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__3884\,
            I => \N__3865\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__3881\,
            I => \N__3865\
        );

    \I__583\ : Span4Mux_v
    port map (
            O => \N__3878\,
            I => \N__3862\
        );

    \I__582\ : InMux
    port map (
            O => \N__3877\,
            I => \N__3857\
        );

    \I__581\ : InMux
    port map (
            O => \N__3876\,
            I => \N__3857\
        );

    \I__580\ : InMux
    port map (
            O => \N__3875\,
            I => \N__3854\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__3872\,
            I => \N__3851\
        );

    \I__578\ : Span12Mux_h
    port map (
            O => \N__3865\,
            I => \N__3848\
        );

    \I__577\ : Span4Mux_v
    port map (
            O => \N__3862\,
            I => \N__3845\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__3857\,
            I => \N__3838\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__3854\,
            I => \N__3838\
        );

    \I__574\ : Sp12to4
    port map (
            O => \N__3851\,
            I => \N__3838\
        );

    \I__573\ : Span12Mux_v
    port map (
            O => \N__3848\,
            I => \N__3835\
        );

    \I__572\ : Sp12to4
    port map (
            O => \N__3845\,
            I => \N__3830\
        );

    \I__571\ : Span12Mux_v
    port map (
            O => \N__3838\,
            I => \N__3830\
        );

    \I__570\ : Odrv12
    port map (
            O => \N__3835\,
            I => \A_c_22\
        );

    \I__569\ : Odrv12
    port map (
            O => \N__3830\,
            I => \A_c_22\
        );

    \I__568\ : CascadeMux
    port map (
            O => \N__3825\,
            I => \N__3820\
        );

    \I__567\ : InMux
    port map (
            O => \N__3824\,
            I => \N__3813\
        );

    \I__566\ : InMux
    port map (
            O => \N__3823\,
            I => \N__3808\
        );

    \I__565\ : InMux
    port map (
            O => \N__3820\,
            I => \N__3808\
        );

    \I__564\ : InMux
    port map (
            O => \N__3819\,
            I => \N__3802\
        );

    \I__563\ : InMux
    port map (
            O => \N__3818\,
            I => \N__3799\
        );

    \I__562\ : InMux
    port map (
            O => \N__3817\,
            I => \N__3794\
        );

    \I__561\ : InMux
    port map (
            O => \N__3816\,
            I => \N__3794\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3813\,
            I => \N__3791\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__3808\,
            I => \N__3788\
        );

    \I__558\ : InMux
    port map (
            O => \N__3807\,
            I => \N__3783\
        );

    \I__557\ : InMux
    port map (
            O => \N__3806\,
            I => \N__3783\
        );

    \I__556\ : InMux
    port map (
            O => \N__3805\,
            I => \N__3780\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__3802\,
            I => \N__3773\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__3799\,
            I => \N__3773\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3794\,
            I => \N__3773\
        );

    \I__552\ : Span4Mux_h
    port map (
            O => \N__3791\,
            I => \N__3764\
        );

    \I__551\ : Span4Mux_h
    port map (
            O => \N__3788\,
            I => \N__3764\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__3783\,
            I => \N__3764\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3780\,
            I => \N__3764\
        );

    \I__548\ : Span4Mux_v
    port map (
            O => \N__3773\,
            I => \N__3761\
        );

    \I__547\ : Span4Mux_v
    port map (
            O => \N__3764\,
            I => \N__3758\
        );

    \I__546\ : Sp12to4
    port map (
            O => \N__3761\,
            I => \N__3753\
        );

    \I__545\ : Sp12to4
    port map (
            O => \N__3758\,
            I => \N__3753\
        );

    \I__544\ : Odrv12
    port map (
            O => \N__3753\,
            I => \A_c_21\
        );

    \I__543\ : CascadeMux
    port map (
            O => \N__3750\,
            I => \U409_ADDRESS_DECODE_un1_RAMSPACEn_cascade_\
        );

    \I__542\ : InMux
    port map (
            O => \N__3747\,
            I => \N__3744\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3744\,
            I => \U409_ADDRESS_DECODE_AUTOCONFIG_SPACE_5\
        );

    \I__540\ : InMux
    port map (
            O => \N__3741\,
            I => \N__3738\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3738\,
            I => \N__3735\
        );

    \I__538\ : Odrv4
    port map (
            O => \N__3735\,
            I => \U409_ADDRESS_DECODE_AUTOCONFIG_SPACE_7\
        );

    \I__537\ : CascadeMux
    port map (
            O => \N__3732\,
            I => \AGNUS_SPACE_0_cascade_\
        );

    \I__536\ : InMux
    port map (
            O => \N__3729\,
            I => \N__3726\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3726\,
            I => \N__3723\
        );

    \I__534\ : Span4Mux_v
    port map (
            O => \N__3723\,
            I => \N__3720\
        );

    \I__533\ : Odrv4
    port map (
            O => \N__3720\,
            I => \U409_ADDRESS_DECODE_AUTOCONFIG_SPACE_6\
        );

    \I__532\ : IoInMux
    port map (
            O => \N__3717\,
            I => \N__3714\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__3714\,
            I => \N__3711\
        );

    \I__530\ : Span4Mux_s3_v
    port map (
            O => \N__3711\,
            I => \N__3708\
        );

    \I__529\ : Span4Mux_h
    port map (
            O => \N__3708\,
            I => \N__3705\
        );

    \I__528\ : Sp12to4
    port map (
            O => \N__3705\,
            I => \N__3702\
        );

    \I__527\ : Span12Mux_h
    port map (
            O => \N__3702\,
            I => \N__3699\
        );

    \I__526\ : Odrv12
    port map (
            O => \N__3699\,
            I => \BUFENn_c\
        );

    \I__525\ : InMux
    port map (
            O => \N__3696\,
            I => \N__3689\
        );

    \I__524\ : InMux
    port map (
            O => \N__3695\,
            I => \N__3689\
        );

    \I__523\ : InMux
    port map (
            O => \N__3694\,
            I => \N__3686\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__3689\,
            I => \N__3681\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3686\,
            I => \N__3678\
        );

    \I__520\ : CascadeMux
    port map (
            O => \N__3685\,
            I => \N__3675\
        );

    \I__519\ : CascadeMux
    port map (
            O => \N__3684\,
            I => \N__3672\
        );

    \I__518\ : Span4Mux_v
    port map (
            O => \N__3681\,
            I => \N__3669\
        );

    \I__517\ : Span4Mux_v
    port map (
            O => \N__3678\,
            I => \N__3666\
        );

    \I__516\ : InMux
    port map (
            O => \N__3675\,
            I => \N__3663\
        );

    \I__515\ : InMux
    port map (
            O => \N__3672\,
            I => \N__3660\
        );

    \I__514\ : Sp12to4
    port map (
            O => \N__3669\,
            I => \N__3650\
        );

    \I__513\ : Sp12to4
    port map (
            O => \N__3666\,
            I => \N__3650\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__3663\,
            I => \N__3650\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3660\,
            I => \N__3650\
        );

    \I__510\ : InMux
    port map (
            O => \N__3659\,
            I => \N__3647\
        );

    \I__509\ : Span12Mux_h
    port map (
            O => \N__3650\,
            I => \N__3644\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__3647\,
            I => \N__3641\
        );

    \I__507\ : Span12Mux_v
    port map (
            O => \N__3644\,
            I => \N__3638\
        );

    \I__506\ : Span12Mux_h
    port map (
            O => \N__3641\,
            I => \N__3635\
        );

    \I__505\ : Odrv12
    port map (
            O => \N__3638\,
            I => \TM_c_0\
        );

    \I__504\ : Odrv12
    port map (
            O => \N__3635\,
            I => \TM_c_0\
        );

    \I__503\ : InMux
    port map (
            O => \N__3630\,
            I => \N__3627\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__3627\,
            I => \N__3623\
        );

    \I__501\ : InMux
    port map (
            O => \N__3626\,
            I => \N__3620\
        );

    \I__500\ : Span4Mux_v
    port map (
            O => \N__3623\,
            I => \N__3615\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__3620\,
            I => \N__3615\
        );

    \I__498\ : Span4Mux_v
    port map (
            O => \N__3615\,
            I => \N__3612\
        );

    \I__497\ : Odrv4
    port map (
            O => \N__3612\,
            I => \U409_ADDRESS_DECODE.un2_REGSPACEn_0\
        );

    \I__496\ : CascadeMux
    port map (
            O => \N__3609\,
            I => \N__3602\
        );

    \I__495\ : InMux
    port map (
            O => \N__3608\,
            I => \N__3599\
        );

    \I__494\ : InMux
    port map (
            O => \N__3607\,
            I => \N__3596\
        );

    \I__493\ : InMux
    port map (
            O => \N__3606\,
            I => \N__3588\
        );

    \I__492\ : InMux
    port map (
            O => \N__3605\,
            I => \N__3588\
        );

    \I__491\ : InMux
    port map (
            O => \N__3602\,
            I => \N__3588\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3599\,
            I => \N__3585\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__3596\,
            I => \N__3582\
        );

    \I__488\ : CascadeMux
    port map (
            O => \N__3595\,
            I => \N__3579\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__3588\,
            I => \N__3576\
        );

    \I__486\ : Span4Mux_h
    port map (
            O => \N__3585\,
            I => \N__3571\
        );

    \I__485\ : Span4Mux_v
    port map (
            O => \N__3582\,
            I => \N__3571\
        );

    \I__484\ : InMux
    port map (
            O => \N__3579\,
            I => \N__3568\
        );

    \I__483\ : Span12Mux_h
    port map (
            O => \N__3576\,
            I => \N__3565\
        );

    \I__482\ : Span4Mux_v
    port map (
            O => \N__3571\,
            I => \N__3562\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__3568\,
            I => \N__3559\
        );

    \I__480\ : Odrv12
    port map (
            O => \N__3565\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0\
        );

    \I__479\ : Odrv4
    port map (
            O => \N__3562\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0\
        );

    \I__478\ : Odrv12
    port map (
            O => \N__3559\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0\
        );

    \I__477\ : CascadeMux
    port map (
            O => \N__3552\,
            I => \N__3549\
        );

    \I__476\ : InMux
    port map (
            O => \N__3549\,
            I => \N__3540\
        );

    \I__475\ : InMux
    port map (
            O => \N__3548\,
            I => \N__3540\
        );

    \I__474\ : InMux
    port map (
            O => \N__3547\,
            I => \N__3537\
        );

    \I__473\ : InMux
    port map (
            O => \N__3546\,
            I => \N__3534\
        );

    \I__472\ : InMux
    port map (
            O => \N__3545\,
            I => \N__3530\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__3540\,
            I => \N__3525\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3537\,
            I => \N__3525\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3534\,
            I => \N__3522\
        );

    \I__468\ : InMux
    port map (
            O => \N__3533\,
            I => \N__3519\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__3530\,
            I => \N__3516\
        );

    \I__466\ : Span4Mux_v
    port map (
            O => \N__3525\,
            I => \N__3509\
        );

    \I__465\ : Span4Mux_h
    port map (
            O => \N__3522\,
            I => \N__3509\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__3519\,
            I => \N__3509\
        );

    \I__463\ : Span4Mux_v
    port map (
            O => \N__3516\,
            I => \N__3506\
        );

    \I__462\ : Span4Mux_h
    port map (
            O => \N__3509\,
            I => \N__3503\
        );

    \I__461\ : Sp12to4
    port map (
            O => \N__3506\,
            I => \N__3500\
        );

    \I__460\ : Sp12to4
    port map (
            O => \N__3503\,
            I => \N__3497\
        );

    \I__459\ : Span12Mux_h
    port map (
            O => \N__3500\,
            I => \N__3494\
        );

    \I__458\ : Odrv12
    port map (
            O => \N__3497\,
            I => \TM_c_1\
        );

    \I__457\ : Odrv12
    port map (
            O => \N__3494\,
            I => \TM_c_1\
        );

    \I__456\ : IoInMux
    port map (
            O => \N__3489\,
            I => \N__3486\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__3486\,
            I => \N__3483\
        );

    \I__454\ : Span4Mux_s1_v
    port map (
            O => \N__3483\,
            I => \N__3480\
        );

    \I__453\ : Span4Mux_h
    port map (
            O => \N__3480\,
            I => \N__3477\
        );

    \I__452\ : Sp12to4
    port map (
            O => \N__3477\,
            I => \N__3474\
        );

    \I__451\ : Span12Mux_h
    port map (
            O => \N__3474\,
            I => \N__3471\
        );

    \I__450\ : Odrv12
    port map (
            O => \N__3471\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\
        );

    \I__449\ : InMux
    port map (
            O => \N__3468\,
            I => \N__3465\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__3465\,
            I => \U409_TRANSFER_ACK.N_38\
        );

    \I__447\ : CascadeMux
    port map (
            O => \N__3462\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3Z0Z_2_cascade_\
        );

    \I__446\ : InMux
    port map (
            O => \N__3459\,
            I => \N__3456\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__3456\,
            I => \N__3451\
        );

    \I__444\ : InMux
    port map (
            O => \N__3455\,
            I => \N__3448\
        );

    \I__443\ : InMux
    port map (
            O => \N__3454\,
            I => \N__3445\
        );

    \I__442\ : Odrv4
    port map (
            O => \N__3451\,
            I => \U409_ADDRESS_DECODE.CIA_SPACE_6\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__3448\,
            I => \U409_ADDRESS_DECODE.CIA_SPACE_6\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__3445\,
            I => \U409_ADDRESS_DECODE.CIA_SPACE_6\
        );

    \I__439\ : CascadeMux
    port map (
            O => \N__3438\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENn_2_cascade_\
        );

    \I__438\ : CascadeMux
    port map (
            O => \N__3435\,
            I => \N__3431\
        );

    \I__437\ : CascadeMux
    port map (
            O => \N__3434\,
            I => \N__3428\
        );

    \I__436\ : InMux
    port map (
            O => \N__3431\,
            I => \N__3423\
        );

    \I__435\ : InMux
    port map (
            O => \N__3428\,
            I => \N__3420\
        );

    \I__434\ : InMux
    port map (
            O => \N__3427\,
            I => \N__3417\
        );

    \I__433\ : InMux
    port map (
            O => \N__3426\,
            I => \N__3414\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__3423\,
            I => \N__3407\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__3420\,
            I => \N__3407\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__3417\,
            I => \N__3402\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__3414\,
            I => \N__3402\
        );

    \I__428\ : InMux
    port map (
            O => \N__3413\,
            I => \N__3397\
        );

    \I__427\ : InMux
    port map (
            O => \N__3412\,
            I => \N__3397\
        );

    \I__426\ : Span4Mux_v
    port map (
            O => \N__3407\,
            I => \N__3393\
        );

    \I__425\ : Span4Mux_v
    port map (
            O => \N__3402\,
            I => \N__3388\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__3397\,
            I => \N__3388\
        );

    \I__423\ : InMux
    port map (
            O => \N__3396\,
            I => \N__3385\
        );

    \I__422\ : Sp12to4
    port map (
            O => \N__3393\,
            I => \N__3378\
        );

    \I__421\ : Sp12to4
    port map (
            O => \N__3388\,
            I => \N__3378\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__3385\,
            I => \N__3378\
        );

    \I__419\ : Odrv12
    port map (
            O => \N__3378\,
            I => \A_c_20\
        );

    \I__418\ : InMux
    port map (
            O => \N__3375\,
            I => \N__3372\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3372\,
            I => \U409_ADDRESS_DECODE.REGISTER_SPACEZ0\
        );

    \I__416\ : CascadeMux
    port map (
            O => \N__3369\,
            I => \U409_ADDRESS_DECODE.RANGER_SPACEZ0Z_2_cascade_\
        );

    \I__415\ : InMux
    port map (
            O => \N__3366\,
            I => \N__3362\
        );

    \I__414\ : InMux
    port map (
            O => \N__3365\,
            I => \N__3358\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__3362\,
            I => \N__3353\
        );

    \I__412\ : InMux
    port map (
            O => \N__3361\,
            I => \N__3350\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__3358\,
            I => \N__3347\
        );

    \I__410\ : InMux
    port map (
            O => \N__3357\,
            I => \N__3344\
        );

    \I__409\ : InMux
    port map (
            O => \N__3356\,
            I => \N__3341\
        );

    \I__408\ : Span4Mux_v
    port map (
            O => \N__3353\,
            I => \N__3336\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__3350\,
            I => \N__3336\
        );

    \I__406\ : Span4Mux_v
    port map (
            O => \N__3347\,
            I => \N__3329\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__3344\,
            I => \N__3329\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__3341\,
            I => \N__3329\
        );

    \I__403\ : Span4Mux_v
    port map (
            O => \N__3336\,
            I => \N__3326\
        );

    \I__402\ : Span4Mux_v
    port map (
            O => \N__3329\,
            I => \N__3323\
        );

    \I__401\ : Sp12to4
    port map (
            O => \N__3326\,
            I => \N__3318\
        );

    \I__400\ : Sp12to4
    port map (
            O => \N__3323\,
            I => \N__3318\
        );

    \I__399\ : Span12Mux_h
    port map (
            O => \N__3318\,
            I => \N__3315\
        );

    \I__398\ : Span12Mux_v
    port map (
            O => \N__3315\,
            I => \N__3312\
        );

    \I__397\ : Odrv12
    port map (
            O => \N__3312\,
            I => \A_c_19\
        );

    \I__396\ : CascadeMux
    port map (
            O => \N__3309\,
            I => \N__3306\
        );

    \I__395\ : InMux
    port map (
            O => \N__3306\,
            I => \N__3299\
        );

    \I__394\ : InMux
    port map (
            O => \N__3305\,
            I => \N__3299\
        );

    \I__393\ : InMux
    port map (
            O => \N__3304\,
            I => \N__3296\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__3299\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__3296\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4\
        );

    \I__390\ : InMux
    port map (
            O => \N__3291\,
            I => \N__3288\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__3288\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_1\
        );

    \I__388\ : CascadeMux
    port map (
            O => \N__3285\,
            I => \N__3282\
        );

    \I__387\ : InMux
    port map (
            O => \N__3282\,
            I => \N__3274\
        );

    \I__386\ : InMux
    port map (
            O => \N__3281\,
            I => \N__3274\
        );

    \I__385\ : InMux
    port map (
            O => \N__3280\,
            I => \N__3269\
        );

    \I__384\ : InMux
    port map (
            O => \N__3279\,
            I => \N__3269\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__3274\,
            I => \N__3264\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__3269\,
            I => \N__3264\
        );

    \I__381\ : Span4Mux_v
    port map (
            O => \N__3264\,
            I => \N__3261\
        );

    \I__380\ : Span4Mux_v
    port map (
            O => \N__3261\,
            I => \N__3258\
        );

    \I__379\ : Span4Mux_v
    port map (
            O => \N__3258\,
            I => \N__3255\
        );

    \I__378\ : Sp12to4
    port map (
            O => \N__3255\,
            I => \N__3252\
        );

    \I__377\ : Odrv12
    port map (
            O => \N__3252\,
            I => \A_c_16\
        );

    \I__376\ : InMux
    port map (
            O => \N__3249\,
            I => \N__3240\
        );

    \I__375\ : InMux
    port map (
            O => \N__3248\,
            I => \N__3240\
        );

    \I__374\ : InMux
    port map (
            O => \N__3247\,
            I => \N__3240\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__3240\,
            I => \N__3237\
        );

    \I__372\ : Span4Mux_v
    port map (
            O => \N__3237\,
            I => \N__3234\
        );

    \I__371\ : Sp12to4
    port map (
            O => \N__3234\,
            I => \N__3231\
        );

    \I__370\ : Span12Mux_v
    port map (
            O => \N__3231\,
            I => \N__3228\
        );

    \I__369\ : Odrv12
    port map (
            O => \N__3228\,
            I => \A_c_17\
        );

    \I__368\ : CascadeMux
    port map (
            O => \N__3225\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3_cascade_\
        );

    \I__367\ : CascadeMux
    port map (
            O => \N__3222\,
            I => \U409_ADDRESS_DECODE_AUTOVECTOR_5_cascade_\
        );

    \I__366\ : CascadeMux
    port map (
            O => \N__3219\,
            I => \N__3216\
        );

    \I__365\ : InMux
    port map (
            O => \N__3216\,
            I => \N__3212\
        );

    \I__364\ : InMux
    port map (
            O => \N__3215\,
            I => \N__3209\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__3212\,
            I => \N__3204\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__3209\,
            I => \N__3204\
        );

    \I__361\ : Span4Mux_v
    port map (
            O => \N__3204\,
            I => \N__3200\
        );

    \I__360\ : InMux
    port map (
            O => \N__3203\,
            I => \N__3197\
        );

    \I__359\ : Sp12to4
    port map (
            O => \N__3200\,
            I => \N__3192\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__3197\,
            I => \N__3192\
        );

    \I__357\ : Span12Mux_h
    port map (
            O => \N__3192\,
            I => \N__3189\
        );

    \I__356\ : Span12Mux_v
    port map (
            O => \N__3189\,
            I => \N__3186\
        );

    \I__355\ : Odrv12
    port map (
            O => \N__3186\,
            I => \A_c_18\
        );

    \I__354\ : InMux
    port map (
            O => \N__3183\,
            I => \N__3179\
        );

    \I__353\ : InMux
    port map (
            O => \N__3182\,
            I => \N__3176\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__3179\,
            I => \N__3173\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__3176\,
            I => \N__3170\
        );

    \I__350\ : Span4Mux_h
    port map (
            O => \N__3173\,
            I => \N__3167\
        );

    \I__349\ : Span12Mux_h
    port map (
            O => \N__3170\,
            I => \N__3164\
        );

    \I__348\ : Span4Mux_v
    port map (
            O => \N__3167\,
            I => \N__3161\
        );

    \I__347\ : Odrv12
    port map (
            O => \N__3164\,
            I => \U409_ADDRESS_DECODE.AUTOVECTOR_16\
        );

    \I__346\ : Odrv4
    port map (
            O => \N__3161\,
            I => \U409_ADDRESS_DECODE.AUTOVECTOR_16\
        );

    \I__345\ : InMux
    port map (
            O => \N__3156\,
            I => \N__3153\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__3153\,
            I => \N__3150\
        );

    \I__343\ : Span4Mux_v
    port map (
            O => \N__3150\,
            I => \N__3147\
        );

    \I__342\ : Span4Mux_v
    port map (
            O => \N__3147\,
            I => \N__3144\
        );

    \I__341\ : IoSpan4Mux
    port map (
            O => \N__3144\,
            I => \N__3141\
        );

    \I__340\ : Odrv4
    port map (
            O => \N__3141\,
            I => \TT_c_1\
        );

    \I__339\ : InMux
    port map (
            O => \N__3138\,
            I => \N__3135\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__3135\,
            I => \N__3132\
        );

    \I__337\ : Span4Mux_v
    port map (
            O => \N__3132\,
            I => \N__3129\
        );

    \I__336\ : Span4Mux_v
    port map (
            O => \N__3129\,
            I => \N__3126\
        );

    \I__335\ : IoSpan4Mux
    port map (
            O => \N__3126\,
            I => \N__3123\
        );

    \I__334\ : Odrv4
    port map (
            O => \N__3123\,
            I => \TT_c_0\
        );

    \I__333\ : InMux
    port map (
            O => \N__3120\,
            I => \N__3117\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__3117\,
            I => \N__3114\
        );

    \I__331\ : Odrv12
    port map (
            O => \N__3114\,
            I => \U409_ADDRESS_DECODE_AUTOVECTOR_4\
        );

    \I__330\ : InMux
    port map (
            O => \N__3111\,
            I => \N__3105\
        );

    \I__329\ : InMux
    port map (
            O => \N__3110\,
            I => \N__3105\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__3105\,
            I => \N__3102\
        );

    \I__327\ : Span4Mux_v
    port map (
            O => \N__3102\,
            I => \N__3099\
        );

    \I__326\ : Span4Mux_h
    port map (
            O => \N__3099\,
            I => \N__3096\
        );

    \I__325\ : Odrv4
    port map (
            O => \N__3096\,
            I => \A_c_31\
        );

    \I__324\ : InMux
    port map (
            O => \N__3093\,
            I => \N__3087\
        );

    \I__323\ : InMux
    port map (
            O => \N__3092\,
            I => \N__3087\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__3087\,
            I => \N__3084\
        );

    \I__321\ : Span4Mux_v
    port map (
            O => \N__3084\,
            I => \N__3081\
        );

    \I__320\ : Sp12to4
    port map (
            O => \N__3081\,
            I => \N__3078\
        );

    \I__319\ : Odrv12
    port map (
            O => \N__3078\,
            I => \A_c_30\
        );

    \I__318\ : InMux
    port map (
            O => \N__3075\,
            I => \N__3072\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__3072\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5\
        );

    \I__316\ : CascadeMux
    port map (
            O => \N__3069\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_\
        );

    \I__315\ : CascadeMux
    port map (
            O => \N__3066\,
            I => \N__3063\
        );

    \I__314\ : InMux
    port map (
            O => \N__3063\,
            I => \N__3057\
        );

    \I__313\ : InMux
    port map (
            O => \N__3062\,
            I => \N__3057\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__3057\,
            I => \N__3054\
        );

    \I__311\ : Span4Mux_v
    port map (
            O => \N__3054\,
            I => \N__3051\
        );

    \I__310\ : Span4Mux_v
    port map (
            O => \N__3051\,
            I => \N__3048\
        );

    \I__309\ : Sp12to4
    port map (
            O => \N__3048\,
            I => \N__3045\
        );

    \I__308\ : Odrv12
    port map (
            O => \N__3045\,
            I => \A_c_26\
        );

    \I__307\ : InMux
    port map (
            O => \N__3042\,
            I => \N__3036\
        );

    \I__306\ : InMux
    port map (
            O => \N__3041\,
            I => \N__3036\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__3036\,
            I => \N__3033\
        );

    \I__304\ : Span4Mux_h
    port map (
            O => \N__3033\,
            I => \N__3030\
        );

    \I__303\ : Span4Mux_v
    port map (
            O => \N__3030\,
            I => \N__3027\
        );

    \I__302\ : Odrv4
    port map (
            O => \N__3027\,
            I => \A_c_24\
        );

    \I__301\ : CascadeMux
    port map (
            O => \N__3024\,
            I => \N__3020\
        );

    \I__300\ : InMux
    port map (
            O => \N__3023\,
            I => \N__3017\
        );

    \I__299\ : InMux
    port map (
            O => \N__3020\,
            I => \N__3014\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__3017\,
            I => \N__3009\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__3014\,
            I => \N__3009\
        );

    \I__296\ : Span4Mux_v
    port map (
            O => \N__3009\,
            I => \N__3006\
        );

    \I__295\ : Sp12to4
    port map (
            O => \N__3006\,
            I => \N__3003\
        );

    \I__294\ : Odrv12
    port map (
            O => \N__3003\,
            I => \A_c_27\
        );

    \I__293\ : InMux
    port map (
            O => \N__3000\,
            I => \N__2994\
        );

    \I__292\ : InMux
    port map (
            O => \N__2999\,
            I => \N__2994\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__2994\,
            I => \N__2991\
        );

    \I__290\ : Span4Mux_v
    port map (
            O => \N__2991\,
            I => \N__2988\
        );

    \I__289\ : Span4Mux_h
    port map (
            O => \N__2988\,
            I => \N__2985\
        );

    \I__288\ : Odrv4
    port map (
            O => \N__2985\,
            I => \A_c_25\
        );

    \I__287\ : InMux
    port map (
            O => \N__2982\,
            I => \N__2979\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__2979\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_3\
        );

    \I__285\ : InMux
    port map (
            O => \N__2976\,
            I => \N__2970\
        );

    \I__284\ : InMux
    port map (
            O => \N__2975\,
            I => \N__2970\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__2970\,
            I => \N__2967\
        );

    \I__282\ : Span4Mux_h
    port map (
            O => \N__2967\,
            I => \N__2964\
        );

    \I__281\ : Span4Mux_v
    port map (
            O => \N__2964\,
            I => \N__2961\
        );

    \I__280\ : Odrv4
    port map (
            O => \N__2961\,
            I => \A_c_29\
        );

    \I__279\ : CascadeMux
    port map (
            O => \N__2958\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_4_cascade_\
        );

    \I__278\ : InMux
    port map (
            O => \N__2955\,
            I => \N__2949\
        );

    \I__277\ : InMux
    port map (
            O => \N__2954\,
            I => \N__2949\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__2949\,
            I => \N__2946\
        );

    \I__275\ : Span4Mux_v
    port map (
            O => \N__2946\,
            I => \N__2943\
        );

    \I__274\ : Span4Mux_v
    port map (
            O => \N__2943\,
            I => \N__2940\
        );

    \I__273\ : Sp12to4
    port map (
            O => \N__2940\,
            I => \N__2937\
        );

    \I__272\ : Odrv12
    port map (
            O => \N__2937\,
            I => \A_c_28\
        );

    \I__271\ : IoInMux
    port map (
            O => \N__2934\,
            I => \N__2931\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2931\,
            I => \N__2928\
        );

    \I__269\ : Span12Mux_s11_h
    port map (
            O => \N__2928\,
            I => \N__2925\
        );

    \I__268\ : Span12Mux_h
    port map (
            O => \N__2925\,
            I => \N__2922\
        );

    \I__267\ : Odrv12
    port map (
            O => \N__2922\,
            I => \U409_ADDRESS_DECODE_un1_RTC_ENn_i\
        );

    \I__266\ : InMux
    port map (
            O => \N__2919\,
            I => \N__2916\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__2916\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_1\
        );

    \I__264\ : CascadeMux
    port map (
            O => \N__2913\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_1_cascade_\
        );

    \I__263\ : InMux
    port map (
            O => \N__2910\,
            I => \N__2904\
        );

    \I__262\ : InMux
    port map (
            O => \N__2909\,
            I => \N__2904\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__2904\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3\
        );

    \I__260\ : ClkMux
    port map (
            O => \N__2901\,
            I => \N__2868\
        );

    \I__259\ : ClkMux
    port map (
            O => \N__2900\,
            I => \N__2868\
        );

    \I__258\ : ClkMux
    port map (
            O => \N__2899\,
            I => \N__2868\
        );

    \I__257\ : ClkMux
    port map (
            O => \N__2898\,
            I => \N__2868\
        );

    \I__256\ : ClkMux
    port map (
            O => \N__2897\,
            I => \N__2868\
        );

    \I__255\ : ClkMux
    port map (
            O => \N__2896\,
            I => \N__2868\
        );

    \I__254\ : ClkMux
    port map (
            O => \N__2895\,
            I => \N__2868\
        );

    \I__253\ : ClkMux
    port map (
            O => \N__2894\,
            I => \N__2868\
        );

    \I__252\ : ClkMux
    port map (
            O => \N__2893\,
            I => \N__2868\
        );

    \I__251\ : ClkMux
    port map (
            O => \N__2892\,
            I => \N__2868\
        );

    \I__250\ : ClkMux
    port map (
            O => \N__2891\,
            I => \N__2868\
        );

    \I__249\ : GlobalMux
    port map (
            O => \N__2868\,
            I => \CLK80_OUT\
        );

    \INVU409_TRANSFER_ACK.TACK_EN_iC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            I => \N__2898\
        );

    \INVU409_TRANSFER_ACK.TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            I => \N__2896\
        );

    \INVU409_TRANSFER_ACK.IRQ_TACK_EN_nesrC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.IRQ_TACK_EN_nesrC_net\,
            I => \N__2894\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            I => \N__2892\
        );

    \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            I => \N__2897\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            I => \N__2895\
        );

    \INVU409_TRANSFER_ACK.CIA_ENABLED_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\,
            I => \N__2893\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            I => \N__2891\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net\,
            I => \N__2901\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            I => \N__2899\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            I => \N__2900\
        );

    \IN_MUX_bfv_14_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_4_0_\
        );

    \IN_MUX_bfv_14_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un3_COUNTER60_1_cry_8\,
            carryinitout => \bfn_14_5_0_\
        );

    \IN_MUX_bfv_14_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_1_0_\
        );

    \IN_MUX_bfv_14_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un2_COUNTER50_1_cry_8\,
            carryinitout => \bfn_14_2_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_8_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__5886\,
            in1 => \N__3023\,
            in2 => \N__3066\,
            in3 => \N__3000\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_3_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3092\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3110\,
            lcout => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__3111\,
            in1 => \N__3042\,
            in2 => \_gnd_net_\,
            in3 => \N__3093\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__3075\,
            in1 => \N__2976\,
            in2 => \N__3069\,
            in3 => \N__2955\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_4_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3062\,
            in1 => \N__3041\,
            in2 => \N__3024\,
            in3 => \N__2999\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2982\,
            in1 => \N__2975\,
            in2 => \N__2958\,
            in3 => \N__2954\,
            lcout => \U409_ADDRESS_DECODE.AUTOVECTOR_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__3280\,
            in1 => \N__2910\,
            in2 => \N__3309\,
            in3 => \N__2919\,
            lcout => \U409_ADDRESS_DECODE_un1_RTC_ENn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_1_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3203\,
            in1 => \N__3898\,
            in2 => \N__3435\,
            in3 => \N__3356\,
            lcout => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_1\,
            ltout => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__2909\,
            in1 => \N__3279\,
            in2 => \N__2913\,
            in3 => \N__3305\,
            lcout => \U409_ADDRESS_DECODE_un1_RTC_ENn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_3_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__3607\,
            in1 => \N__3249\,
            in2 => \_gnd_net_\,
            in3 => \N__3807\,
            lcout => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_6_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3281\,
            in1 => \N__3806\,
            in2 => \N__3434\,
            in3 => \N__3247\,
            lcout => \U409_ADDRESS_DECODE_AUTOCONFIG_SPACE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3357\,
            in1 => \N__3215\,
            in2 => \N__3285\,
            in3 => \N__3248\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3805\,
            in2 => \_gnd_net_\,
            in3 => \N__3396\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_5_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3454\,
            in1 => \N__3182\,
            in2 => \N__3225\,
            in3 => \N__3964\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE_AUTOVECTOR_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__3120\,
            in1 => \N__4019\,
            in2 => \N__3222\,
            in3 => \N__5870\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_7_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__3365\,
            in1 => \N__3963\,
            in2 => \N__3219\,
            in3 => \N__3183\,
            lcout => \U409_ADDRESS_DECODE_AUTOCONFIG_SPACE_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_4_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3894\,
            in1 => \N__3156\,
            in2 => \N__5885\,
            in3 => \N__3138\,
            lcout => \U409_ADDRESS_DECODE_AUTOVECTOR_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_0_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__4083\,
            in1 => \N__3979\,
            in2 => \N__3825\,
            in3 => \N__3899\,
            lcout => \U409_TRANSFER_ACK.N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__3547\,
            in1 => \N__3978\,
            in2 => \_gnd_net_\,
            in3 => \N__3694\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_2_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3980\,
            in1 => \N__3427\,
            in2 => \_gnd_net_\,
            in3 => \N__3823\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__3468\,
            in1 => \N__3361\,
            in2 => \N__3462\,
            in3 => \N__3900\,
            lcout => \U409_TRANSFER_ACK.N_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_1_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3455\,
            in1 => \N__3819\,
            in2 => \_gnd_net_\,
            in3 => \N__3426\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.REGISTER_SPACE_3_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3876\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3413\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.un1_RTC_ENn_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.REGISTER_SPACE_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__3459\,
            in1 => \N__3817\,
            in2 => \N__3438\,
            in3 => \N__3976\,
            lcout => \U409_ADDRESS_DECODE.REGISTER_SPACEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.RANGER_SPACE_2_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__3412\,
            in1 => \N__3975\,
            in2 => \_gnd_net_\,
            in3 => \N__3816\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.RANGER_SPACEZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un2_REGSPACEn_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__3877\,
            in1 => \N__3375\,
            in2 => \N__3369\,
            in3 => \N__3366\,
            lcout => \U409_ADDRESS_DECODE.un2_REGSPACEn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_5_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000000000"
        )
    port map (
            in0 => \N__3533\,
            in1 => \N__3875\,
            in2 => \N__3684\,
            in3 => \N__5878\,
            lcout => \U409_ADDRESS_DECODE_AUTOCONFIG_SPACE_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__3304\,
            in1 => \N__3901\,
            in2 => \N__3609\,
            in3 => \N__3291\,
            lcout => \CIA_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_1_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__3695\,
            in1 => \N__3605\,
            in2 => \_gnd_net_\,
            in3 => \N__3548\,
            lcout => \U409_ADDRESS_DECODE_ROMEN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_0_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__3606\,
            in1 => \N__3696\,
            in2 => \N__3552\,
            in3 => \N__4079\,
            lcout => \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0\,
            ltout => \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__3902\,
            in1 => \N__3981\,
            in2 => \N__4047\,
            in3 => \N__3824\,
            lcout => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4124\,
            in1 => \N__4023\,
            in2 => \_gnd_net_\,
            in3 => \N__4209\,
            lcout => \PORTSIZE_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__3977\,
            in1 => \N__3918\,
            in2 => \N__3909\,
            in3 => \N__3818\,
            lcout => \U409_ADDRESS_DECODE_un1_RAMSPACEn\,
            ltout => \U409_ADDRESS_DECODE_un1_RAMSPACEn_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__4207\,
            in1 => \_gnd_net_\,
            in2 => \N__3750\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \AGNUS_SPACE_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_DATA_BUFFERS.un1_BUFENn_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__3747\,
            in1 => \N__3741\,
            in2 => \N__3732\,
            in3 => \N__3729\,
            lcout => \BUFENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__3626\,
            in1 => \N__3608\,
            in2 => \N__3685\,
            in3 => \N__3546\,
            lcout => \U409_ADDRESS_DECODE_un1_REGSPACEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__3659\,
            in1 => \N__3630\,
            in2 => \N__3595\,
            in3 => \N__3545\,
            lcout => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_0_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__4104\,
            in1 => \N__4275\,
            in2 => \N__4428\,
            in3 => \N__4475\,
            lcout => OPEN,
            ltout => \U409_CIA.VMA_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__4476\,
            in1 => \N__4128\,
            in2 => \N__4107\,
            in3 => \N__5155\,
            lcout => \U409_CIA.VMAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_1_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__4564\,
            in1 => \N__4635\,
            in2 => \N__4506\,
            in3 => \N__4538\,
            lcout => \U409_CIA.un1_CIA_CLK_COUNT_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4463\,
            in2 => \N__4542\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_2_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4631\,
            in2 => \_gnd_net_\,
            in3 => \N__4098\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            clk => \N__4583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4380\,
            in2 => \_gnd_net_\,
            in3 => \N__4095\,
            lcout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_4_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4415\,
            in2 => \_gnd_net_\,
            in3 => \N__4092\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            clk => \N__4583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4610\,
            in2 => \_gnd_net_\,
            in3 => \N__4089\,
            lcout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_6_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4566\,
            in2 => \_gnd_net_\,
            in3 => \N__4086\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\,
            clk => \N__4583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_7_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4504\,
            in2 => \_gnd_net_\,
            in3 => \N__4227\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_1_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4541\,
            in2 => \_gnd_net_\,
            in3 => \N__4473\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__4884\,
            in1 => \N__4350\,
            in2 => \_gnd_net_\,
            in3 => \N__4682\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__4987\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4217\,
            in2 => \N__4689\,
            in3 => \N__4861\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__4987\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__4862\,
            in1 => \N__4878\,
            in2 => \N__4221\,
            in3 => \N__4686\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__4987\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIF4AR_5_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4816\,
            in2 => \_gnd_net_\,
            in3 => \N__4348\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1\,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_3_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4783\,
            in2 => \N__4224\,
            in3 => \N__4798\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__4208\,
            in1 => \N__4191\,
            in2 => \N__5877\,
            in3 => \N__4182\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_10_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4164\,
            in2 => \_gnd_net_\,
            in3 => \N__4290\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS1n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4286\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4323\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS0n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNI692L_0_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5837\,
            in1 => \N__5156\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CIA_ENABLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNICGRM_3_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4604\,
            in2 => \_gnd_net_\,
            in3 => \N__4379\,
            lcout => \U409_CIA.CLK_CIA6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_0_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__4274\,
            in1 => \N__4634\,
            in2 => \N__4424\,
            in3 => \N__4437\,
            lcout => OPEN,
            ltout => \U409_CIA.CLK_CIA6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4903\,
            in2 => \N__4263\,
            in3 => \N__4356\,
            lcout => \CLK_CIA_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_3_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100101010"
        )
    port map (
            in0 => \N__4383\,
            in1 => \N__4254\,
            in2 => \N__4239\,
            in3 => \N__4260\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_3_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__4633\,
            in1 => \N__4382\,
            in2 => \N__4611\,
            in3 => \N__4539\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_2_0\,
            ltout => \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_5_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001101001100"
        )
    port map (
            in0 => \N__4238\,
            in1 => \N__4609\,
            in2 => \N__4248\,
            in3 => \N__4245\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__4565\,
            in1 => \N__4503\,
            in2 => \N__4474\,
            in3 => \N__4420\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_2_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4632\,
            in2 => \_gnd_net_\,
            in3 => \N__4605\,
            lcout => \U409_CIA.un1_CIA_CLK_COUNT_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_0_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4540\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIMUMD1_7_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4563\,
            in1 => \N__4537\,
            in2 => \N__4505\,
            in3 => \N__4464\,
            lcout => \U409_CIA.CLK_CIA6_3\,
            ltout => \U409_CIA.CLK_CIA6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_1_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4416\,
            in1 => \N__4392\,
            in2 => \N__4386\,
            in3 => \N__4381\,
            lcout => \U409_CIA.CLK_CIA_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__5292\,
            in1 => \N__4733\,
            in2 => \_gnd_net_\,
            in3 => \N__4833\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            ce => 'H',
            sr => \N__4995\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_5_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4876\,
            in1 => \N__4823\,
            in2 => \N__4863\,
            in3 => \N__4349\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_0_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4781\,
            in1 => \N__4716\,
            in2 => \N__4332\,
            in3 => \N__4329\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4652\,
            in2 => \_gnd_net_\,
            in3 => \N__4749\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010000000"
        )
    port map (
            in0 => \N__4653\,
            in1 => \N__4714\,
            in2 => \N__4758\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4824\,
            in2 => \N__4887\,
            in3 => \N__4782\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__4654\,
            in1 => \N__4877\,
            in2 => \N__4757\,
            in3 => \N__4857\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4715\,
            in1 => \N__4780\,
            in2 => \N__4842\,
            in3 => \N__4839\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_0_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__5523\,
            in1 => \N__5590\,
            in2 => \N__4827\,
            in3 => \N__4732\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__4800\,
            in1 => \N__4785\,
            in2 => \N__4688\,
            in3 => \N__4822\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net\,
            ce => 'H',
            sr => \N__4994\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__4784\,
            in1 => \N__4799\,
            in2 => \_gnd_net_\,
            in3 => \N__4675\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net\,
            ce => 'H',
            sr => \N__4994\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__4655\,
            in1 => \N__4713\,
            in2 => \_gnd_net_\,
            in3 => \N__4756\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net\,
            ce => 'H',
            sr => \N__4994\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001110011"
        )
    port map (
            in0 => \N__5583\,
            in1 => \N__4734\,
            in2 => \N__5528\,
            in3 => \N__4711\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net\,
            ce => 'H',
            sr => \N__4994\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__4712\,
            in1 => \_gnd_net_\,
            in2 => \N__4687\,
            in3 => \N__4656\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net\,
            ce => 'H',
            sr => \N__4994\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_1_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5490\,
            in1 => \N__5119\,
            in2 => \_gnd_net_\,
            in3 => \N__5099\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.m8_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100100111"
        )
    port map (
            in0 => \N__5067\,
            in1 => \N__4931\,
            in2 => \N__4962\,
            in3 => \N__5137\,
            lcout => \U409_TRANSFER_ACK.N_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000110111"
        )
    port map (
            in0 => \N__5138\,
            in1 => \N__5048\,
            in2 => \N__4935\,
            in3 => \N__4950\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.i6_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101000001000"
        )
    port map (
            in0 => \N__5822\,
            in1 => \N__5076\,
            in2 => \N__4959\,
            in3 => \N__5050\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000000100000"
        )
    port map (
            in0 => \N__5049\,
            in1 => \N__4956\,
            in2 => \N__5846\,
            in3 => \N__4941\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5118\,
            in2 => \_gnd_net_\,
            in3 => \N__5098\,
            lcout => \U409_TRANSFER_ACK.N_4\,
            ltout => \U409_TRANSFER_ACK.N_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m4_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111000001010"
        )
    port map (
            in0 => \N__5068\,
            in1 => \N__4930\,
            in2 => \N__4944\,
            in3 => \N__5136\,
            lcout => \U409_TRANSFER_ACK.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5139\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\,
            ce => 'H',
            sr => \N__5351\
        );

    \U409_TRANSFER_ACK.LASTCLK_0_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4904\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\,
            ce => 'H',
            sr => \N__5351\
        );

    \U409_TRANSFER_ACK.LASTCLK_1_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5121\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\,
            ce => 'H',
            sr => \N__5351\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5163\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5838\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\,
            ce => 'H',
            sr => \N__5351\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5682\,
            in2 => \_gnd_net_\,
            in3 => \N__5622\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_EN_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__5051\,
            in1 => \N__5120\,
            in2 => \N__5507\,
            in3 => \N__5100\,
            lcout => \U409_TRANSFER_ACK.N_138\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111100100000"
        )
    port map (
            in0 => \N__5436\,
            in1 => \N__5655\,
            in2 => \N__5085\,
            in3 => \N__5279\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            ce => 'H',
            sr => \N__5362\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100011101000000"
        )
    port map (
            in0 => \N__5075\,
            in1 => \N__5052\,
            in2 => \N__5022\,
            in3 => \N__5265\,
            lcout => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            ce => 'H',
            sr => \N__5362\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__5012\,
            in1 => \N__5495\,
            in2 => \N__5591\,
            in3 => \N__5393\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNIG3KDC_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__5013\,
            in1 => \N__5494\,
            in2 => \N__5592\,
            in3 => \N__5392\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_RNO_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5295\,
            in3 => \N__5363\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_RNIECRR_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5379\,
            in1 => \N__5291\,
            in2 => \N__5280\,
            in3 => \N__5264\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5788\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__5677\,
            in1 => \N__5619\,
            in2 => \_gnd_net_\,
            in3 => \N__5649\,
            lcout => \U409_TRANSFER_ACK.N_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5621\,
            in1 => \N__5430\,
            in2 => \N__5689\,
            in3 => \N__5650\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5681\,
            in1 => \N__5620\,
            in2 => \N__5238\,
            in3 => \N__5651\,
            lcout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__5403\,
            in1 => \N__5435\,
            in2 => \N__5237\,
            in3 => \N__5211\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5358\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100010110000"
        )
    port map (
            in0 => \N__5625\,
            in1 => \N__5434\,
            in2 => \N__5691\,
            in3 => \N__5654\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5358\
        );

    \U409_TRANSFER_ACK.ROMENn_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101110000"
        )
    port map (
            in0 => \N__5205\,
            in1 => \N__5402\,
            in2 => \N__5180\,
            in3 => \N__5199\,
            lcout => \ROMENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5358\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110001100"
        )
    port map (
            in0 => \N__5623\,
            in1 => \N__5432\,
            in2 => \N__5690\,
            in3 => \N__5652\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5358\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__5624\,
            in1 => \N__5433\,
            in2 => \_gnd_net_\,
            in3 => \N__5653\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5358\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIPTM34_0_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5571\,
            in1 => \N__5541\,
            in2 => \N__5524\,
            in3 => \N__5431\,
            lcout => \U409_TRANSFER_ACK.N_28_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5394\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_EN_nesrC_net\,
            ce => \N__5373\,
            sr => \N__5364\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011010000"
        )
    port map (
            in0 => \N__5723\,
            in1 => \N__5931\,
            in2 => \N__5847\,
            in3 => \N__5906\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100100111"
        )
    port map (
            in0 => \N__5903\,
            in1 => \N__5308\,
            in2 => \N__5933\,
            in3 => \N__5721\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111110101010"
        )
    port map (
            in0 => \N__5309\,
            in1 => \_gnd_net_\,
            in2 => \N__5322\,
            in3 => \N__5828\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__5826\,
            in1 => \N__5930\,
            in2 => \_gnd_net_\,
            in3 => \N__5905\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110110111"
        )
    port map (
            in0 => \N__5904\,
            in1 => \N__5827\,
            in2 => \N__5934\,
            in3 => \N__5722\,
            lcout => \U409_TRANSFER_ACK.TACK_OUTn_0_sqmuxa_0_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__5932\,
            in1 => \N__5907\,
            in2 => \N__5848\,
            in3 => \N__5727\,
            lcout => \TACK_EN_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            ce => \N__5706\,
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_8_LC_13_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6008\,
            in1 => \N__6039\,
            in2 => \N__5976\,
            in3 => \N__6294\,
            lcout => \U409_TICK.COUNTER60Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6770\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_4_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__5965\,
            in1 => \N__6035\,
            in2 => \N__6114\,
            in3 => \N__6001\,
            lcout => \U409_TICK.COUNTER60Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6773\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_6_LC_13_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6033\,
            in1 => \N__5966\,
            in2 => \N__6009\,
            in3 => \N__6336\,
            lcout => \U409_TICK.COUNTER60Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6773\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIHJU51_4_LC_13_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6363\,
            in1 => \N__6126\,
            in2 => \_gnd_net_\,
            in3 => \N__6174\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK603_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI335G2_11_LC_13_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6246\,
            in1 => \N__6045\,
            in2 => \N__5697\,
            in3 => \N__6141\,
            lcout => \U409_TICK.TICK603_14\,
            ltout => \U409_TICK.TICK603_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_0_LC_13_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__5964\,
            in1 => \N__6000\,
            in2 => \N__5694\,
            in3 => \N__6175\,
            lcout => \U409_TICK.COUNTER60Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6773\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_1_LC_13_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__6176\,
            in1 => \_gnd_net_\,
            in2 => \N__6201\,
            in3 => \_gnd_net_\,
            lcout => \U409_TICK.COUNTER60Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6773\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNICDC71_14_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6285\,
            in1 => \N__6486\,
            in2 => \N__6309\,
            in3 => \N__6348\,
            lcout => \U409_TICK.TICK603_9\,
            ltout => \U409_TICK.TICK603_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK60_LC_13_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__6034\,
            in1 => \N__6059\,
            in2 => \N__6075\,
            in3 => \N__5967\,
            lcout => \TICK60_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6773\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_9_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__6007\,
            in1 => \N__5968\,
            in2 => \N__6273\,
            in3 => \N__6038\,
            lcout => \U409_TICK.COUNTER60Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6775\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI2USG_10_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__6501\,
            in1 => \N__6261\,
            in2 => \N__6327\,
            in3 => \N__6465\,
            lcout => \U409_TICK.TICK603_10\,
            ltout => \U409_TICK.TICK603_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_14_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6005\,
            in1 => \N__6037\,
            in2 => \N__6048\,
            in3 => \N__6474\,
            lcout => \U409_TICK.COUNTER60Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6775\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6231\,
            in1 => \N__6156\,
            in2 => \N__6200\,
            in3 => \N__6440\,
            lcout => \U409_TICK.TICK603_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_15_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6036\,
            in1 => \N__6006\,
            in2 => \N__5975\,
            in3 => \N__6453\,
            lcout => \U409_TICK.COUNTER60Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6775\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6655\,
            in2 => \N__6411\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_1_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_2_LC_14_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6674\,
            in2 => \_gnd_net_\,
            in3 => \N__5937\,
            lcout => \U409_TICK.COUNTER50Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_1\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_2\,
            clk => \N__6769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_3_LC_14_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6422\,
            in2 => \_gnd_net_\,
            in3 => \N__6102\,
            lcout => \U409_TICK.COUNTER50Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_2\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_3\,
            clk => \N__6769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_4_LC_14_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6533\,
            in2 => \_gnd_net_\,
            in3 => \N__6099\,
            lcout => \U409_TICK.COUNTER50Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_3\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_4\,
            clk => \N__6769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_5_LC_14_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6698\,
            in2 => \_gnd_net_\,
            in3 => \N__6096\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_4\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_6_LC_14_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6578\,
            in2 => \_gnd_net_\,
            in3 => \N__6093\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_5\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_7_LC_14_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6545\,
            in2 => \_gnd_net_\,
            in3 => \N__6090\,
            lcout => \U409_TICK.COUNTER50Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_6\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_7\,
            clk => \N__6769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_8_LC_14_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6686\,
            in2 => \_gnd_net_\,
            in3 => \N__6087\,
            lcout => \U409_TICK.COUNTER50Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_7\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_8\,
            clk => \N__6769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_9_LC_14_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6593\,
            in2 => \_gnd_net_\,
            in3 => \N__6084\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_2_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_10_LC_14_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6374\,
            in2 => \_gnd_net_\,
            in3 => \N__6081\,
            lcout => \U409_TICK.COUNTER50Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_9\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_10\,
            clk => \N__6771\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_11_LC_14_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6512\,
            in2 => \_gnd_net_\,
            in3 => \N__6078\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_10\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_12_LC_14_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6389\,
            in2 => \_gnd_net_\,
            in3 => \N__6216\,
            lcout => \U409_TICK.COUNTER50Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_11\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_12\,
            clk => \N__6771\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_13_LC_14_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6557\,
            in2 => \_gnd_net_\,
            in3 => \N__6213\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_12\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_14_LC_14_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6788\,
            in2 => \_gnd_net_\,
            in3 => \N__6210\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_13\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_15_LC_14_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6923\,
            in2 => \_gnd_net_\,
            in3 => \N__6207\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_14\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_16_LC_14_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6642\,
            in2 => \_gnd_net_\,
            in3 => \N__6204\,
            lcout => \U409_TICK.COUNTER50Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6771\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6193\,
            in2 => \N__6177\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_4_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_2_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6155\,
            in2 => \_gnd_net_\,
            in3 => \N__6144\,
            lcout => \U409_TICK.COUNTER60Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_1\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_2\,
            clk => \N__6776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_3_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6140\,
            in2 => \_gnd_net_\,
            in3 => \N__6129\,
            lcout => \U409_TICK.COUNTER60Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_2\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_3\,
            clk => \N__6776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_4_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6125\,
            in2 => \_gnd_net_\,
            in3 => \N__6105\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_3\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_5_LC_14_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6362\,
            in2 => \_gnd_net_\,
            in3 => \N__6351\,
            lcout => \U409_TICK.COUNTER60Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_4\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_5\,
            clk => \N__6776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_6_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6347\,
            in2 => \_gnd_net_\,
            in3 => \N__6330\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_5\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_7_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6323\,
            in2 => \_gnd_net_\,
            in3 => \N__6312\,
            lcout => \U409_TICK.COUNTER60Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_6\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_7\,
            clk => \N__6776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_8_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6305\,
            in2 => \_gnd_net_\,
            in3 => \N__6288\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_7\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_9_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6284\,
            in2 => \_gnd_net_\,
            in3 => \N__6264\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_5_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_10_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6260\,
            in2 => \_gnd_net_\,
            in3 => \N__6249\,
            lcout => \U409_TICK.COUNTER60Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_9\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_10\,
            clk => \N__6777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_11_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6245\,
            in2 => \_gnd_net_\,
            in3 => \N__6234\,
            lcout => \U409_TICK.COUNTER60Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_10\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_11\,
            clk => \N__6777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_12_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6230\,
            in2 => \_gnd_net_\,
            in3 => \N__6219\,
            lcout => \U409_TICK.COUNTER60Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_11\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_12\,
            clk => \N__6777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_13_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6500\,
            in2 => \_gnd_net_\,
            in3 => \N__6489\,
            lcout => \U409_TICK.COUNTER60Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_12\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_13\,
            clk => \N__6777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_14_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6485\,
            in2 => \_gnd_net_\,
            in3 => \N__6468\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_13\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_15_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6464\,
            in2 => \_gnd_net_\,
            in3 => \N__6447\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_14\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_16_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6441\,
            in2 => \_gnd_net_\,
            in3 => \N__6444\,
            lcout => \U409_TICK.COUNTER60Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_6_LC_15_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6906\,
            in1 => \N__6881\,
            in2 => \N__6843\,
            in3 => \N__6429\,
            lcout => \U409_TICK.COUNTER50Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6772\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_0_LC_15_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__6879\,
            in1 => \N__6905\,
            in2 => \N__6837\,
            in3 => \N__6409\,
            lcout => \U409_TICK.COUNTER50Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6772\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_1_LC_15_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__6410\,
            in1 => \_gnd_net_\,
            in2 => \N__6663\,
            in3 => \_gnd_net_\,
            lcout => \U409_TICK.COUNTER50Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6772\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNID6CP_3_LC_15_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__6699\,
            in1 => \N__6423\,
            in2 => \_gnd_net_\,
            in3 => \N__6408\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK503_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNITU182_10_LC_15_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__6630\,
            in1 => \N__6390\,
            in2 => \N__6378\,
            in3 => \N__6375\,
            lcout => \U409_TICK.TICK503_14\,
            ltout => \U409_TICK.TICK503_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_5_LC_15_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6880\,
            in1 => \N__6839\,
            in2 => \N__6708\,
            in3 => \N__6705\,
            lcout => \U409_TICK.COUNTER50Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6772\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIUHF01_16_LC_15_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6687\,
            in1 => \N__6675\,
            in2 => \N__6662\,
            in3 => \N__6641\,
            lcout => \U409_TICK.TICK503_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK50_LC_15_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__6882\,
            in1 => \N__6614\,
            in2 => \N__6838\,
            in3 => \N__6907\,
            lcout => \TICK50_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6772\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_9_LC_15_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__6878\,
            in1 => \N__6603\,
            in2 => \N__6836\,
            in3 => \N__6912\,
            lcout => \U409_TICK.COUNTER50Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6774\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIH14V_11_LC_15_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6513\,
            in1 => \N__6594\,
            in2 => \N__6582\,
            in3 => \N__6558\,
            lcout => \U409_TICK.TICK503_9\,
            ltout => \U409_TICK.TICK503_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_13_LC_15_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6909\,
            in1 => \N__6875\,
            in2 => \N__6567\,
            in3 => \N__6564\,
            lcout => \U409_TICK.COUNTER50Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6774\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNII24V_14_LC_15_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__6924\,
            in1 => \N__6546\,
            in2 => \N__6792\,
            in3 => \N__6534\,
            lcout => \U409_TICK.TICK503_10\,
            ltout => \U409_TICK.TICK503_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_11_LC_15_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6908\,
            in1 => \N__6819\,
            in2 => \N__6522\,
            in3 => \N__6519\,
            lcout => \U409_TICK.COUNTER50Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6774\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_15_LC_15_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6877\,
            in1 => \N__6911\,
            in2 => \N__6835\,
            in3 => \N__6930\,
            lcout => \U409_TICK.COUNTER50Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6774\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_14_LC_15_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__6910\,
            in1 => \N__6876\,
            in2 => \N__6852\,
            in3 => \N__6820\,
            lcout => \U409_TICK.COUNTER50Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6774\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_iobuf_RNO_LC_19_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6744\,
            lcout => \N_475_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

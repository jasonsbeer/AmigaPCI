-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 25 2025 20:17:12

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    A : in std_logic_vector(20 downto 0);
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    DBRn : in std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__12003\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11714\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \N_882_i\ : std_logic;
signal \U712_REG_SM.N_71_i_cascade_\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \U712_REG_SM.N_265_cascade_\ : std_logic;
signal \ASn_c\ : std_logic;
signal \INVU712_REG_SM.STATE_COUNTER_9C_net\ : std_logic;
signal \REGENn_c\ : std_logic;
signal \INVU712_REG_SM.REGENnC_net\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_REG_SM.N_330_cascade_\ : std_logic;
signal \INVU712_REG_SM.LDSnC_net\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_REG_SM.N_295_cascade_\ : std_logic;
signal \U712_REG_SM.LDSn_6_iv_i_0_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_REG_SM.N_332\ : std_logic;
signal \U712_REG_SM.UDSn_6_iv_i_0_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTER_RNI7KTS1Z0Z_9\ : std_logic;
signal \UDSn_c\ : std_logic;
signal \U712_REG_SM.N_266\ : std_logic;
signal \U712_REG_SM.STATE_COUNTER_srsts_i_i_i_a3_3_0_cascade_\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.CYCLE_RUNZ0\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \INVU712_REG_SM.UDSnC_net\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_9\ : std_logic;
signal \U712_REG_SM.N_71_i\ : std_logic;
signal \REG_CPU_CYCLE\ : std_logic;
signal \INVU712_REG_SM.LATCH_REGC_net\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \INVU712_REG_SM.C3_SYNC_0C_net\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.N_241_cascade_\ : std_logic;
signal \U712_BYTE_ENABLE.N_276\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0Z0Z_0_cascade_\ : std_logic;
signal \N_47_i\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \A_c_14\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5_cascade_\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.N_361_cascade_\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \U712_CHIP_RAM.N_452\ : std_logic;
signal \U712_CHIP_RAM.N_452_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0\ : std_logic;
signal \LDSn_c\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_309\ : std_logic;
signal \U712_REG_SM.STATE_COUNTER_srsts_i_i_i_a3_2_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_5\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_7\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_3\ : std_logic;
signal \U712_REG_SM.un18_0_i_0_0_1_cascade_\ : std_logic;
signal \INVU712_REG_SM.STATE_COUNTER_5C_net\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_8\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_4\ : std_logic;
signal \U712_REG_SM.N_442_cascade_\ : std_logic;
signal \U712_REG_SM.REG_CPU_CYCLE_e_1\ : std_logic;
signal \U712_REG_SM.N_84\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_447\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_6\ : std_logic;
signal \U712_REG_SM.N_288\ : std_logic;
signal \LATCH_REG\ : std_logic;
signal \LATCH_CLK_0_i\ : std_logic;
signal \A_c_8\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\ : std_logic;
signal \A_c_13\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i\ : std_logic;
signal \A_c_11\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_325_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_301\ : std_logic;
signal \U712_CHIP_RAM.N_392_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_449\ : std_logic;
signal \U712_CHIP_RAM.N_376_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_45_i_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_324_2\ : std_logic;
signal \U712_CHIP_RAM.N_324_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_450\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNIVIFVCZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.N_252\ : std_logic;
signal \U712_CHIP_RAM.N_252_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_365_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0\ : std_logic;
signal \RnW_c\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\ : std_logic;
signal \LATCH_RAM\ : std_logic;
signal \U712_REG_SM.N_265\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_2\ : std_logic;
signal \U712_REG_SM.DBR_SYNCZ0Z_1\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \U712_REG_SM.DBR_SYNCZ0Z_0\ : std_logic;
signal \INVU712_REG_SM.STATE_COUNTER_2C_net\ : std_logic;
signal \REG_WRITE_CYCLE\ : std_logic;
signal \N_289\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lt7\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.N_324\ : std_logic;
signal \U712_CHIP_RAM.N_456_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.N_363\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.N_384_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_448_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_255\ : std_logic;
signal \U712_CHIP_RAM.N_255_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_269\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_444\ : std_logic;
signal \U712_CHIP_RAM.N_392\ : std_logic;
signal \U712_CHIP_RAM.N_444_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.N_334\ : std_logic;
signal \U712_CHIP_RAM.N_334_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_448\ : std_logic;
signal \U712_CHIP_RAM.N_323\ : std_logic;
signal \U712_CHIP_RAM.N_323_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un3_DMA_CYCLE_START\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \N_46_i\ : std_logic;
signal \U712_BYTE_ENABLE.UUBE_cascade_\ : std_logic;
signal \N_48_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_278\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0Z0Z_0\ : std_logic;
signal \N_49_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_277\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_2_0\ : std_logic;
signal \U712_CHIP_RAM.N_325_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_365_1\ : std_logic;
signal \U712_CHIP_RAM.N_294\ : std_logic;
signal \DMA_CYCLE\ : std_logic;
signal \U712_CHIP_RAM.N_305_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_388\ : std_logic;
signal \U712_CHIP_RAM.N_45_i\ : std_logic;
signal \U712_CHIP_RAM.N_346_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_180_i_2\ : std_logic;
signal \U712_CHIP_RAM.N_407\ : std_logic;
signal \U712_CHIP_RAM.N_407_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_400\ : std_logic;
signal \WRITE_CYCLE\ : std_logic;
signal \U712_CHIP_RAM.N_257_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.N_396_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_436\ : std_logic;
signal \U712_CHIP_RAM.N_436_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_257\ : std_logic;
signal \U712_CHIP_RAM.N_357\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_396\ : std_logic;
signal \U712_CHIP_RAM.N_384\ : std_logic;
signal \U712_CHIP_RAM.N_351\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_117\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_63_i_a2_0_0_a2_0_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.N_274_i_0_0_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_274_i_0_en_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_274_i_0_en_0\ : std_logic;
signal \U712_CHIP_RAM.N_456\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \U712_CHIP_RAM.N_202\ : std_logic;
signal \U712_CHIP_RAM.N_359\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \CLK40_PLL\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \U712_CYCLE_TERM.N_8\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \CPU_TACK\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \REG_CYCLE\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \CLK40_PLL_g\ : std_logic;
signal \CLK40_PLL_iso_i\ : std_logic;
signal \U712_BYTE_ENABLE_UUBE_i\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\ : std_logic;
signal \N_276_i\ : std_logic;
signal \N_278_i\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \A_c_1\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \N_277_i\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \RASn_c\ : std_logic;
signal \CASn_c\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_0\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \CPU_CYCLE\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z20\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A20C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL\,
            REFERENCECLK => \N__4061\,
            RESETB => \N__6878\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12003\,
            DIN => \N__12002\,
            DOUT => \N__12001\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12003\,
            PADOUT => \N__12002\,
            PADIN => \N__12001\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6959\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11994\,
            DIN => \N__11993\,
            DOUT => \N__11992\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11994\,
            PADOUT => \N__11993\,
            PADIN => \N__11992\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11985\,
            DIN => \N__11984\,
            DOUT => \N__11983\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11985\,
            PADOUT => \N__11984\,
            PADIN => \N__11983\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8897\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11976\,
            DIN => \N__11975\,
            DOUT => \N__11974\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11976\,
            PADOUT => \N__11975\,
            PADIN => \N__11974\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5867\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11967\,
            DIN => \N__11966\,
            DOUT => \N__11965\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11967\,
            PADOUT => \N__11966\,
            PADIN => \N__11965\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11958\,
            DIN => \N__11957\,
            DOUT => \N__11956\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11958\,
            PADOUT => \N__11957\,
            PADIN => \N__11956\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11949\,
            DIN => \N__11948\,
            DOUT => \N__11947\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11949\,
            PADOUT => \N__11948\,
            PADIN => \N__11947\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11940\,
            DIN => \N__11939\,
            DOUT => \N__11938\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11940\,
            PADOUT => \N__11939\,
            PADIN => \N__11938\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11931\,
            DIN => \N__11930\,
            DOUT => \N__11929\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11931\,
            PADOUT => \N__11930\,
            PADIN => \N__11929\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11922\,
            DIN => \N__11921\,
            DOUT => \N__11920\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11922\,
            PADOUT => \N__11921\,
            PADIN => \N__11920\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11913\,
            DIN => \N__11912\,
            DOUT => \N__11911\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11913\,
            PADOUT => \N__11912\,
            PADIN => \N__11911\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6857\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11904\,
            DIN => \N__11903\,
            DOUT => \N__11902\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11904\,
            PADOUT => \N__11903\,
            PADIN => \N__11902\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8780\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11895\,
            DIN => \N__11894\,
            DOUT => \N__11893\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11895\,
            PADOUT => \N__11894\,
            PADIN => \N__11893\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11886\,
            DIN => \N__11885\,
            DOUT => \N__11884\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11886\,
            PADOUT => \N__11885\,
            PADIN => \N__11884\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11877\,
            DIN => \N__11876\,
            DOUT => \N__11875\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11877\,
            PADOUT => \N__11876\,
            PADIN => \N__11875\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11868\,
            DIN => \N__11867\,
            DOUT => \N__11866\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11868\,
            PADOUT => \N__11867\,
            PADIN => \N__11866\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4139\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11859\,
            DIN => \N__11858\,
            DOUT => \N__11857\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11859\,
            PADOUT => \N__11858\,
            PADIN => \N__11857\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11850\,
            DIN => \N__11849\,
            DOUT => \N__11848\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11850\,
            PADOUT => \N__11849\,
            PADIN => \N__11848\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11841\,
            DIN => \N__11840\,
            DOUT => \N__11839\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11841\,
            PADOUT => \N__11840\,
            PADIN => \N__11839\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9947\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11832\,
            DIN => \N__11831\,
            DOUT => \N__11830\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11832\,
            PADOUT => \N__11831\,
            PADIN => \N__11830\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11823\,
            DIN => \N__11822\,
            DOUT => \N__11821\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11823\,
            PADOUT => \N__11822\,
            PADIN => \N__11821\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8936\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11814\,
            DIN => \N__11813\,
            DOUT => \N__11812\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11814\,
            PADOUT => \N__11813\,
            PADIN => \N__11812\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11805\,
            DIN => \N__11804\,
            DOUT => \N__11803\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11805\,
            PADOUT => \N__11804\,
            PADIN => \N__11803\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9314\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11796\,
            DIN => \N__11795\,
            DOUT => \N__11794\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11796\,
            PADOUT => \N__11795\,
            PADIN => \N__11794\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11787\,
            DIN => \N__11786\,
            DOUT => \N__11785\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11787\,
            PADOUT => \N__11786\,
            PADIN => \N__11785\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11778\,
            DIN => \N__11777\,
            DOUT => \N__11776\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11778\,
            PADOUT => \N__11777\,
            PADIN => \N__11776\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11769\,
            DIN => \N__11768\,
            DOUT => \N__11767\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11769\,
            PADOUT => \N__11768\,
            PADIN => \N__11767\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11760\,
            DIN => \N__11759\,
            DOUT => \N__11758\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11760\,
            PADOUT => \N__11759\,
            PADIN => \N__11758\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11751\,
            DIN => \N__11750\,
            DOUT => \N__11749\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11751\,
            PADOUT => \N__11750\,
            PADIN => \N__11749\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5863\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11742\,
            DIN => \N__11741\,
            DOUT => \N__11740\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11742\,
            PADOUT => \N__11741\,
            PADIN => \N__11740\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11733\,
            DIN => \N__11732\,
            DOUT => \N__11731\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11733\,
            PADOUT => \N__11732\,
            PADIN => \N__11731\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11724\,
            DIN => \N__11723\,
            DOUT => \N__11722\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11724\,
            PADOUT => \N__11723\,
            PADIN => \N__11722\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11715\,
            DIN => \N__11714\,
            DOUT => \N__11713\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11715\,
            PADOUT => \N__11714\,
            PADIN => \N__11713\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11706\,
            DIN => \N__11705\,
            DOUT => \N__11704\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11706\,
            PADOUT => \N__11705\,
            PADIN => \N__11704\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11697\,
            DIN => \N__11696\,
            DOUT => \N__11695\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11697\,
            PADOUT => \N__11696\,
            PADIN => \N__11695\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8918\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11688\,
            DIN => \N__11687\,
            DOUT => \N__11686\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11688\,
            PADOUT => \N__11687\,
            PADIN => \N__11686\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4733\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11679\,
            DIN => \N__11678\,
            DOUT => \N__11677\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11679\,
            PADOUT => \N__11678\,
            PADIN => \N__11677\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8827\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11670\,
            DIN => \N__11669\,
            DOUT => \N__11668\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11670\,
            PADOUT => \N__11669\,
            PADIN => \N__11668\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4115\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11661\,
            DIN => \N__11660\,
            DOUT => \N__11659\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11661\,
            PADOUT => \N__11660\,
            PADIN => \N__11659\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11652\,
            DIN => \N__11651\,
            DOUT => \N__11650\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11652\,
            PADOUT => \N__11651\,
            PADIN => \N__11650\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4196\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11643\,
            DIN => \N__11642\,
            DOUT => \N__11641\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11643\,
            PADOUT => \N__11642\,
            PADIN => \N__11641\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6803\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11634\,
            DIN => \N__11633\,
            DOUT => \N__11632\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11634\,
            PADOUT => \N__11633\,
            PADIN => \N__11632\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11625\,
            DIN => \N__11624\,
            DOUT => \N__11623\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11625\,
            PADOUT => \N__11624\,
            PADIN => \N__11623\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11616\,
            DIN => \N__11615\,
            DOUT => \N__11614\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11616\,
            PADOUT => \N__11615\,
            PADIN => \N__11614\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11607\,
            DIN => \N__11606\,
            DOUT => \N__11605\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11607\,
            PADOUT => \N__11606\,
            PADIN => \N__11605\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11598\,
            DIN => \N__11597\,
            DOUT => \N__11596\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11598\,
            PADOUT => \N__11597\,
            PADIN => \N__11596\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10172\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11589\,
            DIN => \N__11588\,
            DOUT => \N__11587\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11589\,
            PADOUT => \N__11588\,
            PADIN => \N__11587\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11580\,
            DIN => \N__11579\,
            DOUT => \N__11578\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11580\,
            PADOUT => \N__11579\,
            PADIN => \N__11578\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8820\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11571\,
            DIN => \N__11570\,
            DOUT => \N__11569\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11571\,
            PADOUT => \N__11570\,
            PADIN => \N__11569\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6830\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11562\,
            DIN => \N__11561\,
            DOUT => \N__11560\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11562\,
            PADOUT => \N__11561\,
            PADIN => \N__11560\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7976\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11553\,
            DIN => \N__11552\,
            DOUT => \N__11551\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11553\,
            PADOUT => \N__11552\,
            PADIN => \N__11551\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4622\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11544\,
            DIN => \N__11543\,
            DOUT => \N__11542\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11544\,
            PADOUT => \N__11543\,
            PADIN => \N__11542\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6734\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11535\,
            DIN => \N__11534\,
            DOUT => \N__11533\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11535\,
            PADOUT => \N__11534\,
            PADIN => \N__11533\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4166\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11526\,
            DIN => \N__11525\,
            DOUT => \N__11524\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11526\,
            PADOUT => \N__11525\,
            PADIN => \N__11524\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11517\,
            DIN => \N__11516\,
            DOUT => \N__11515\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11517\,
            PADOUT => \N__11516\,
            PADIN => \N__11515\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11508\,
            DIN => \N__11507\,
            DOUT => \N__11506\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11508\,
            PADOUT => \N__11507\,
            PADIN => \N__11506\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6986\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11499\,
            DIN => \N__11498\,
            DOUT => \N__11497\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11499\,
            PADOUT => \N__11498\,
            PADIN => \N__11497\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10340\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11490\,
            DIN => \N__11489\,
            DOUT => \N__11488\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11490\,
            PADOUT => \N__11489\,
            PADIN => \N__11488\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6233\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11481\,
            DIN => \N__11480\,
            DOUT => \N__11479\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11481\,
            PADOUT => \N__11480\,
            PADIN => \N__11479\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6692\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11472\,
            DIN => \N__11471\,
            DOUT => \N__11470\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11472\,
            PADOUT => \N__11471\,
            PADIN => \N__11470\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11463\,
            DIN => \N__11462\,
            DOUT => \N__11461\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11463\,
            PADOUT => \N__11462\,
            PADIN => \N__11461\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11454\,
            DIN => \N__11453\,
            DOUT => \N__11452\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11454\,
            PADOUT => \N__11453\,
            PADIN => \N__11452\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11445\,
            DIN => \N__11444\,
            DOUT => \N__11443\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11445\,
            PADOUT => \N__11444\,
            PADIN => \N__11443\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11436\,
            DIN => \N__11435\,
            DOUT => \N__11434\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11436\,
            PADOUT => \N__11435\,
            PADIN => \N__11434\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5315\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11427\,
            DIN => \N__11426\,
            DOUT => \N__11425\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11427\,
            PADOUT => \N__11426\,
            PADIN => \N__11425\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9299\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11418\,
            DIN => \N__11417\,
            DOUT => \N__11416\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11418\,
            PADOUT => \N__11417\,
            PADIN => \N__11416\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11409\,
            DIN => \N__11408\,
            DOUT => \N__11407\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11409\,
            PADOUT => \N__11408\,
            PADIN => \N__11407\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7031\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11400\,
            DIN => \N__11399\,
            DOUT => \N__11398\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11400\,
            PADOUT => \N__11399\,
            PADIN => \N__11398\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4100\,
            DIN0 => OPEN,
            DOUT0 => \N__4361\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11391\,
            DIN => \N__11390\,
            DOUT => \N__11389\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11391\,
            PADOUT => \N__11390\,
            PADIN => \N__11389\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6713\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11382\,
            DIN => \N__11381\,
            DOUT => \N__11380\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11382\,
            PADOUT => \N__11381\,
            PADIN => \N__11380\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11373\,
            DIN => \N__11372\,
            DOUT => \N__11371\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11373\,
            PADOUT => \N__11372\,
            PADIN => \N__11371\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11364\,
            DIN => \N__11363\,
            DOUT => \N__11362\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11364\,
            PADOUT => \N__11363\,
            PADIN => \N__11362\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8717\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11355\,
            DIN => \N__11354\,
            DOUT => \N__11353\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11355\,
            PADOUT => \N__11354\,
            PADIN => \N__11353\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11346\,
            DIN => \N__11345\,
            DOUT => \N__11344\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11346\,
            PADOUT => \N__11345\,
            PADIN => \N__11344\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11337\,
            DIN => \N__11336\,
            DOUT => \N__11335\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11337\,
            PADOUT => \N__11336\,
            PADIN => \N__11335\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11328\,
            DIN => \N__11327\,
            DOUT => \N__11326\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11328\,
            PADOUT => \N__11327\,
            PADIN => \N__11326\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11319\,
            DIN => \N__11318\,
            DOUT => \N__11317\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11319\,
            PADOUT => \N__11318\,
            PADIN => \N__11317\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5342\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11310\,
            DIN => \N__11309\,
            DOUT => \N__11308\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11310\,
            PADOUT => \N__11309\,
            PADIN => \N__11308\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4283\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11301\,
            DIN => \N__11300\,
            DOUT => \N__11299\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11301\,
            PADOUT => \N__11300\,
            PADIN => \N__11299\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8954\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11292\,
            DIN => \N__11291\,
            DOUT => \N__11290\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11292\,
            PADOUT => \N__11291\,
            PADIN => \N__11290\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5702\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11283\,
            DIN => \N__11282\,
            DOUT => \N__11281\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11283\,
            PADOUT => \N__11282\,
            PADIN => \N__11281\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11274\,
            DIN => \N__11273\,
            DOUT => \N__11272\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11274\,
            PADOUT => \N__11273\,
            PADIN => \N__11272\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11265\,
            DIN => \N__11264\,
            DOUT => \N__11263\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11265\,
            PADOUT => \N__11264\,
            PADIN => \N__11263\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6773\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11256\,
            DIN => \N__11255\,
            DOUT => \N__11254\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11256\,
            PADOUT => \N__11255\,
            PADIN => \N__11254\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11247\,
            DIN => \N__11246\,
            DOUT => \N__11245\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11247\,
            PADOUT => \N__11246\,
            PADIN => \N__11245\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11238\,
            DIN => \N__11237\,
            DOUT => \N__11236\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11238\,
            PADOUT => \N__11237\,
            PADIN => \N__11236\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4943\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11229\,
            DIN => \N__11228\,
            DOUT => \N__11227\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11229\,
            PADOUT => \N__11228\,
            PADIN => \N__11227\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4907\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11220\,
            DIN => \N__11219\,
            DOUT => \N__11218\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11220\,
            PADOUT => \N__11219\,
            PADIN => \N__11218\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8831\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11211\,
            DIN => \N__11210\,
            DOUT => \N__11209\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11211\,
            PADOUT => \N__11210\,
            PADIN => \N__11209\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2739\ : CascadeMux
    port map (
            O => \N__11192\,
            I => \N__11189\
        );

    \I__2738\ : InMux
    port map (
            O => \N__11189\,
            I => \N__11185\
        );

    \I__2737\ : CascadeMux
    port map (
            O => \N__11188\,
            I => \N__11178\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__11185\,
            I => \N__11174\
        );

    \I__2735\ : InMux
    port map (
            O => \N__11184\,
            I => \N__11169\
        );

    \I__2734\ : InMux
    port map (
            O => \N__11183\,
            I => \N__11169\
        );

    \I__2733\ : InMux
    port map (
            O => \N__11182\,
            I => \N__11164\
        );

    \I__2732\ : InMux
    port map (
            O => \N__11181\,
            I => \N__11164\
        );

    \I__2731\ : InMux
    port map (
            O => \N__11178\,
            I => \N__11158\
        );

    \I__2730\ : InMux
    port map (
            O => \N__11177\,
            I => \N__11158\
        );

    \I__2729\ : Span4Mux_v
    port map (
            O => \N__11174\,
            I => \N__11147\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__11169\,
            I => \N__11142\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__11164\,
            I => \N__11142\
        );

    \I__2726\ : InMux
    port map (
            O => \N__11163\,
            I => \N__11139\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__11158\,
            I => \N__11136\
        );

    \I__2724\ : InMux
    port map (
            O => \N__11157\,
            I => \N__11133\
        );

    \I__2723\ : InMux
    port map (
            O => \N__11156\,
            I => \N__11126\
        );

    \I__2722\ : InMux
    port map (
            O => \N__11155\,
            I => \N__11126\
        );

    \I__2721\ : InMux
    port map (
            O => \N__11154\,
            I => \N__11126\
        );

    \I__2720\ : InMux
    port map (
            O => \N__11153\,
            I => \N__11123\
        );

    \I__2719\ : InMux
    port map (
            O => \N__11152\,
            I => \N__11120\
        );

    \I__2718\ : InMux
    port map (
            O => \N__11151\,
            I => \N__11117\
        );

    \I__2717\ : InMux
    port map (
            O => \N__11150\,
            I => \N__11114\
        );

    \I__2716\ : Span4Mux_h
    port map (
            O => \N__11147\,
            I => \N__11105\
        );

    \I__2715\ : Span4Mux_v
    port map (
            O => \N__11142\,
            I => \N__11105\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__11139\,
            I => \N__11105\
        );

    \I__2713\ : Span4Mux_h
    port map (
            O => \N__11136\,
            I => \N__11100\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__11133\,
            I => \N__11100\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__11126\,
            I => \N__11088\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__11123\,
            I => \N__11088\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__11120\,
            I => \N__11088\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__11117\,
            I => \N__11088\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__11114\,
            I => \N__11088\
        );

    \I__2706\ : InMux
    port map (
            O => \N__11113\,
            I => \N__11084\
        );

    \I__2705\ : InMux
    port map (
            O => \N__11112\,
            I => \N__11080\
        );

    \I__2704\ : Span4Mux_h
    port map (
            O => \N__11105\,
            I => \N__11075\
        );

    \I__2703\ : Span4Mux_v
    port map (
            O => \N__11100\,
            I => \N__11075\
        );

    \I__2702\ : InMux
    port map (
            O => \N__11099\,
            I => \N__11072\
        );

    \I__2701\ : Span4Mux_v
    port map (
            O => \N__11088\,
            I => \N__11069\
        );

    \I__2700\ : InMux
    port map (
            O => \N__11087\,
            I => \N__11066\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__11084\,
            I => \N__11063\
        );

    \I__2698\ : InMux
    port map (
            O => \N__11083\,
            I => \N__11060\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__11080\,
            I => \N__11057\
        );

    \I__2696\ : Sp12to4
    port map (
            O => \N__11075\,
            I => \N__11048\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__11072\,
            I => \N__11048\
        );

    \I__2694\ : Sp12to4
    port map (
            O => \N__11069\,
            I => \N__11048\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__11066\,
            I => \N__11048\
        );

    \I__2692\ : Sp12to4
    port map (
            O => \N__11063\,
            I => \N__11043\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__11060\,
            I => \N__11043\
        );

    \I__2690\ : Span12Mux_h
    port map (
            O => \N__11057\,
            I => \N__11040\
        );

    \I__2689\ : Span12Mux_h
    port map (
            O => \N__11048\,
            I => \N__11037\
        );

    \I__2688\ : Span12Mux_v
    port map (
            O => \N__11043\,
            I => \N__11034\
        );

    \I__2687\ : Span12Mux_v
    port map (
            O => \N__11040\,
            I => \N__11031\
        );

    \I__2686\ : Span12Mux_v
    port map (
            O => \N__11037\,
            I => \N__11026\
        );

    \I__2685\ : Span12Mux_h
    port map (
            O => \N__11034\,
            I => \N__11026\
        );

    \I__2684\ : Odrv12
    port map (
            O => \N__11031\,
            I => \AGNUS_REV_c\
        );

    \I__2683\ : Odrv12
    port map (
            O => \N__11026\,
            I => \AGNUS_REV_c\
        );

    \I__2682\ : InMux
    port map (
            O => \N__11021\,
            I => \N__11017\
        );

    \I__2681\ : InMux
    port map (
            O => \N__11020\,
            I => \N__11014\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__11017\,
            I => \N__11009\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__11014\,
            I => \N__11009\
        );

    \I__2678\ : Sp12to4
    port map (
            O => \N__11009\,
            I => \N__11006\
        );

    \I__2677\ : Span12Mux_v
    port map (
            O => \N__11006\,
            I => \N__11003\
        );

    \I__2676\ : Span12Mux_h
    port map (
            O => \N__11003\,
            I => \N__11000\
        );

    \I__2675\ : Odrv12
    port map (
            O => \N__11000\,
            I => \DRA_c_0\
        );

    \I__2674\ : InMux
    port map (
            O => \N__10997\,
            I => \N__10992\
        );

    \I__2673\ : InMux
    port map (
            O => \N__10996\,
            I => \N__10988\
        );

    \I__2672\ : InMux
    port map (
            O => \N__10995\,
            I => \N__10985\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__10992\,
            I => \N__10982\
        );

    \I__2670\ : InMux
    port map (
            O => \N__10991\,
            I => \N__10979\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__10988\,
            I => \N__10972\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__10985\,
            I => \N__10972\
        );

    \I__2667\ : Span4Mux_v
    port map (
            O => \N__10982\,
            I => \N__10972\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__10979\,
            I => \N__10969\
        );

    \I__2665\ : Sp12to4
    port map (
            O => \N__10972\,
            I => \N__10966\
        );

    \I__2664\ : Span4Mux_h
    port map (
            O => \N__10969\,
            I => \N__10963\
        );

    \I__2663\ : Span12Mux_h
    port map (
            O => \N__10966\,
            I => \N__10958\
        );

    \I__2662\ : Sp12to4
    port map (
            O => \N__10963\,
            I => \N__10958\
        );

    \I__2661\ : Span12Mux_v
    port map (
            O => \N__10958\,
            I => \N__10955\
        );

    \I__2660\ : Odrv12
    port map (
            O => \N__10955\,
            I => \DRA_c_1\
        );

    \I__2659\ : InMux
    port map (
            O => \N__10952\,
            I => \N__10949\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__10949\,
            I => \N__10946\
        );

    \I__2657\ : Odrv4
    port map (
            O => \N__10946\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2656\ : ClkMux
    port map (
            O => \N__10943\,
            I => \N__10925\
        );

    \I__2655\ : ClkMux
    port map (
            O => \N__10942\,
            I => \N__10925\
        );

    \I__2654\ : ClkMux
    port map (
            O => \N__10941\,
            I => \N__10925\
        );

    \I__2653\ : ClkMux
    port map (
            O => \N__10940\,
            I => \N__10925\
        );

    \I__2652\ : ClkMux
    port map (
            O => \N__10939\,
            I => \N__10925\
        );

    \I__2651\ : ClkMux
    port map (
            O => \N__10938\,
            I => \N__10925\
        );

    \I__2650\ : GlobalMux
    port map (
            O => \N__10925\,
            I => \N__10922\
        );

    \I__2649\ : gio2CtrlBuf
    port map (
            O => \N__10922\,
            I => \C3_c_g\
        );

    \I__2648\ : CEMux
    port map (
            O => \N__10919\,
            I => \N__10880\
        );

    \I__2647\ : CEMux
    port map (
            O => \N__10918\,
            I => \N__10880\
        );

    \I__2646\ : CEMux
    port map (
            O => \N__10917\,
            I => \N__10880\
        );

    \I__2645\ : CEMux
    port map (
            O => \N__10916\,
            I => \N__10880\
        );

    \I__2644\ : CEMux
    port map (
            O => \N__10915\,
            I => \N__10880\
        );

    \I__2643\ : CEMux
    port map (
            O => \N__10914\,
            I => \N__10880\
        );

    \I__2642\ : CEMux
    port map (
            O => \N__10913\,
            I => \N__10880\
        );

    \I__2641\ : CEMux
    port map (
            O => \N__10912\,
            I => \N__10880\
        );

    \I__2640\ : CEMux
    port map (
            O => \N__10911\,
            I => \N__10880\
        );

    \I__2639\ : CEMux
    port map (
            O => \N__10910\,
            I => \N__10880\
        );

    \I__2638\ : CEMux
    port map (
            O => \N__10909\,
            I => \N__10880\
        );

    \I__2637\ : CEMux
    port map (
            O => \N__10908\,
            I => \N__10880\
        );

    \I__2636\ : CEMux
    port map (
            O => \N__10907\,
            I => \N__10880\
        );

    \I__2635\ : GlobalMux
    port map (
            O => \N__10880\,
            I => \N__10877\
        );

    \I__2634\ : gio2CtrlBuf
    port map (
            O => \N__10877\,
            I => \DBRn_c_i_0_g\
        );

    \I__2633\ : InMux
    port map (
            O => \N__10874\,
            I => \N__10867\
        );

    \I__2632\ : InMux
    port map (
            O => \N__10873\,
            I => \N__10864\
        );

    \I__2631\ : InMux
    port map (
            O => \N__10872\,
            I => \N__10861\
        );

    \I__2630\ : InMux
    port map (
            O => \N__10871\,
            I => \N__10858\
        );

    \I__2629\ : InMux
    port map (
            O => \N__10870\,
            I => \N__10855\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__10867\,
            I => \N__10841\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__10864\,
            I => \N__10833\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__10861\,
            I => \N__10825\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__10858\,
            I => \N__10816\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__10855\,
            I => \N__10803\
        );

    \I__2623\ : SRMux
    port map (
            O => \N__10854\,
            I => \N__10703\
        );

    \I__2622\ : SRMux
    port map (
            O => \N__10853\,
            I => \N__10703\
        );

    \I__2621\ : SRMux
    port map (
            O => \N__10852\,
            I => \N__10703\
        );

    \I__2620\ : SRMux
    port map (
            O => \N__10851\,
            I => \N__10703\
        );

    \I__2619\ : SRMux
    port map (
            O => \N__10850\,
            I => \N__10703\
        );

    \I__2618\ : SRMux
    port map (
            O => \N__10849\,
            I => \N__10703\
        );

    \I__2617\ : SRMux
    port map (
            O => \N__10848\,
            I => \N__10703\
        );

    \I__2616\ : SRMux
    port map (
            O => \N__10847\,
            I => \N__10703\
        );

    \I__2615\ : SRMux
    port map (
            O => \N__10846\,
            I => \N__10703\
        );

    \I__2614\ : SRMux
    port map (
            O => \N__10845\,
            I => \N__10703\
        );

    \I__2613\ : SRMux
    port map (
            O => \N__10844\,
            I => \N__10703\
        );

    \I__2612\ : Glb2LocalMux
    port map (
            O => \N__10841\,
            I => \N__10703\
        );

    \I__2611\ : SRMux
    port map (
            O => \N__10840\,
            I => \N__10703\
        );

    \I__2610\ : SRMux
    port map (
            O => \N__10839\,
            I => \N__10703\
        );

    \I__2609\ : SRMux
    port map (
            O => \N__10838\,
            I => \N__10703\
        );

    \I__2608\ : SRMux
    port map (
            O => \N__10837\,
            I => \N__10703\
        );

    \I__2607\ : SRMux
    port map (
            O => \N__10836\,
            I => \N__10703\
        );

    \I__2606\ : Glb2LocalMux
    port map (
            O => \N__10833\,
            I => \N__10703\
        );

    \I__2605\ : SRMux
    port map (
            O => \N__10832\,
            I => \N__10703\
        );

    \I__2604\ : SRMux
    port map (
            O => \N__10831\,
            I => \N__10703\
        );

    \I__2603\ : SRMux
    port map (
            O => \N__10830\,
            I => \N__10703\
        );

    \I__2602\ : SRMux
    port map (
            O => \N__10829\,
            I => \N__10703\
        );

    \I__2601\ : SRMux
    port map (
            O => \N__10828\,
            I => \N__10703\
        );

    \I__2600\ : Glb2LocalMux
    port map (
            O => \N__10825\,
            I => \N__10703\
        );

    \I__2599\ : SRMux
    port map (
            O => \N__10824\,
            I => \N__10703\
        );

    \I__2598\ : SRMux
    port map (
            O => \N__10823\,
            I => \N__10703\
        );

    \I__2597\ : SRMux
    port map (
            O => \N__10822\,
            I => \N__10703\
        );

    \I__2596\ : SRMux
    port map (
            O => \N__10821\,
            I => \N__10703\
        );

    \I__2595\ : SRMux
    port map (
            O => \N__10820\,
            I => \N__10703\
        );

    \I__2594\ : SRMux
    port map (
            O => \N__10819\,
            I => \N__10703\
        );

    \I__2593\ : Glb2LocalMux
    port map (
            O => \N__10816\,
            I => \N__10703\
        );

    \I__2592\ : SRMux
    port map (
            O => \N__10815\,
            I => \N__10703\
        );

    \I__2591\ : SRMux
    port map (
            O => \N__10814\,
            I => \N__10703\
        );

    \I__2590\ : SRMux
    port map (
            O => \N__10813\,
            I => \N__10703\
        );

    \I__2589\ : SRMux
    port map (
            O => \N__10812\,
            I => \N__10703\
        );

    \I__2588\ : SRMux
    port map (
            O => \N__10811\,
            I => \N__10703\
        );

    \I__2587\ : SRMux
    port map (
            O => \N__10810\,
            I => \N__10703\
        );

    \I__2586\ : SRMux
    port map (
            O => \N__10809\,
            I => \N__10703\
        );

    \I__2585\ : SRMux
    port map (
            O => \N__10808\,
            I => \N__10703\
        );

    \I__2584\ : SRMux
    port map (
            O => \N__10807\,
            I => \N__10703\
        );

    \I__2583\ : SRMux
    port map (
            O => \N__10806\,
            I => \N__10703\
        );

    \I__2582\ : Glb2LocalMux
    port map (
            O => \N__10803\,
            I => \N__10703\
        );

    \I__2581\ : SRMux
    port map (
            O => \N__10802\,
            I => \N__10703\
        );

    \I__2580\ : SRMux
    port map (
            O => \N__10801\,
            I => \N__10703\
        );

    \I__2579\ : SRMux
    port map (
            O => \N__10800\,
            I => \N__10703\
        );

    \I__2578\ : SRMux
    port map (
            O => \N__10799\,
            I => \N__10703\
        );

    \I__2577\ : SRMux
    port map (
            O => \N__10798\,
            I => \N__10703\
        );

    \I__2576\ : GlobalMux
    port map (
            O => \N__10703\,
            I => \N__10700\
        );

    \I__2575\ : gio2CtrlBuf
    port map (
            O => \N__10700\,
            I => \RESETn_c_i_g\
        );

    \I__2574\ : CascadeMux
    port map (
            O => \N__10697\,
            I => \N__10694\
        );

    \I__2573\ : InMux
    port map (
            O => \N__10694\,
            I => \N__10690\
        );

    \I__2572\ : InMux
    port map (
            O => \N__10693\,
            I => \N__10687\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__10690\,
            I => \N__10680\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__10687\,
            I => \N__10680\
        );

    \I__2569\ : InMux
    port map (
            O => \N__10686\,
            I => \N__10677\
        );

    \I__2568\ : InMux
    port map (
            O => \N__10685\,
            I => \N__10674\
        );

    \I__2567\ : Sp12to4
    port map (
            O => \N__10680\,
            I => \N__10667\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__10677\,
            I => \N__10667\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__10674\,
            I => \N__10667\
        );

    \I__2564\ : Span12Mux_v
    port map (
            O => \N__10667\,
            I => \N__10664\
        );

    \I__2563\ : Span12Mux_h
    port map (
            O => \N__10664\,
            I => \N__10661\
        );

    \I__2562\ : Odrv12
    port map (
            O => \N__10661\,
            I => \DRA_c_6\
        );

    \I__2561\ : InMux
    port map (
            O => \N__10658\,
            I => \N__10655\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__10655\,
            I => \N__10652\
        );

    \I__2559\ : Span4Mux_h
    port map (
            O => \N__10652\,
            I => \N__10649\
        );

    \I__2558\ : Odrv4
    port map (
            O => \N__10649\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2557\ : InMux
    port map (
            O => \N__10646\,
            I => \N__10643\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__10643\,
            I => \N__10640\
        );

    \I__2555\ : Span4Mux_h
    port map (
            O => \N__10640\,
            I => \N__10636\
        );

    \I__2554\ : InMux
    port map (
            O => \N__10639\,
            I => \N__10633\
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__10636\,
            I => \DBRn_c_i\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__10633\,
            I => \DBRn_c_i\
        );

    \I__2551\ : InMux
    port map (
            O => \N__10628\,
            I => \N__10624\
        );

    \I__2550\ : InMux
    port map (
            O => \N__10627\,
            I => \N__10621\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__10624\,
            I => \N__10618\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__10621\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__2547\ : Odrv12
    port map (
            O => \N__10618\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__2546\ : InMux
    port map (
            O => \N__10613\,
            I => \N__10610\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__10610\,
            I => \N__10607\
        );

    \I__2544\ : Span4Mux_h
    port map (
            O => \N__10607\,
            I => \N__10604\
        );

    \I__2543\ : Odrv4
    port map (
            O => \N__10604\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2542\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10596\
        );

    \I__2541\ : InMux
    port map (
            O => \N__10600\,
            I => \N__10593\
        );

    \I__2540\ : InMux
    port map (
            O => \N__10599\,
            I => \N__10590\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__10596\,
            I => \N__10587\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__10593\,
            I => \N__10581\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__10590\,
            I => \N__10581\
        );

    \I__2536\ : Span4Mux_v
    port map (
            O => \N__10587\,
            I => \N__10578\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__10586\,
            I => \N__10575\
        );

    \I__2534\ : Span4Mux_h
    port map (
            O => \N__10581\,
            I => \N__10572\
        );

    \I__2533\ : Span4Mux_v
    port map (
            O => \N__10578\,
            I => \N__10569\
        );

    \I__2532\ : InMux
    port map (
            O => \N__10575\,
            I => \N__10566\
        );

    \I__2531\ : Span4Mux_v
    port map (
            O => \N__10572\,
            I => \N__10563\
        );

    \I__2530\ : Sp12to4
    port map (
            O => \N__10569\,
            I => \N__10558\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__10566\,
            I => \N__10558\
        );

    \I__2528\ : Sp12to4
    port map (
            O => \N__10563\,
            I => \N__10555\
        );

    \I__2527\ : Span12Mux_h
    port map (
            O => \N__10558\,
            I => \N__10552\
        );

    \I__2526\ : Span12Mux_v
    port map (
            O => \N__10555\,
            I => \N__10549\
        );

    \I__2525\ : Span12Mux_v
    port map (
            O => \N__10552\,
            I => \N__10546\
        );

    \I__2524\ : Odrv12
    port map (
            O => \N__10549\,
            I => \DRA_c_9\
        );

    \I__2523\ : Odrv12
    port map (
            O => \N__10546\,
            I => \DRA_c_9\
        );

    \I__2522\ : InMux
    port map (
            O => \N__10541\,
            I => \N__10538\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__10538\,
            I => \N__10535\
        );

    \I__2520\ : Span4Mux_h
    port map (
            O => \N__10535\,
            I => \N__10532\
        );

    \I__2519\ : Odrv4
    port map (
            O => \N__10532\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__2518\ : InMux
    port map (
            O => \N__10529\,
            I => \N__10523\
        );

    \I__2517\ : InMux
    port map (
            O => \N__10528\,
            I => \N__10520\
        );

    \I__2516\ : InMux
    port map (
            O => \N__10527\,
            I => \N__10517\
        );

    \I__2515\ : InMux
    port map (
            O => \N__10526\,
            I => \N__10514\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__10523\,
            I => \N__10511\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__10520\,
            I => \N__10508\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__10517\,
            I => \N__10503\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__10514\,
            I => \N__10503\
        );

    \I__2510\ : Span4Mux_v
    port map (
            O => \N__10511\,
            I => \N__10500\
        );

    \I__2509\ : Span4Mux_v
    port map (
            O => \N__10508\,
            I => \N__10495\
        );

    \I__2508\ : Span4Mux_v
    port map (
            O => \N__10503\,
            I => \N__10495\
        );

    \I__2507\ : Sp12to4
    port map (
            O => \N__10500\,
            I => \N__10492\
        );

    \I__2506\ : Sp12to4
    port map (
            O => \N__10495\,
            I => \N__10489\
        );

    \I__2505\ : Span12Mux_h
    port map (
            O => \N__10492\,
            I => \N__10486\
        );

    \I__2504\ : Span12Mux_h
    port map (
            O => \N__10489\,
            I => \N__10483\
        );

    \I__2503\ : Odrv12
    port map (
            O => \N__10486\,
            I => \DRA_c_7\
        );

    \I__2502\ : Odrv12
    port map (
            O => \N__10483\,
            I => \DRA_c_7\
        );

    \I__2501\ : InMux
    port map (
            O => \N__10478\,
            I => \N__10473\
        );

    \I__2500\ : InMux
    port map (
            O => \N__10477\,
            I => \N__10470\
        );

    \I__2499\ : InMux
    port map (
            O => \N__10476\,
            I => \N__10467\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__10473\,
            I => \N__10460\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__10470\,
            I => \N__10460\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__10467\,
            I => \N__10460\
        );

    \I__2495\ : Span4Mux_v
    port map (
            O => \N__10460\,
            I => \N__10456\
        );

    \I__2494\ : InMux
    port map (
            O => \N__10459\,
            I => \N__10453\
        );

    \I__2493\ : Sp12to4
    port map (
            O => \N__10456\,
            I => \N__10448\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__10453\,
            I => \N__10448\
        );

    \I__2491\ : Span12Mux_h
    port map (
            O => \N__10448\,
            I => \N__10445\
        );

    \I__2490\ : Odrv12
    port map (
            O => \N__10445\,
            I => \DRA_c_8\
        );

    \I__2489\ : InMux
    port map (
            O => \N__10442\,
            I => \N__10439\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__10439\,
            I => \N__10436\
        );

    \I__2487\ : Span4Mux_h
    port map (
            O => \N__10436\,
            I => \N__10433\
        );

    \I__2486\ : Span4Mux_h
    port map (
            O => \N__10433\,
            I => \N__10430\
        );

    \I__2485\ : Odrv4
    port map (
            O => \N__10430\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__2484\ : InMux
    port map (
            O => \N__10427\,
            I => \N__10424\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__10424\,
            I => \N__10421\
        );

    \I__2482\ : Odrv12
    port map (
            O => \N__10421\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2481\ : InMux
    port map (
            O => \N__10418\,
            I => \N__10415\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__10415\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__2479\ : InMux
    port map (
            O => \N__10412\,
            I => \N__10407\
        );

    \I__2478\ : InMux
    port map (
            O => \N__10411\,
            I => \N__10404\
        );

    \I__2477\ : InMux
    port map (
            O => \N__10410\,
            I => \N__10401\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__10407\,
            I => \N__10397\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__10404\,
            I => \N__10394\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__10401\,
            I => \N__10391\
        );

    \I__2473\ : InMux
    port map (
            O => \N__10400\,
            I => \N__10388\
        );

    \I__2472\ : Span4Mux_v
    port map (
            O => \N__10397\,
            I => \N__10385\
        );

    \I__2471\ : Span4Mux_v
    port map (
            O => \N__10394\,
            I => \N__10378\
        );

    \I__2470\ : Span4Mux_h
    port map (
            O => \N__10391\,
            I => \N__10378\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__10388\,
            I => \N__10378\
        );

    \I__2468\ : Span4Mux_v
    port map (
            O => \N__10385\,
            I => \N__10375\
        );

    \I__2467\ : Span4Mux_h
    port map (
            O => \N__10378\,
            I => \N__10372\
        );

    \I__2466\ : Sp12to4
    port map (
            O => \N__10375\,
            I => \N__10369\
        );

    \I__2465\ : Sp12to4
    port map (
            O => \N__10372\,
            I => \N__10366\
        );

    \I__2464\ : Span12Mux_h
    port map (
            O => \N__10369\,
            I => \N__10363\
        );

    \I__2463\ : Span12Mux_v
    port map (
            O => \N__10366\,
            I => \N__10360\
        );

    \I__2462\ : Odrv12
    port map (
            O => \N__10363\,
            I => \DRA_c_2\
        );

    \I__2461\ : Odrv12
    port map (
            O => \N__10360\,
            I => \DRA_c_2\
        );

    \I__2460\ : InMux
    port map (
            O => \N__10355\,
            I => \N__10349\
        );

    \I__2459\ : InMux
    port map (
            O => \N__10354\,
            I => \N__10349\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__10349\,
            I => \N__10346\
        );

    \I__2457\ : Span4Mux_h
    port map (
            O => \N__10346\,
            I => \N__10343\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__10343\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2455\ : IoInMux
    port map (
            O => \N__10340\,
            I => \N__10337\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__10337\,
            I => \N__10334\
        );

    \I__2453\ : Span4Mux_s2_h
    port map (
            O => \N__10334\,
            I => \N__10331\
        );

    \I__2452\ : Sp12to4
    port map (
            O => \N__10331\,
            I => \N__10328\
        );

    \I__2451\ : Span12Mux_s10_v
    port map (
            O => \N__10328\,
            I => \N__10325\
        );

    \I__2450\ : Odrv12
    port map (
            O => \N__10325\,
            I => \WEn_c\
        );

    \I__2449\ : InMux
    port map (
            O => \N__10322\,
            I => \N__10318\
        );

    \I__2448\ : InMux
    port map (
            O => \N__10321\,
            I => \N__10315\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__10318\,
            I => \N__10312\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__10315\,
            I => \N__10306\
        );

    \I__2445\ : Span4Mux_h
    port map (
            O => \N__10312\,
            I => \N__10306\
        );

    \I__2444\ : InMux
    port map (
            O => \N__10311\,
            I => \N__10303\
        );

    \I__2443\ : Span4Mux_v
    port map (
            O => \N__10306\,
            I => \N__10296\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__10303\,
            I => \N__10296\
        );

    \I__2441\ : InMux
    port map (
            O => \N__10302\,
            I => \N__10291\
        );

    \I__2440\ : InMux
    port map (
            O => \N__10301\,
            I => \N__10288\
        );

    \I__2439\ : Span4Mux_h
    port map (
            O => \N__10296\,
            I => \N__10285\
        );

    \I__2438\ : InMux
    port map (
            O => \N__10295\,
            I => \N__10280\
        );

    \I__2437\ : InMux
    port map (
            O => \N__10294\,
            I => \N__10280\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__10291\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__10288\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__10285\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__10280\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__10271\,
            I => \N__10268\
        );

    \I__2431\ : InMux
    port map (
            O => \N__10268\,
            I => \N__10264\
        );

    \I__2430\ : InMux
    port map (
            O => \N__10267\,
            I => \N__10261\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__10264\,
            I => \N__10255\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__10261\,
            I => \N__10255\
        );

    \I__2427\ : InMux
    port map (
            O => \N__10260\,
            I => \N__10252\
        );

    \I__2426\ : Span4Mux_v
    port map (
            O => \N__10255\,
            I => \N__10249\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__10252\,
            I => \N__10242\
        );

    \I__2424\ : Span4Mux_h
    port map (
            O => \N__10249\,
            I => \N__10242\
        );

    \I__2423\ : InMux
    port map (
            O => \N__10248\,
            I => \N__10237\
        );

    \I__2422\ : InMux
    port map (
            O => \N__10247\,
            I => \N__10237\
        );

    \I__2421\ : Odrv4
    port map (
            O => \N__10242\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__10237\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2419\ : InMux
    port map (
            O => \N__10232\,
            I => \N__10228\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10231\,
            I => \N__10225\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__10228\,
            I => \N__10221\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__10225\,
            I => \N__10218\
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__10224\,
            I => \N__10212\
        );

    \I__2414\ : Span4Mux_v
    port map (
            O => \N__10221\,
            I => \N__10206\
        );

    \I__2413\ : Span4Mux_v
    port map (
            O => \N__10218\,
            I => \N__10206\
        );

    \I__2412\ : InMux
    port map (
            O => \N__10217\,
            I => \N__10203\
        );

    \I__2411\ : CascadeMux
    port map (
            O => \N__10216\,
            I => \N__10200\
        );

    \I__2410\ : CascadeMux
    port map (
            O => \N__10215\,
            I => \N__10197\
        );

    \I__2409\ : InMux
    port map (
            O => \N__10212\,
            I => \N__10194\
        );

    \I__2408\ : InMux
    port map (
            O => \N__10211\,
            I => \N__10191\
        );

    \I__2407\ : Span4Mux_h
    port map (
            O => \N__10206\,
            I => \N__10186\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__10203\,
            I => \N__10186\
        );

    \I__2405\ : InMux
    port map (
            O => \N__10200\,
            I => \N__10181\
        );

    \I__2404\ : InMux
    port map (
            O => \N__10197\,
            I => \N__10181\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__10194\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__10191\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__10186\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__10181\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__2399\ : IoInMux
    port map (
            O => \N__10172\,
            I => \N__10169\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__10169\,
            I => \N__10166\
        );

    \I__2397\ : IoSpan4Mux
    port map (
            O => \N__10166\,
            I => \N__10163\
        );

    \I__2396\ : Span4Mux_s1_v
    port map (
            O => \N__10163\,
            I => \N__10160\
        );

    \I__2395\ : Sp12to4
    port map (
            O => \N__10160\,
            I => \N__10157\
        );

    \I__2394\ : Span12Mux_v
    port map (
            O => \N__10157\,
            I => \N__10154\
        );

    \I__2393\ : Odrv12
    port map (
            O => \N__10154\,
            I => \CMA_c_10\
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__10151\,
            I => \N__10148\
        );

    \I__2391\ : InMux
    port map (
            O => \N__10148\,
            I => \N__10145\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__10145\,
            I => \N__10142\
        );

    \I__2389\ : Span4Mux_v
    port map (
            O => \N__10142\,
            I => \N__10139\
        );

    \I__2388\ : Odrv4
    port map (
            O => \N__10139\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2387\ : InMux
    port map (
            O => \N__10136\,
            I => \N__10131\
        );

    \I__2386\ : InMux
    port map (
            O => \N__10135\,
            I => \N__10126\
        );

    \I__2385\ : InMux
    port map (
            O => \N__10134\,
            I => \N__10126\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__10131\,
            I => \N__10120\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__10126\,
            I => \N__10120\
        );

    \I__2382\ : InMux
    port map (
            O => \N__10125\,
            I => \N__10117\
        );

    \I__2381\ : Sp12to4
    port map (
            O => \N__10120\,
            I => \N__10112\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__10117\,
            I => \N__10112\
        );

    \I__2379\ : Span12Mux_v
    port map (
            O => \N__10112\,
            I => \N__10109\
        );

    \I__2378\ : Span12Mux_h
    port map (
            O => \N__10109\,
            I => \N__10106\
        );

    \I__2377\ : Odrv12
    port map (
            O => \N__10106\,
            I => \DRA_c_5\
        );

    \I__2376\ : InMux
    port map (
            O => \N__10103\,
            I => \N__10099\
        );

    \I__2375\ : InMux
    port map (
            O => \N__10102\,
            I => \N__10096\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__10099\,
            I => \N__10093\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__10096\,
            I => \N__10090\
        );

    \I__2372\ : Span4Mux_h
    port map (
            O => \N__10093\,
            I => \N__10087\
        );

    \I__2371\ : Odrv12
    port map (
            O => \N__10090\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2370\ : Odrv4
    port map (
            O => \N__10087\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2369\ : InMux
    port map (
            O => \N__10082\,
            I => \N__10079\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__10079\,
            I => \N__10076\
        );

    \I__2367\ : Span12Mux_h
    port map (
            O => \N__10076\,
            I => \N__10073\
        );

    \I__2366\ : Odrv12
    port map (
            O => \N__10073\,
            I => \RAS0n_c\
        );

    \I__2365\ : InMux
    port map (
            O => \N__10070\,
            I => \N__10067\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__10067\,
            I => \N__10064\
        );

    \I__2363\ : Span4Mux_h
    port map (
            O => \N__10064\,
            I => \N__10061\
        );

    \I__2362\ : Odrv4
    port map (
            O => \N__10061\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2361\ : CascadeMux
    port map (
            O => \N__10058\,
            I => \N__10055\
        );

    \I__2360\ : InMux
    port map (
            O => \N__10055\,
            I => \N__10045\
        );

    \I__2359\ : InMux
    port map (
            O => \N__10054\,
            I => \N__10045\
        );

    \I__2358\ : InMux
    port map (
            O => \N__10053\,
            I => \N__10040\
        );

    \I__2357\ : InMux
    port map (
            O => \N__10052\,
            I => \N__10040\
        );

    \I__2356\ : InMux
    port map (
            O => \N__10051\,
            I => \N__10037\
        );

    \I__2355\ : InMux
    port map (
            O => \N__10050\,
            I => \N__10033\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__10045\,
            I => \N__10028\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__10040\,
            I => \N__10028\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__10037\,
            I => \N__10025\
        );

    \I__2351\ : InMux
    port map (
            O => \N__10036\,
            I => \N__10021\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__10033\,
            I => \N__10018\
        );

    \I__2349\ : Span4Mux_h
    port map (
            O => \N__10028\,
            I => \N__10015\
        );

    \I__2348\ : Span4Mux_h
    port map (
            O => \N__10025\,
            I => \N__10012\
        );

    \I__2347\ : InMux
    port map (
            O => \N__10024\,
            I => \N__10009\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__10021\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2345\ : Odrv12
    port map (
            O => \N__10018\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2344\ : Odrv4
    port map (
            O => \N__10015\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2343\ : Odrv4
    port map (
            O => \N__10012\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__10009\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2341\ : CascadeMux
    port map (
            O => \N__9998\,
            I => \N__9992\
        );

    \I__2340\ : CascadeMux
    port map (
            O => \N__9997\,
            I => \N__9989\
        );

    \I__2339\ : CascadeMux
    port map (
            O => \N__9996\,
            I => \N__9984\
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__9995\,
            I => \N__9981\
        );

    \I__2337\ : InMux
    port map (
            O => \N__9992\,
            I => \N__9978\
        );

    \I__2336\ : InMux
    port map (
            O => \N__9989\,
            I => \N__9975\
        );

    \I__2335\ : InMux
    port map (
            O => \N__9988\,
            I => \N__9966\
        );

    \I__2334\ : InMux
    port map (
            O => \N__9987\,
            I => \N__9966\
        );

    \I__2333\ : InMux
    port map (
            O => \N__9984\,
            I => \N__9966\
        );

    \I__2332\ : InMux
    port map (
            O => \N__9981\,
            I => \N__9966\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__9978\,
            I => \N__9963\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__9975\,
            I => \N__9960\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__9966\,
            I => \N__9957\
        );

    \I__2328\ : Span4Mux_h
    port map (
            O => \N__9963\,
            I => \N__9954\
        );

    \I__2327\ : Odrv4
    port map (
            O => \N__9960\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__2326\ : Odrv12
    port map (
            O => \N__9957\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__9954\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__2324\ : IoInMux
    port map (
            O => \N__9947\,
            I => \N__9944\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__9944\,
            I => \N__9941\
        );

    \I__2322\ : Span4Mux_s2_v
    port map (
            O => \N__9941\,
            I => \N__9938\
        );

    \I__2321\ : Span4Mux_v
    port map (
            O => \N__9938\,
            I => \N__9935\
        );

    \I__2320\ : Span4Mux_v
    port map (
            O => \N__9935\,
            I => \N__9932\
        );

    \I__2319\ : Span4Mux_h
    port map (
            O => \N__9932\,
            I => \N__9929\
        );

    \I__2318\ : Odrv4
    port map (
            O => \N__9929\,
            I => \CMA_c_0\
        );

    \I__2317\ : InMux
    port map (
            O => \N__9926\,
            I => \N__9923\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__9923\,
            I => \N__9904\
        );

    \I__2315\ : ClkMux
    port map (
            O => \N__9922\,
            I => \N__9842\
        );

    \I__2314\ : ClkMux
    port map (
            O => \N__9921\,
            I => \N__9842\
        );

    \I__2313\ : ClkMux
    port map (
            O => \N__9920\,
            I => \N__9842\
        );

    \I__2312\ : ClkMux
    port map (
            O => \N__9919\,
            I => \N__9842\
        );

    \I__2311\ : ClkMux
    port map (
            O => \N__9918\,
            I => \N__9842\
        );

    \I__2310\ : ClkMux
    port map (
            O => \N__9917\,
            I => \N__9842\
        );

    \I__2309\ : ClkMux
    port map (
            O => \N__9916\,
            I => \N__9842\
        );

    \I__2308\ : ClkMux
    port map (
            O => \N__9915\,
            I => \N__9842\
        );

    \I__2307\ : ClkMux
    port map (
            O => \N__9914\,
            I => \N__9842\
        );

    \I__2306\ : ClkMux
    port map (
            O => \N__9913\,
            I => \N__9842\
        );

    \I__2305\ : ClkMux
    port map (
            O => \N__9912\,
            I => \N__9842\
        );

    \I__2304\ : ClkMux
    port map (
            O => \N__9911\,
            I => \N__9842\
        );

    \I__2303\ : ClkMux
    port map (
            O => \N__9910\,
            I => \N__9842\
        );

    \I__2302\ : ClkMux
    port map (
            O => \N__9909\,
            I => \N__9842\
        );

    \I__2301\ : ClkMux
    port map (
            O => \N__9908\,
            I => \N__9842\
        );

    \I__2300\ : ClkMux
    port map (
            O => \N__9907\,
            I => \N__9842\
        );

    \I__2299\ : Glb2LocalMux
    port map (
            O => \N__9904\,
            I => \N__9842\
        );

    \I__2298\ : ClkMux
    port map (
            O => \N__9903\,
            I => \N__9842\
        );

    \I__2297\ : ClkMux
    port map (
            O => \N__9902\,
            I => \N__9842\
        );

    \I__2296\ : ClkMux
    port map (
            O => \N__9901\,
            I => \N__9842\
        );

    \I__2295\ : ClkMux
    port map (
            O => \N__9900\,
            I => \N__9842\
        );

    \I__2294\ : ClkMux
    port map (
            O => \N__9899\,
            I => \N__9842\
        );

    \I__2293\ : ClkMux
    port map (
            O => \N__9898\,
            I => \N__9842\
        );

    \I__2292\ : ClkMux
    port map (
            O => \N__9897\,
            I => \N__9842\
        );

    \I__2291\ : ClkMux
    port map (
            O => \N__9896\,
            I => \N__9842\
        );

    \I__2290\ : ClkMux
    port map (
            O => \N__9895\,
            I => \N__9842\
        );

    \I__2289\ : GlobalMux
    port map (
            O => \N__9842\,
            I => \CLK80_PLL\
        );

    \I__2288\ : CEMux
    port map (
            O => \N__9839\,
            I => \N__9834\
        );

    \I__2287\ : CEMux
    port map (
            O => \N__9838\,
            I => \N__9830\
        );

    \I__2286\ : CEMux
    port map (
            O => \N__9837\,
            I => \N__9826\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__9834\,
            I => \N__9823\
        );

    \I__2284\ : CEMux
    port map (
            O => \N__9833\,
            I => \N__9820\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__9830\,
            I => \N__9817\
        );

    \I__2282\ : CEMux
    port map (
            O => \N__9829\,
            I => \N__9814\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__9826\,
            I => \N__9811\
        );

    \I__2280\ : Span4Mux_v
    port map (
            O => \N__9823\,
            I => \N__9808\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__9820\,
            I => \N__9801\
        );

    \I__2278\ : Span4Mux_h
    port map (
            O => \N__9817\,
            I => \N__9801\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__9814\,
            I => \N__9801\
        );

    \I__2276\ : Span4Mux_v
    port map (
            O => \N__9811\,
            I => \N__9798\
        );

    \I__2275\ : Span4Mux_h
    port map (
            O => \N__9808\,
            I => \N__9793\
        );

    \I__2274\ : Span4Mux_v
    port map (
            O => \N__9801\,
            I => \N__9793\
        );

    \I__2273\ : Sp12to4
    port map (
            O => \N__9798\,
            I => \N__9787\
        );

    \I__2272\ : Sp12to4
    port map (
            O => \N__9793\,
            I => \N__9787\
        );

    \I__2271\ : CEMux
    port map (
            O => \N__9792\,
            I => \N__9784\
        );

    \I__2270\ : Span12Mux_h
    port map (
            O => \N__9787\,
            I => \N__9779\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__9784\,
            I => \N__9779\
        );

    \I__2268\ : Odrv12
    port map (
            O => \N__9779\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2267\ : InMux
    port map (
            O => \N__9776\,
            I => \N__9773\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__9773\,
            I => \N__9770\
        );

    \I__2265\ : Span12Mux_h
    port map (
            O => \N__9770\,
            I => \N__9767\
        );

    \I__2264\ : Odrv12
    port map (
            O => \N__9767\,
            I => \A_c_9\
        );

    \I__2263\ : InMux
    port map (
            O => \N__9764\,
            I => \N__9761\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__9761\,
            I => \N__9758\
        );

    \I__2261\ : Span4Mux_v
    port map (
            O => \N__9758\,
            I => \N__9755\
        );

    \I__2260\ : Sp12to4
    port map (
            O => \N__9755\,
            I => \N__9752\
        );

    \I__2259\ : Span12Mux_h
    port map (
            O => \N__9752\,
            I => \N__9749\
        );

    \I__2258\ : Span12Mux_v
    port map (
            O => \N__9749\,
            I => \N__9746\
        );

    \I__2257\ : Odrv12
    port map (
            O => \N__9746\,
            I => \A_c_2\
        );

    \I__2256\ : InMux
    port map (
            O => \N__9743\,
            I => \N__9737\
        );

    \I__2255\ : InMux
    port map (
            O => \N__9742\,
            I => \N__9732\
        );

    \I__2254\ : CascadeMux
    port map (
            O => \N__9741\,
            I => \N__9728\
        );

    \I__2253\ : CascadeMux
    port map (
            O => \N__9740\,
            I => \N__9720\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__9737\,
            I => \N__9711\
        );

    \I__2251\ : InMux
    port map (
            O => \N__9736\,
            I => \N__9704\
        );

    \I__2250\ : InMux
    port map (
            O => \N__9735\,
            I => \N__9704\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__9732\,
            I => \N__9699\
        );

    \I__2248\ : InMux
    port map (
            O => \N__9731\,
            I => \N__9696\
        );

    \I__2247\ : InMux
    port map (
            O => \N__9728\,
            I => \N__9693\
        );

    \I__2246\ : InMux
    port map (
            O => \N__9727\,
            I => \N__9690\
        );

    \I__2245\ : InMux
    port map (
            O => \N__9726\,
            I => \N__9681\
        );

    \I__2244\ : InMux
    port map (
            O => \N__9725\,
            I => \N__9681\
        );

    \I__2243\ : InMux
    port map (
            O => \N__9724\,
            I => \N__9681\
        );

    \I__2242\ : InMux
    port map (
            O => \N__9723\,
            I => \N__9681\
        );

    \I__2241\ : InMux
    port map (
            O => \N__9720\,
            I => \N__9678\
        );

    \I__2240\ : InMux
    port map (
            O => \N__9719\,
            I => \N__9671\
        );

    \I__2239\ : InMux
    port map (
            O => \N__9718\,
            I => \N__9671\
        );

    \I__2238\ : InMux
    port map (
            O => \N__9717\,
            I => \N__9671\
        );

    \I__2237\ : InMux
    port map (
            O => \N__9716\,
            I => \N__9666\
        );

    \I__2236\ : InMux
    port map (
            O => \N__9715\,
            I => \N__9666\
        );

    \I__2235\ : InMux
    port map (
            O => \N__9714\,
            I => \N__9661\
        );

    \I__2234\ : Span12Mux_v
    port map (
            O => \N__9711\,
            I => \N__9658\
        );

    \I__2233\ : InMux
    port map (
            O => \N__9710\,
            I => \N__9653\
        );

    \I__2232\ : InMux
    port map (
            O => \N__9709\,
            I => \N__9653\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__9704\,
            I => \N__9650\
        );

    \I__2230\ : InMux
    port map (
            O => \N__9703\,
            I => \N__9645\
        );

    \I__2229\ : InMux
    port map (
            O => \N__9702\,
            I => \N__9645\
        );

    \I__2228\ : Span4Mux_v
    port map (
            O => \N__9699\,
            I => \N__9640\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__9696\,
            I => \N__9640\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__9693\,
            I => \N__9633\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__9690\,
            I => \N__9633\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__9681\,
            I => \N__9633\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__9678\,
            I => \N__9626\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__9671\,
            I => \N__9626\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__9666\,
            I => \N__9626\
        );

    \I__2220\ : InMux
    port map (
            O => \N__9665\,
            I => \N__9621\
        );

    \I__2219\ : InMux
    port map (
            O => \N__9664\,
            I => \N__9621\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__9661\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2217\ : Odrv12
    port map (
            O => \N__9658\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__9653\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2215\ : Odrv12
    port map (
            O => \N__9650\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__9645\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2213\ : Odrv4
    port map (
            O => \N__9640\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2212\ : Odrv4
    port map (
            O => \N__9633\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__9626\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__9621\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__9602\,
            I => \N__9599\
        );

    \I__2208\ : InMux
    port map (
            O => \N__9599\,
            I => \N__9594\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__9598\,
            I => \N__9585\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__9597\,
            I => \N__9578\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__9594\,
            I => \N__9572\
        );

    \I__2204\ : InMux
    port map (
            O => \N__9593\,
            I => \N__9569\
        );

    \I__2203\ : InMux
    port map (
            O => \N__9592\,
            I => \N__9563\
        );

    \I__2202\ : InMux
    port map (
            O => \N__9591\,
            I => \N__9560\
        );

    \I__2201\ : InMux
    port map (
            O => \N__9590\,
            I => \N__9557\
        );

    \I__2200\ : InMux
    port map (
            O => \N__9589\,
            I => \N__9554\
        );

    \I__2199\ : InMux
    port map (
            O => \N__9588\,
            I => \N__9551\
        );

    \I__2198\ : InMux
    port map (
            O => \N__9585\,
            I => \N__9548\
        );

    \I__2197\ : InMux
    port map (
            O => \N__9584\,
            I => \N__9541\
        );

    \I__2196\ : InMux
    port map (
            O => \N__9583\,
            I => \N__9541\
        );

    \I__2195\ : InMux
    port map (
            O => \N__9582\,
            I => \N__9541\
        );

    \I__2194\ : InMux
    port map (
            O => \N__9581\,
            I => \N__9536\
        );

    \I__2193\ : InMux
    port map (
            O => \N__9578\,
            I => \N__9536\
        );

    \I__2192\ : InMux
    port map (
            O => \N__9577\,
            I => \N__9529\
        );

    \I__2191\ : InMux
    port map (
            O => \N__9576\,
            I => \N__9529\
        );

    \I__2190\ : InMux
    port map (
            O => \N__9575\,
            I => \N__9529\
        );

    \I__2189\ : Span4Mux_h
    port map (
            O => \N__9572\,
            I => \N__9524\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__9569\,
            I => \N__9524\
        );

    \I__2187\ : InMux
    port map (
            O => \N__9568\,
            I => \N__9521\
        );

    \I__2186\ : InMux
    port map (
            O => \N__9567\,
            I => \N__9514\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9566\,
            I => \N__9514\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__9563\,
            I => \N__9507\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__9560\,
            I => \N__9507\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__9557\,
            I => \N__9507\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__9554\,
            I => \N__9496\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__9551\,
            I => \N__9496\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__9548\,
            I => \N__9496\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__9541\,
            I => \N__9496\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__9536\,
            I => \N__9496\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__9529\,
            I => \N__9492\
        );

    \I__2175\ : Span4Mux_v
    port map (
            O => \N__9524\,
            I => \N__9487\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__9521\,
            I => \N__9487\
        );

    \I__2173\ : InMux
    port map (
            O => \N__9520\,
            I => \N__9484\
        );

    \I__2172\ : InMux
    port map (
            O => \N__9519\,
            I => \N__9480\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__9514\,
            I => \N__9473\
        );

    \I__2170\ : Span4Mux_h
    port map (
            O => \N__9507\,
            I => \N__9473\
        );

    \I__2169\ : Span4Mux_v
    port map (
            O => \N__9496\,
            I => \N__9473\
        );

    \I__2168\ : InMux
    port map (
            O => \N__9495\,
            I => \N__9470\
        );

    \I__2167\ : Span4Mux_v
    port map (
            O => \N__9492\,
            I => \N__9463\
        );

    \I__2166\ : Span4Mux_h
    port map (
            O => \N__9487\,
            I => \N__9463\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__9484\,
            I => \N__9463\
        );

    \I__2164\ : InMux
    port map (
            O => \N__9483\,
            I => \N__9460\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__9480\,
            I => \N__9457\
        );

    \I__2162\ : Span4Mux_v
    port map (
            O => \N__9473\,
            I => \N__9454\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__9470\,
            I => \N__9449\
        );

    \I__2160\ : Span4Mux_h
    port map (
            O => \N__9463\,
            I => \N__9449\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__9460\,
            I => \CPU_CYCLE\
        );

    \I__2158\ : Odrv12
    port map (
            O => \N__9457\,
            I => \CPU_CYCLE\
        );

    \I__2157\ : Odrv4
    port map (
            O => \N__9454\,
            I => \CPU_CYCLE\
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__9449\,
            I => \CPU_CYCLE\
        );

    \I__2155\ : CascadeMux
    port map (
            O => \N__9440\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\
        );

    \I__2154\ : InMux
    port map (
            O => \N__9437\,
            I => \N__9434\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__9434\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__2152\ : InMux
    port map (
            O => \N__9431\,
            I => \N__9428\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__9428\,
            I => \N__9425\
        );

    \I__2150\ : Odrv4
    port map (
            O => \N__9425\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2149\ : InMux
    port map (
            O => \N__9422\,
            I => \N__9418\
        );

    \I__2148\ : InMux
    port map (
            O => \N__9421\,
            I => \N__9415\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__9418\,
            I => \N__9408\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__9415\,
            I => \N__9408\
        );

    \I__2145\ : InMux
    port map (
            O => \N__9414\,
            I => \N__9405\
        );

    \I__2144\ : InMux
    port map (
            O => \N__9413\,
            I => \N__9402\
        );

    \I__2143\ : Span4Mux_h
    port map (
            O => \N__9408\,
            I => \N__9395\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__9405\,
            I => \N__9395\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__9402\,
            I => \N__9395\
        );

    \I__2140\ : Span4Mux_v
    port map (
            O => \N__9395\,
            I => \N__9392\
        );

    \I__2139\ : Span4Mux_v
    port map (
            O => \N__9392\,
            I => \N__9389\
        );

    \I__2138\ : Sp12to4
    port map (
            O => \N__9389\,
            I => \N__9386\
        );

    \I__2137\ : Span12Mux_h
    port map (
            O => \N__9386\,
            I => \N__9383\
        );

    \I__2136\ : Odrv12
    port map (
            O => \N__9383\,
            I => \DRA_c_4\
        );

    \I__2135\ : InMux
    port map (
            O => \N__9380\,
            I => \N__9377\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__9377\,
            I => \N__9374\
        );

    \I__2133\ : Span4Mux_v
    port map (
            O => \N__9374\,
            I => \N__9371\
        );

    \I__2132\ : Odrv4
    port map (
            O => \N__9371\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__2131\ : InMux
    port map (
            O => \N__9368\,
            I => \N__9364\
        );

    \I__2130\ : InMux
    port map (
            O => \N__9367\,
            I => \N__9361\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__9364\,
            I => \N__9356\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__9361\,
            I => \N__9353\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9360\,
            I => \N__9350\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9359\,
            I => \N__9347\
        );

    \I__2125\ : Span4Mux_v
    port map (
            O => \N__9356\,
            I => \N__9338\
        );

    \I__2124\ : Span4Mux_h
    port map (
            O => \N__9353\,
            I => \N__9338\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__9350\,
            I => \N__9338\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__9347\,
            I => \N__9338\
        );

    \I__2121\ : Sp12to4
    port map (
            O => \N__9338\,
            I => \N__9335\
        );

    \I__2120\ : Span12Mux_v
    port map (
            O => \N__9335\,
            I => \N__9332\
        );

    \I__2119\ : Span12Mux_h
    port map (
            O => \N__9332\,
            I => \N__9329\
        );

    \I__2118\ : Odrv12
    port map (
            O => \N__9329\,
            I => \DRA_c_3\
        );

    \I__2117\ : InMux
    port map (
            O => \N__9326\,
            I => \N__9323\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__9323\,
            I => \N__9320\
        );

    \I__2115\ : Span4Mux_v
    port map (
            O => \N__9320\,
            I => \N__9317\
        );

    \I__2114\ : Odrv4
    port map (
            O => \N__9317\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__2113\ : IoInMux
    port map (
            O => \N__9314\,
            I => \N__9311\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__9311\,
            I => \N__9308\
        );

    \I__2111\ : Span4Mux_s2_v
    port map (
            O => \N__9308\,
            I => \N__9305\
        );

    \I__2110\ : Span4Mux_v
    port map (
            O => \N__9305\,
            I => \N__9302\
        );

    \I__2109\ : Odrv4
    port map (
            O => \N__9302\,
            I => \N_276_i\
        );

    \I__2108\ : IoInMux
    port map (
            O => \N__9299\,
            I => \N__9296\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__9296\,
            I => \N__9293\
        );

    \I__2106\ : Span4Mux_s2_v
    port map (
            O => \N__9293\,
            I => \N__9290\
        );

    \I__2105\ : Span4Mux_v
    port map (
            O => \N__9290\,
            I => \N__9287\
        );

    \I__2104\ : Odrv4
    port map (
            O => \N__9287\,
            I => \N_278_i\
        );

    \I__2103\ : InMux
    port map (
            O => \N__9284\,
            I => \N__9275\
        );

    \I__2102\ : InMux
    port map (
            O => \N__9283\,
            I => \N__9275\
        );

    \I__2101\ : InMux
    port map (
            O => \N__9282\,
            I => \N__9275\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__9275\,
            I => \N__9268\
        );

    \I__2099\ : InMux
    port map (
            O => \N__9274\,
            I => \N__9265\
        );

    \I__2098\ : InMux
    port map (
            O => \N__9273\,
            I => \N__9262\
        );

    \I__2097\ : InMux
    port map (
            O => \N__9272\,
            I => \N__9255\
        );

    \I__2096\ : InMux
    port map (
            O => \N__9271\,
            I => \N__9255\
        );

    \I__2095\ : Span4Mux_v
    port map (
            O => \N__9268\,
            I => \N__9250\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__9265\,
            I => \N__9250\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__9262\,
            I => \N__9247\
        );

    \I__2092\ : InMux
    port map (
            O => \N__9261\,
            I => \N__9242\
        );

    \I__2091\ : InMux
    port map (
            O => \N__9260\,
            I => \N__9239\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__9255\,
            I => \N__9236\
        );

    \I__2089\ : Span4Mux_h
    port map (
            O => \N__9250\,
            I => \N__9233\
        );

    \I__2088\ : Span4Mux_v
    port map (
            O => \N__9247\,
            I => \N__9230\
        );

    \I__2087\ : InMux
    port map (
            O => \N__9246\,
            I => \N__9227\
        );

    \I__2086\ : InMux
    port map (
            O => \N__9245\,
            I => \N__9224\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__9242\,
            I => \N__9221\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__9239\,
            I => \N__9218\
        );

    \I__2083\ : Span12Mux_v
    port map (
            O => \N__9236\,
            I => \N__9215\
        );

    \I__2082\ : Span4Mux_v
    port map (
            O => \N__9233\,
            I => \N__9210\
        );

    \I__2081\ : Span4Mux_v
    port map (
            O => \N__9230\,
            I => \N__9210\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__9227\,
            I => \N__9205\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__9224\,
            I => \N__9205\
        );

    \I__2078\ : Span4Mux_v
    port map (
            O => \N__9221\,
            I => \N__9200\
        );

    \I__2077\ : Span4Mux_v
    port map (
            O => \N__9218\,
            I => \N__9200\
        );

    \I__2076\ : Span12Mux_h
    port map (
            O => \N__9215\,
            I => \N__9197\
        );

    \I__2075\ : Sp12to4
    port map (
            O => \N__9210\,
            I => \N__9190\
        );

    \I__2074\ : Span12Mux_v
    port map (
            O => \N__9205\,
            I => \N__9190\
        );

    \I__2073\ : Sp12to4
    port map (
            O => \N__9200\,
            I => \N__9190\
        );

    \I__2072\ : Odrv12
    port map (
            O => \N__9197\,
            I => \A_c_0\
        );

    \I__2071\ : Odrv12
    port map (
            O => \N__9190\,
            I => \A_c_0\
        );

    \I__2070\ : CascadeMux
    port map (
            O => \N__9185\,
            I => \N__9181\
        );

    \I__2069\ : InMux
    port map (
            O => \N__9184\,
            I => \N__9174\
        );

    \I__2068\ : InMux
    port map (
            O => \N__9181\,
            I => \N__9171\
        );

    \I__2067\ : InMux
    port map (
            O => \N__9180\,
            I => \N__9168\
        );

    \I__2066\ : InMux
    port map (
            O => \N__9179\,
            I => \N__9160\
        );

    \I__2065\ : InMux
    port map (
            O => \N__9178\,
            I => \N__9160\
        );

    \I__2064\ : InMux
    port map (
            O => \N__9177\,
            I => \N__9160\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__9174\,
            I => \N__9157\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__9171\,
            I => \N__9152\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__9168\,
            I => \N__9152\
        );

    \I__2060\ : CascadeMux
    port map (
            O => \N__9167\,
            I => \N__9149\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__9160\,
            I => \N__9146\
        );

    \I__2058\ : Span4Mux_v
    port map (
            O => \N__9157\,
            I => \N__9143\
        );

    \I__2057\ : Span4Mux_v
    port map (
            O => \N__9152\,
            I => \N__9140\
        );

    \I__2056\ : InMux
    port map (
            O => \N__9149\,
            I => \N__9137\
        );

    \I__2055\ : Span4Mux_h
    port map (
            O => \N__9146\,
            I => \N__9134\
        );

    \I__2054\ : Sp12to4
    port map (
            O => \N__9143\,
            I => \N__9127\
        );

    \I__2053\ : Sp12to4
    port map (
            O => \N__9140\,
            I => \N__9127\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__9137\,
            I => \N__9127\
        );

    \I__2051\ : Span4Mux_v
    port map (
            O => \N__9134\,
            I => \N__9124\
        );

    \I__2050\ : Span12Mux_h
    port map (
            O => \N__9127\,
            I => \N__9121\
        );

    \I__2049\ : Sp12to4
    port map (
            O => \N__9124\,
            I => \N__9118\
        );

    \I__2048\ : Span12Mux_v
    port map (
            O => \N__9121\,
            I => \N__9113\
        );

    \I__2047\ : Span12Mux_h
    port map (
            O => \N__9118\,
            I => \N__9113\
        );

    \I__2046\ : Odrv12
    port map (
            O => \N__9113\,
            I => \SIZ_c_0\
        );

    \I__2045\ : InMux
    port map (
            O => \N__9110\,
            I => \N__9105\
        );

    \I__2044\ : CascadeMux
    port map (
            O => \N__9109\,
            I => \N__9101\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__9108\,
            I => \N__9098\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__9105\,
            I => \N__9095\
        );

    \I__2041\ : InMux
    port map (
            O => \N__9104\,
            I => \N__9085\
        );

    \I__2040\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9085\
        );

    \I__2039\ : InMux
    port map (
            O => \N__9098\,
            I => \N__9085\
        );

    \I__2038\ : Span4Mux_v
    port map (
            O => \N__9095\,
            I => \N__9081\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__9094\,
            I => \N__9078\
        );

    \I__2036\ : InMux
    port map (
            O => \N__9093\,
            I => \N__9073\
        );

    \I__2035\ : InMux
    port map (
            O => \N__9092\,
            I => \N__9073\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__9085\,
            I => \N__9070\
        );

    \I__2033\ : InMux
    port map (
            O => \N__9084\,
            I => \N__9067\
        );

    \I__2032\ : Span4Mux_v
    port map (
            O => \N__9081\,
            I => \N__9064\
        );

    \I__2031\ : InMux
    port map (
            O => \N__9078\,
            I => \N__9061\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__9073\,
            I => \N__9058\
        );

    \I__2029\ : Span4Mux_v
    port map (
            O => \N__9070\,
            I => \N__9055\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__9067\,
            I => \N__9052\
        );

    \I__2027\ : Span4Mux_v
    port map (
            O => \N__9064\,
            I => \N__9049\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__9061\,
            I => \N__9046\
        );

    \I__2025\ : Span12Mux_v
    port map (
            O => \N__9058\,
            I => \N__9039\
        );

    \I__2024\ : Sp12to4
    port map (
            O => \N__9055\,
            I => \N__9039\
        );

    \I__2023\ : Span12Mux_s7_v
    port map (
            O => \N__9052\,
            I => \N__9039\
        );

    \I__2022\ : Sp12to4
    port map (
            O => \N__9049\,
            I => \N__9034\
        );

    \I__2021\ : Span12Mux_v
    port map (
            O => \N__9046\,
            I => \N__9034\
        );

    \I__2020\ : Span12Mux_h
    port map (
            O => \N__9039\,
            I => \N__9031\
        );

    \I__2019\ : Odrv12
    port map (
            O => \N__9034\,
            I => \A_c_1\
        );

    \I__2018\ : Odrv12
    port map (
            O => \N__9031\,
            I => \A_c_1\
        );

    \I__2017\ : CascadeMux
    port map (
            O => \N__9026\,
            I => \N__9023\
        );

    \I__2016\ : InMux
    port map (
            O => \N__9023\,
            I => \N__9017\
        );

    \I__2015\ : InMux
    port map (
            O => \N__9022\,
            I => \N__9014\
        );

    \I__2014\ : InMux
    port map (
            O => \N__9021\,
            I => \N__9011\
        );

    \I__2013\ : CascadeMux
    port map (
            O => \N__9020\,
            I => \N__9008\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__9017\,
            I => \N__9003\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__9014\,
            I => \N__8998\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__9011\,
            I => \N__8998\
        );

    \I__2009\ : InMux
    port map (
            O => \N__9008\,
            I => \N__8990\
        );

    \I__2008\ : InMux
    port map (
            O => \N__9007\,
            I => \N__8990\
        );

    \I__2007\ : InMux
    port map (
            O => \N__9006\,
            I => \N__8990\
        );

    \I__2006\ : Span4Mux_v
    port map (
            O => \N__9003\,
            I => \N__8987\
        );

    \I__2005\ : Span4Mux_v
    port map (
            O => \N__8998\,
            I => \N__8984\
        );

    \I__2004\ : InMux
    port map (
            O => \N__8997\,
            I => \N__8981\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__8990\,
            I => \N__8978\
        );

    \I__2002\ : Sp12to4
    port map (
            O => \N__8987\,
            I => \N__8971\
        );

    \I__2001\ : Sp12to4
    port map (
            O => \N__8984\,
            I => \N__8971\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__8981\,
            I => \N__8971\
        );

    \I__1999\ : Sp12to4
    port map (
            O => \N__8978\,
            I => \N__8968\
        );

    \I__1998\ : Span12Mux_h
    port map (
            O => \N__8971\,
            I => \N__8965\
        );

    \I__1997\ : Span12Mux_v
    port map (
            O => \N__8968\,
            I => \N__8962\
        );

    \I__1996\ : Span12Mux_v
    port map (
            O => \N__8965\,
            I => \N__8957\
        );

    \I__1995\ : Span12Mux_h
    port map (
            O => \N__8962\,
            I => \N__8957\
        );

    \I__1994\ : Odrv12
    port map (
            O => \N__8957\,
            I => \SIZ_c_1\
        );

    \I__1993\ : IoInMux
    port map (
            O => \N__8954\,
            I => \N__8951\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__8951\,
            I => \N__8948\
        );

    \I__1991\ : Span4Mux_s2_v
    port map (
            O => \N__8948\,
            I => \N__8945\
        );

    \I__1990\ : Span4Mux_h
    port map (
            O => \N__8945\,
            I => \N__8942\
        );

    \I__1989\ : Span4Mux_v
    port map (
            O => \N__8942\,
            I => \N__8939\
        );

    \I__1988\ : Odrv4
    port map (
            O => \N__8939\,
            I => \N_277_i\
        );

    \I__1987\ : IoInMux
    port map (
            O => \N__8936\,
            I => \N__8933\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__8933\,
            I => \N__8930\
        );

    \I__1985\ : IoSpan4Mux
    port map (
            O => \N__8930\,
            I => \N__8927\
        );

    \I__1984\ : Sp12to4
    port map (
            O => \N__8927\,
            I => \N__8924\
        );

    \I__1983\ : Span12Mux_s9_v
    port map (
            O => \N__8924\,
            I => \N__8921\
        );

    \I__1982\ : Odrv12
    port map (
            O => \N__8921\,
            I => \CRCSn_c\
        );

    \I__1981\ : IoInMux
    port map (
            O => \N__8918\,
            I => \N__8915\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__8915\,
            I => \N__8912\
        );

    \I__1979\ : Span4Mux_s1_v
    port map (
            O => \N__8912\,
            I => \N__8909\
        );

    \I__1978\ : Span4Mux_v
    port map (
            O => \N__8909\,
            I => \N__8906\
        );

    \I__1977\ : Span4Mux_v
    port map (
            O => \N__8906\,
            I => \N__8903\
        );

    \I__1976\ : Sp12to4
    port map (
            O => \N__8903\,
            I => \N__8900\
        );

    \I__1975\ : Odrv12
    port map (
            O => \N__8900\,
            I => \RASn_c\
        );

    \I__1974\ : IoInMux
    port map (
            O => \N__8897\,
            I => \N__8894\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__8894\,
            I => \N__8891\
        );

    \I__1972\ : Span4Mux_s1_v
    port map (
            O => \N__8891\,
            I => \N__8888\
        );

    \I__1971\ : Sp12to4
    port map (
            O => \N__8888\,
            I => \N__8885\
        );

    \I__1970\ : Span12Mux_h
    port map (
            O => \N__8885\,
            I => \N__8882\
        );

    \I__1969\ : Odrv12
    port map (
            O => \N__8882\,
            I => \CASn_c\
        );

    \I__1968\ : InMux
    port map (
            O => \N__8879\,
            I => \N__8875\
        );

    \I__1967\ : InMux
    port map (
            O => \N__8878\,
            I => \N__8872\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__8875\,
            I => \N__8866\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__8872\,
            I => \N__8858\
        );

    \I__1964\ : ClkMux
    port map (
            O => \N__8871\,
            I => \N__8837\
        );

    \I__1963\ : ClkMux
    port map (
            O => \N__8870\,
            I => \N__8837\
        );

    \I__1962\ : ClkMux
    port map (
            O => \N__8869\,
            I => \N__8837\
        );

    \I__1961\ : Glb2LocalMux
    port map (
            O => \N__8866\,
            I => \N__8837\
        );

    \I__1960\ : ClkMux
    port map (
            O => \N__8865\,
            I => \N__8837\
        );

    \I__1959\ : ClkMux
    port map (
            O => \N__8864\,
            I => \N__8837\
        );

    \I__1958\ : ClkMux
    port map (
            O => \N__8863\,
            I => \N__8837\
        );

    \I__1957\ : ClkMux
    port map (
            O => \N__8862\,
            I => \N__8837\
        );

    \I__1956\ : ClkMux
    port map (
            O => \N__8861\,
            I => \N__8837\
        );

    \I__1955\ : Glb2LocalMux
    port map (
            O => \N__8858\,
            I => \N__8837\
        );

    \I__1954\ : GlobalMux
    port map (
            O => \N__8837\,
            I => \N__8834\
        );

    \I__1953\ : gio2CtrlBuf
    port map (
            O => \N__8834\,
            I => \CLK40_PLL_g\
        );

    \I__1952\ : IoInMux
    port map (
            O => \N__8831\,
            I => \N__8828\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__8828\,
            I => \N__8824\
        );

    \I__1950\ : IoInMux
    port map (
            O => \N__8827\,
            I => \N__8821\
        );

    \I__1949\ : IoSpan4Mux
    port map (
            O => \N__8824\,
            I => \N__8817\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__8821\,
            I => \N__8814\
        );

    \I__1947\ : IoInMux
    port map (
            O => \N__8820\,
            I => \N__8811\
        );

    \I__1946\ : IoSpan4Mux
    port map (
            O => \N__8817\,
            I => \N__8808\
        );

    \I__1945\ : Span4Mux_s3_v
    port map (
            O => \N__8814\,
            I => \N__8805\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__8811\,
            I => \N__8802\
        );

    \I__1943\ : Span4Mux_s3_v
    port map (
            O => \N__8808\,
            I => \N__8797\
        );

    \I__1942\ : Span4Mux_h
    port map (
            O => \N__8805\,
            I => \N__8797\
        );

    \I__1941\ : Span12Mux_s3_h
    port map (
            O => \N__8802\,
            I => \N__8794\
        );

    \I__1940\ : Span4Mux_h
    port map (
            O => \N__8797\,
            I => \N__8791\
        );

    \I__1939\ : Span12Mux_h
    port map (
            O => \N__8794\,
            I => \N__8788\
        );

    \I__1938\ : Span4Mux_h
    port map (
            O => \N__8791\,
            I => \N__8785\
        );

    \I__1937\ : Odrv12
    port map (
            O => \N__8788\,
            I => \CLK40_PLL_iso_i\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__8785\,
            I => \CLK40_PLL_iso_i\
        );

    \I__1935\ : IoInMux
    port map (
            O => \N__8780\,
            I => \N__8777\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__8777\,
            I => \N__8774\
        );

    \I__1933\ : IoSpan4Mux
    port map (
            O => \N__8774\,
            I => \N__8771\
        );

    \I__1932\ : Span4Mux_s3_v
    port map (
            O => \N__8771\,
            I => \N__8768\
        );

    \I__1931\ : Odrv4
    port map (
            O => \N__8768\,
            I => \U712_BYTE_ENABLE_UUBE_i\
        );

    \I__1930\ : InMux
    port map (
            O => \N__8765\,
            I => \N__8761\
        );

    \I__1929\ : CascadeMux
    port map (
            O => \N__8764\,
            I => \N__8758\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__8761\,
            I => \N__8755\
        );

    \I__1927\ : InMux
    port map (
            O => \N__8758\,
            I => \N__8751\
        );

    \I__1926\ : Span4Mux_h
    port map (
            O => \N__8755\,
            I => \N__8748\
        );

    \I__1925\ : InMux
    port map (
            O => \N__8754\,
            I => \N__8745\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__8751\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1923\ : Odrv4
    port map (
            O => \N__8748\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__8745\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1921\ : InMux
    port map (
            O => \N__8738\,
            I => \N__8735\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__8735\,
            I => \N__8732\
        );

    \I__1919\ : Span4Mux_v
    port map (
            O => \N__8732\,
            I => \N__8729\
        );

    \I__1918\ : Span4Mux_v
    port map (
            O => \N__8729\,
            I => \N__8726\
        );

    \I__1917\ : Sp12to4
    port map (
            O => \N__8726\,
            I => \N__8723\
        );

    \I__1916\ : Span12Mux_h
    port map (
            O => \N__8723\,
            I => \N__8720\
        );

    \I__1915\ : Odrv12
    port map (
            O => \N__8720\,
            I => \A_c_17\
        );

    \I__1914\ : IoInMux
    port map (
            O => \N__8717\,
            I => \N__8714\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__8714\,
            I => \N__8711\
        );

    \I__1912\ : Span12Mux_s3_h
    port map (
            O => \N__8711\,
            I => \N__8708\
        );

    \I__1911\ : Span12Mux_h
    port map (
            O => \N__8708\,
            I => \N__8705\
        );

    \I__1910\ : Odrv12
    port map (
            O => \N__8705\,
            I => \CMA_c_8\
        );

    \I__1909\ : InMux
    port map (
            O => \N__8702\,
            I => \N__8699\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8699\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__1907\ : InMux
    port map (
            O => \N__8696\,
            I => \N__8693\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__8693\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__1905\ : InMux
    port map (
            O => \N__8690\,
            I => \N__8687\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__8687\,
            I => \N__8684\
        );

    \I__1903\ : Span4Mux_v
    port map (
            O => \N__8684\,
            I => \N__8681\
        );

    \I__1902\ : Odrv4
    port map (
            O => \N__8681\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__1901\ : InMux
    port map (
            O => \N__8678\,
            I => \N__8675\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__8675\,
            I => \N__8672\
        );

    \I__1899\ : Span4Mux_v
    port map (
            O => \N__8672\,
            I => \N__8669\
        );

    \I__1898\ : Odrv4
    port map (
            O => \N__8669\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__1897\ : InMux
    port map (
            O => \N__8666\,
            I => \N__8663\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__8663\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__1895\ : InMux
    port map (
            O => \N__8660\,
            I => \N__8657\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__8657\,
            I => \N__8654\
        );

    \I__1893\ : Span4Mux_h
    port map (
            O => \N__8654\,
            I => \N__8651\
        );

    \I__1892\ : Odrv4
    port map (
            O => \N__8651\,
            I => \U712_CHIP_RAM.N_456\
        );

    \I__1891\ : InMux
    port map (
            O => \N__8648\,
            I => \N__8645\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__8645\,
            I => \N__8642\
        );

    \I__1889\ : Odrv4
    port map (
            O => \N__8642\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__1888\ : CascadeMux
    port map (
            O => \N__8639\,
            I => \N__8636\
        );

    \I__1887\ : InMux
    port map (
            O => \N__8636\,
            I => \N__8631\
        );

    \I__1886\ : CascadeMux
    port map (
            O => \N__8635\,
            I => \N__8625\
        );

    \I__1885\ : CascadeMux
    port map (
            O => \N__8634\,
            I => \N__8620\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__8631\,
            I => \N__8617\
        );

    \I__1883\ : InMux
    port map (
            O => \N__8630\,
            I => \N__8608\
        );

    \I__1882\ : InMux
    port map (
            O => \N__8629\,
            I => \N__8608\
        );

    \I__1881\ : InMux
    port map (
            O => \N__8628\,
            I => \N__8608\
        );

    \I__1880\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8608\
        );

    \I__1879\ : InMux
    port map (
            O => \N__8624\,
            I => \N__8601\
        );

    \I__1878\ : InMux
    port map (
            O => \N__8623\,
            I => \N__8601\
        );

    \I__1877\ : InMux
    port map (
            O => \N__8620\,
            I => \N__8601\
        );

    \I__1876\ : Odrv4
    port map (
            O => \N__8617\,
            I => \U712_CHIP_RAM.N_202\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__8608\,
            I => \U712_CHIP_RAM.N_202\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__8601\,
            I => \U712_CHIP_RAM.N_202\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8594\,
            I => \N__8591\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__8591\,
            I => \N__8588\
        );

    \I__1871\ : Span4Mux_h
    port map (
            O => \N__8588\,
            I => \N__8585\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__8585\,
            I => \U712_CHIP_RAM.N_359\
        );

    \I__1869\ : InMux
    port map (
            O => \N__8582\,
            I => \N__8575\
        );

    \I__1868\ : InMux
    port map (
            O => \N__8581\,
            I => \N__8572\
        );

    \I__1867\ : InMux
    port map (
            O => \N__8580\,
            I => \N__8569\
        );

    \I__1866\ : InMux
    port map (
            O => \N__8579\,
            I => \N__8566\
        );

    \I__1865\ : InMux
    port map (
            O => \N__8578\,
            I => \N__8563\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__8575\,
            I => \N__8548\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__8572\,
            I => \N__8548\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__8569\,
            I => \N__8548\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__8566\,
            I => \N__8548\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__8563\,
            I => \N__8545\
        );

    \I__1859\ : InMux
    port map (
            O => \N__8562\,
            I => \N__8542\
        );

    \I__1858\ : InMux
    port map (
            O => \N__8561\,
            I => \N__8539\
        );

    \I__1857\ : InMux
    port map (
            O => \N__8560\,
            I => \N__8534\
        );

    \I__1856\ : InMux
    port map (
            O => \N__8559\,
            I => \N__8534\
        );

    \I__1855\ : InMux
    port map (
            O => \N__8558\,
            I => \N__8529\
        );

    \I__1854\ : InMux
    port map (
            O => \N__8557\,
            I => \N__8529\
        );

    \I__1853\ : Span4Mux_h
    port map (
            O => \N__8548\,
            I => \N__8526\
        );

    \I__1852\ : Odrv4
    port map (
            O => \N__8545\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__8542\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__8539\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__8534\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__8529\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1847\ : Odrv4
    port map (
            O => \N__8526\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1846\ : CEMux
    port map (
            O => \N__8513\,
            I => \N__8510\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__8510\,
            I => \N__8506\
        );

    \I__1844\ : CEMux
    port map (
            O => \N__8509\,
            I => \N__8503\
        );

    \I__1843\ : Odrv4
    port map (
            O => \N__8506\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__8503\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__1841\ : InMux
    port map (
            O => \N__8498\,
            I => \N__8494\
        );

    \I__1840\ : InMux
    port map (
            O => \N__8497\,
            I => \N__8489\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__8494\,
            I => \N__8485\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8493\,
            I => \N__8480\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8492\,
            I => \N__8480\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__8489\,
            I => \N__8476\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8488\,
            I => \N__8473\
        );

    \I__1834\ : Span4Mux_v
    port map (
            O => \N__8485\,
            I => \N__8470\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__8480\,
            I => \N__8467\
        );

    \I__1832\ : InMux
    port map (
            O => \N__8479\,
            I => \N__8464\
        );

    \I__1831\ : Span4Mux_v
    port map (
            O => \N__8476\,
            I => \N__8450\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8473\,
            I => \N__8450\
        );

    \I__1829\ : Span4Mux_h
    port map (
            O => \N__8470\,
            I => \N__8443\
        );

    \I__1828\ : Span4Mux_v
    port map (
            O => \N__8467\,
            I => \N__8443\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8464\,
            I => \N__8443\
        );

    \I__1826\ : InMux
    port map (
            O => \N__8463\,
            I => \N__8438\
        );

    \I__1825\ : InMux
    port map (
            O => \N__8462\,
            I => \N__8438\
        );

    \I__1824\ : InMux
    port map (
            O => \N__8461\,
            I => \N__8433\
        );

    \I__1823\ : InMux
    port map (
            O => \N__8460\,
            I => \N__8433\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8459\,
            I => \N__8429\
        );

    \I__1821\ : InMux
    port map (
            O => \N__8458\,
            I => \N__8420\
        );

    \I__1820\ : InMux
    port map (
            O => \N__8457\,
            I => \N__8420\
        );

    \I__1819\ : InMux
    port map (
            O => \N__8456\,
            I => \N__8420\
        );

    \I__1818\ : InMux
    port map (
            O => \N__8455\,
            I => \N__8420\
        );

    \I__1817\ : Span4Mux_v
    port map (
            O => \N__8450\,
            I => \N__8417\
        );

    \I__1816\ : Sp12to4
    port map (
            O => \N__8443\,
            I => \N__8412\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__8438\,
            I => \N__8412\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__8433\,
            I => \N__8409\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8432\,
            I => \N__8406\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__8429\,
            I => \N__8401\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__8420\,
            I => \N__8401\
        );

    \I__1810\ : Sp12to4
    port map (
            O => \N__8417\,
            I => \N__8392\
        );

    \I__1809\ : Span12Mux_v
    port map (
            O => \N__8412\,
            I => \N__8392\
        );

    \I__1808\ : Span12Mux_v
    port map (
            O => \N__8409\,
            I => \N__8392\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__8406\,
            I => \N__8392\
        );

    \I__1806\ : Span12Mux_h
    port map (
            O => \N__8401\,
            I => \N__8389\
        );

    \I__1805\ : Span12Mux_h
    port map (
            O => \N__8392\,
            I => \N__8386\
        );

    \I__1804\ : Odrv12
    port map (
            O => \N__8389\,
            I => \RESETn_c\
        );

    \I__1803\ : Odrv12
    port map (
            O => \N__8386\,
            I => \RESETn_c\
        );

    \I__1802\ : IoInMux
    port map (
            O => \N__8381\,
            I => \N__8378\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__8378\,
            I => \N__8375\
        );

    \I__1800\ : Span12Mux_s8_v
    port map (
            O => \N__8375\,
            I => \N__8371\
        );

    \I__1799\ : InMux
    port map (
            O => \N__8374\,
            I => \N__8368\
        );

    \I__1798\ : Odrv12
    port map (
            O => \N__8371\,
            I => \RESETn_c_i\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__8368\,
            I => \RESETn_c_i\
        );

    \I__1796\ : CascadeMux
    port map (
            O => \N__8363\,
            I => \N__8359\
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__8362\,
            I => \N__8355\
        );

    \I__1794\ : InMux
    port map (
            O => \N__8359\,
            I => \N__8350\
        );

    \I__1793\ : InMux
    port map (
            O => \N__8358\,
            I => \N__8350\
        );

    \I__1792\ : InMux
    port map (
            O => \N__8355\,
            I => \N__8347\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__8350\,
            I => \N__8344\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__8347\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1789\ : Odrv12
    port map (
            O => \N__8344\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1788\ : CascadeMux
    port map (
            O => \N__8339\,
            I => \N__8336\
        );

    \I__1787\ : InMux
    port map (
            O => \N__8336\,
            I => \N__8332\
        );

    \I__1786\ : IoInMux
    port map (
            O => \N__8335\,
            I => \N__8329\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__8332\,
            I => \N__8325\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__8329\,
            I => \N__8322\
        );

    \I__1783\ : InMux
    port map (
            O => \N__8328\,
            I => \N__8319\
        );

    \I__1782\ : Span4Mux_h
    port map (
            O => \N__8325\,
            I => \N__8316\
        );

    \I__1781\ : Span12Mux_s3_h
    port map (
            O => \N__8322\,
            I => \N__8313\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__8319\,
            I => \N__8310\
        );

    \I__1779\ : Span4Mux_h
    port map (
            O => \N__8316\,
            I => \N__8307\
        );

    \I__1778\ : Span12Mux_v
    port map (
            O => \N__8313\,
            I => \N__8304\
        );

    \I__1777\ : Sp12to4
    port map (
            O => \N__8310\,
            I => \N__8299\
        );

    \I__1776\ : Sp12to4
    port map (
            O => \N__8307\,
            I => \N__8299\
        );

    \I__1775\ : Span12Mux_h
    port map (
            O => \N__8304\,
            I => \N__8296\
        );

    \I__1774\ : Span12Mux_v
    port map (
            O => \N__8299\,
            I => \N__8293\
        );

    \I__1773\ : Odrv12
    port map (
            O => \N__8296\,
            I => \CLK40_PLL\
        );

    \I__1772\ : Odrv12
    port map (
            O => \N__8293\,
            I => \CLK40_PLL\
        );

    \I__1771\ : InMux
    port map (
            O => \N__8288\,
            I => \N__8285\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__8285\,
            I => \N__8281\
        );

    \I__1769\ : InMux
    port map (
            O => \N__8284\,
            I => \N__8278\
        );

    \I__1768\ : Span4Mux_v
    port map (
            O => \N__8281\,
            I => \N__8275\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__8278\,
            I => \N__8272\
        );

    \I__1766\ : Sp12to4
    port map (
            O => \N__8275\,
            I => \N__8267\
        );

    \I__1765\ : Span12Mux_v
    port map (
            O => \N__8272\,
            I => \N__8267\
        );

    \I__1764\ : Odrv12
    port map (
            O => \N__8267\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__1763\ : InMux
    port map (
            O => \N__8264\,
            I => \N__8261\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__8261\,
            I => \U712_CYCLE_TERM.N_8\
        );

    \I__1761\ : CascadeMux
    port map (
            O => \N__8258\,
            I => \N__8253\
        );

    \I__1760\ : InMux
    port map (
            O => \N__8257\,
            I => \N__8250\
        );

    \I__1759\ : InMux
    port map (
            O => \N__8256\,
            I => \N__8245\
        );

    \I__1758\ : InMux
    port map (
            O => \N__8253\,
            I => \N__8242\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__8250\,
            I => \N__8239\
        );

    \I__1756\ : InMux
    port map (
            O => \N__8249\,
            I => \N__8236\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8248\,
            I => \N__8233\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__8245\,
            I => \N__8228\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__8242\,
            I => \N__8228\
        );

    \I__1752\ : Span4Mux_h
    port map (
            O => \N__8239\,
            I => \N__8225\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__8236\,
            I => \REG_TACK\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__8233\,
            I => \REG_TACK\
        );

    \I__1749\ : Odrv12
    port map (
            O => \N__8228\,
            I => \REG_TACK\
        );

    \I__1748\ : Odrv4
    port map (
            O => \N__8225\,
            I => \REG_TACK\
        );

    \I__1747\ : InMux
    port map (
            O => \N__8216\,
            I => \N__8213\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__8213\,
            I => \N__8208\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__8212\,
            I => \N__8205\
        );

    \I__1744\ : InMux
    port map (
            O => \N__8211\,
            I => \N__8201\
        );

    \I__1743\ : Span4Mux_h
    port map (
            O => \N__8208\,
            I => \N__8198\
        );

    \I__1742\ : InMux
    port map (
            O => \N__8205\,
            I => \N__8195\
        );

    \I__1741\ : InMux
    port map (
            O => \N__8204\,
            I => \N__8191\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__8201\,
            I => \N__8186\
        );

    \I__1739\ : Span4Mux_h
    port map (
            O => \N__8198\,
            I => \N__8186\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__8195\,
            I => \N__8183\
        );

    \I__1737\ : InMux
    port map (
            O => \N__8194\,
            I => \N__8180\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__8191\,
            I => \CPU_TACK\
        );

    \I__1735\ : Odrv4
    port map (
            O => \N__8186\,
            I => \CPU_TACK\
        );

    \I__1734\ : Odrv12
    port map (
            O => \N__8183\,
            I => \CPU_TACK\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__8180\,
            I => \CPU_TACK\
        );

    \I__1732\ : InMux
    port map (
            O => \N__8171\,
            I => \N__8164\
        );

    \I__1731\ : InMux
    port map (
            O => \N__8170\,
            I => \N__8164\
        );

    \I__1730\ : InMux
    port map (
            O => \N__8169\,
            I => \N__8161\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__8164\,
            I => \N__8158\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__8161\,
            I => \N__8155\
        );

    \I__1727\ : Span4Mux_v
    port map (
            O => \N__8158\,
            I => \N__8148\
        );

    \I__1726\ : Span4Mux_h
    port map (
            O => \N__8155\,
            I => \N__8148\
        );

    \I__1725\ : InMux
    port map (
            O => \N__8154\,
            I => \N__8142\
        );

    \I__1724\ : InMux
    port map (
            O => \N__8153\,
            I => \N__8142\
        );

    \I__1723\ : Span4Mux_h
    port map (
            O => \N__8148\,
            I => \N__8139\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8147\,
            I => \N__8136\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__8142\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1720\ : Odrv4
    port map (
            O => \N__8139\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__8136\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8129\,
            I => \N__8126\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__8126\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1716\ : InMux
    port map (
            O => \N__8123\,
            I => \N__8119\
        );

    \I__1715\ : InMux
    port map (
            O => \N__8122\,
            I => \N__8116\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__8119\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__8116\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1712\ : InMux
    port map (
            O => \N__8111\,
            I => \N__8108\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__8108\,
            I => \N__8104\
        );

    \I__1710\ : InMux
    port map (
            O => \N__8107\,
            I => \N__8101\
        );

    \I__1709\ : Span4Mux_v
    port map (
            O => \N__8104\,
            I => \N__8098\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__8101\,
            I => \N__8095\
        );

    \I__1707\ : Span4Mux_h
    port map (
            O => \N__8098\,
            I => \N__8090\
        );

    \I__1706\ : Span4Mux_v
    port map (
            O => \N__8095\,
            I => \N__8087\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8094\,
            I => \N__8084\
        );

    \I__1704\ : InMux
    port map (
            O => \N__8093\,
            I => \N__8081\
        );

    \I__1703\ : Sp12to4
    port map (
            O => \N__8090\,
            I => \N__8078\
        );

    \I__1702\ : Sp12to4
    port map (
            O => \N__8087\,
            I => \N__8071\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__8084\,
            I => \N__8071\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8081\,
            I => \N__8071\
        );

    \I__1699\ : Span12Mux_h
    port map (
            O => \N__8078\,
            I => \N__8068\
        );

    \I__1698\ : Span12Mux_v
    port map (
            O => \N__8071\,
            I => \N__8065\
        );

    \I__1697\ : Span12Mux_v
    port map (
            O => \N__8068\,
            I => \N__8060\
        );

    \I__1696\ : Span12Mux_h
    port map (
            O => \N__8065\,
            I => \N__8060\
        );

    \I__1695\ : Odrv12
    port map (
            O => \N__8060\,
            I => \CASLn_c\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8057\,
            I => \N__8053\
        );

    \I__1693\ : InMux
    port map (
            O => \N__8056\,
            I => \N__8050\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__8053\,
            I => \N__8046\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__8050\,
            I => \N__8043\
        );

    \I__1690\ : InMux
    port map (
            O => \N__8049\,
            I => \N__8040\
        );

    \I__1689\ : Span4Mux_v
    port map (
            O => \N__8046\,
            I => \N__8034\
        );

    \I__1688\ : Span4Mux_v
    port map (
            O => \N__8043\,
            I => \N__8034\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__8040\,
            I => \N__8031\
        );

    \I__1686\ : InMux
    port map (
            O => \N__8039\,
            I => \N__8028\
        );

    \I__1685\ : Span4Mux_v
    port map (
            O => \N__8034\,
            I => \N__8021\
        );

    \I__1684\ : Span4Mux_h
    port map (
            O => \N__8031\,
            I => \N__8021\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__8028\,
            I => \N__8021\
        );

    \I__1682\ : Span4Mux_v
    port map (
            O => \N__8021\,
            I => \N__8018\
        );

    \I__1681\ : Span4Mux_v
    port map (
            O => \N__8018\,
            I => \N__8015\
        );

    \I__1680\ : Sp12to4
    port map (
            O => \N__8015\,
            I => \N__8012\
        );

    \I__1679\ : Span12Mux_h
    port map (
            O => \N__8012\,
            I => \N__8009\
        );

    \I__1678\ : Odrv12
    port map (
            O => \N__8009\,
            I => \CASUn_c\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8006\,
            I => \N__8002\
        );

    \I__1676\ : InMux
    port map (
            O => \N__8005\,
            I => \N__7999\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__8002\,
            I => \N__7996\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__7999\,
            I => \N__7993\
        );

    \I__1673\ : Span4Mux_v
    port map (
            O => \N__7996\,
            I => \N__7989\
        );

    \I__1672\ : Span4Mux_v
    port map (
            O => \N__7993\,
            I => \N__7986\
        );

    \I__1671\ : InMux
    port map (
            O => \N__7992\,
            I => \N__7983\
        );

    \I__1670\ : Odrv4
    port map (
            O => \N__7989\,
            I => \REG_CYCLE\
        );

    \I__1669\ : Odrv4
    port map (
            O => \N__7986\,
            I => \REG_CYCLE\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__7983\,
            I => \REG_CYCLE\
        );

    \I__1667\ : IoInMux
    port map (
            O => \N__7976\,
            I => \N__7973\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__7973\,
            I => \N__7970\
        );

    \I__1665\ : IoSpan4Mux
    port map (
            O => \N__7970\,
            I => \N__7967\
        );

    \I__1664\ : Span4Mux_s1_v
    port map (
            O => \N__7967\,
            I => \N__7964\
        );

    \I__1663\ : Sp12to4
    port map (
            O => \N__7964\,
            I => \N__7961\
        );

    \I__1662\ : Span12Mux_h
    port map (
            O => \N__7961\,
            I => \N__7958\
        );

    \I__1661\ : Odrv12
    port map (
            O => \N__7958\,
            I => \DRDENn_c\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__7955\,
            I => \N__7949\
        );

    \I__1659\ : CascadeMux
    port map (
            O => \N__7954\,
            I => \N__7943\
        );

    \I__1658\ : InMux
    port map (
            O => \N__7953\,
            I => \N__7935\
        );

    \I__1657\ : InMux
    port map (
            O => \N__7952\,
            I => \N__7932\
        );

    \I__1656\ : InMux
    port map (
            O => \N__7949\,
            I => \N__7927\
        );

    \I__1655\ : InMux
    port map (
            O => \N__7948\,
            I => \N__7927\
        );

    \I__1654\ : InMux
    port map (
            O => \N__7947\,
            I => \N__7924\
        );

    \I__1653\ : InMux
    port map (
            O => \N__7946\,
            I => \N__7919\
        );

    \I__1652\ : InMux
    port map (
            O => \N__7943\,
            I => \N__7919\
        );

    \I__1651\ : InMux
    port map (
            O => \N__7942\,
            I => \N__7916\
        );

    \I__1650\ : InMux
    port map (
            O => \N__7941\,
            I => \N__7913\
        );

    \I__1649\ : InMux
    port map (
            O => \N__7940\,
            I => \N__7908\
        );

    \I__1648\ : InMux
    port map (
            O => \N__7939\,
            I => \N__7908\
        );

    \I__1647\ : InMux
    port map (
            O => \N__7938\,
            I => \N__7905\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__7935\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__7932\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__7927\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__7924\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__7919\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__7916\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__7913\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__7908\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__7905\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1637\ : CascadeMux
    port map (
            O => \N__7886\,
            I => \N__7883\
        );

    \I__1636\ : InMux
    port map (
            O => \N__7883\,
            I => \N__7878\
        );

    \I__1635\ : InMux
    port map (
            O => \N__7882\,
            I => \N__7873\
        );

    \I__1634\ : InMux
    port map (
            O => \N__7881\,
            I => \N__7870\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__7878\,
            I => \N__7864\
        );

    \I__1632\ : InMux
    port map (
            O => \N__7877\,
            I => \N__7861\
        );

    \I__1631\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7858\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__7873\,
            I => \N__7847\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__7870\,
            I => \N__7847\
        );

    \I__1628\ : InMux
    port map (
            O => \N__7869\,
            I => \N__7840\
        );

    \I__1627\ : InMux
    port map (
            O => \N__7868\,
            I => \N__7840\
        );

    \I__1626\ : InMux
    port map (
            O => \N__7867\,
            I => \N__7840\
        );

    \I__1625\ : Span4Mux_v
    port map (
            O => \N__7864\,
            I => \N__7832\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__7861\,
            I => \N__7832\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__7858\,
            I => \N__7832\
        );

    \I__1622\ : InMux
    port map (
            O => \N__7857\,
            I => \N__7829\
        );

    \I__1621\ : InMux
    port map (
            O => \N__7856\,
            I => \N__7823\
        );

    \I__1620\ : InMux
    port map (
            O => \N__7855\,
            I => \N__7823\
        );

    \I__1619\ : InMux
    port map (
            O => \N__7854\,
            I => \N__7816\
        );

    \I__1618\ : InMux
    port map (
            O => \N__7853\,
            I => \N__7816\
        );

    \I__1617\ : InMux
    port map (
            O => \N__7852\,
            I => \N__7816\
        );

    \I__1616\ : Span4Mux_v
    port map (
            O => \N__7847\,
            I => \N__7811\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__7840\,
            I => \N__7811\
        );

    \I__1614\ : InMux
    port map (
            O => \N__7839\,
            I => \N__7808\
        );

    \I__1613\ : Span4Mux_h
    port map (
            O => \N__7832\,
            I => \N__7803\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__7829\,
            I => \N__7803\
        );

    \I__1611\ : InMux
    port map (
            O => \N__7828\,
            I => \N__7800\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__7823\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__7816\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1608\ : Odrv4
    port map (
            O => \N__7811\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__7808\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1606\ : Odrv4
    port map (
            O => \N__7803\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__7800\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__7787\,
            I => \U712_CHIP_RAM.N_396_cascade_\
        );

    \I__1603\ : InMux
    port map (
            O => \N__7784\,
            I => \N__7781\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__7781\,
            I => \N__7778\
        );

    \I__1601\ : Span4Mux_v
    port map (
            O => \N__7778\,
            I => \N__7772\
        );

    \I__1600\ : InMux
    port map (
            O => \N__7777\,
            I => \N__7767\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7776\,
            I => \N__7767\
        );

    \I__1598\ : InMux
    port map (
            O => \N__7775\,
            I => \N__7764\
        );

    \I__1597\ : Odrv4
    port map (
            O => \N__7772\,
            I => \U712_CHIP_RAM.N_436\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__7767\,
            I => \U712_CHIP_RAM.N_436\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__7764\,
            I => \U712_CHIP_RAM.N_436\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__7757\,
            I => \U712_CHIP_RAM.N_436_cascade_\
        );

    \I__1593\ : InMux
    port map (
            O => \N__7754\,
            I => \N__7751\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__7751\,
            I => \N__7748\
        );

    \I__1591\ : Span4Mux_h
    port map (
            O => \N__7748\,
            I => \N__7742\
        );

    \I__1590\ : InMux
    port map (
            O => \N__7747\,
            I => \N__7737\
        );

    \I__1589\ : InMux
    port map (
            O => \N__7746\,
            I => \N__7737\
        );

    \I__1588\ : InMux
    port map (
            O => \N__7745\,
            I => \N__7734\
        );

    \I__1587\ : Odrv4
    port map (
            O => \N__7742\,
            I => \U712_CHIP_RAM.N_257\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__7737\,
            I => \U712_CHIP_RAM.N_257\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__7734\,
            I => \U712_CHIP_RAM.N_257\
        );

    \I__1584\ : InMux
    port map (
            O => \N__7727\,
            I => \N__7724\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__7724\,
            I => \N__7721\
        );

    \I__1582\ : Odrv4
    port map (
            O => \N__7721\,
            I => \U712_CHIP_RAM.N_357\
        );

    \I__1581\ : InMux
    port map (
            O => \N__7718\,
            I => \N__7715\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__7715\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0_1\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__7712\,
            I => \N__7708\
        );

    \I__1578\ : InMux
    port map (
            O => \N__7711\,
            I => \N__7704\
        );

    \I__1577\ : InMux
    port map (
            O => \N__7708\,
            I => \N__7700\
        );

    \I__1576\ : CascadeMux
    port map (
            O => \N__7707\,
            I => \N__7697\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__7704\,
            I => \N__7694\
        );

    \I__1574\ : InMux
    port map (
            O => \N__7703\,
            I => \N__7691\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__7700\,
            I => \N__7688\
        );

    \I__1572\ : InMux
    port map (
            O => \N__7697\,
            I => \N__7685\
        );

    \I__1571\ : Span4Mux_v
    port map (
            O => \N__7694\,
            I => \N__7677\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__7691\,
            I => \N__7677\
        );

    \I__1569\ : Span4Mux_v
    port map (
            O => \N__7688\,
            I => \N__7677\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__7685\,
            I => \N__7674\
        );

    \I__1567\ : InMux
    port map (
            O => \N__7684\,
            I => \N__7671\
        );

    \I__1566\ : Odrv4
    port map (
            O => \N__7677\,
            I => \U712_CHIP_RAM.N_396\
        );

    \I__1565\ : Odrv4
    port map (
            O => \N__7674\,
            I => \U712_CHIP_RAM.N_396\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__7671\,
            I => \U712_CHIP_RAM.N_396\
        );

    \I__1563\ : InMux
    port map (
            O => \N__7664\,
            I => \N__7661\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__7661\,
            I => \N__7655\
        );

    \I__1561\ : InMux
    port map (
            O => \N__7660\,
            I => \N__7652\
        );

    \I__1560\ : InMux
    port map (
            O => \N__7659\,
            I => \N__7648\
        );

    \I__1559\ : CascadeMux
    port map (
            O => \N__7658\,
            I => \N__7645\
        );

    \I__1558\ : Span4Mux_h
    port map (
            O => \N__7655\,
            I => \N__7638\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__7652\,
            I => \N__7635\
        );

    \I__1556\ : InMux
    port map (
            O => \N__7651\,
            I => \N__7632\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__7648\,
            I => \N__7629\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7645\,
            I => \N__7626\
        );

    \I__1553\ : InMux
    port map (
            O => \N__7644\,
            I => \N__7621\
        );

    \I__1552\ : InMux
    port map (
            O => \N__7643\,
            I => \N__7621\
        );

    \I__1551\ : InMux
    port map (
            O => \N__7642\,
            I => \N__7616\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7641\,
            I => \N__7616\
        );

    \I__1549\ : Odrv4
    port map (
            O => \N__7638\,
            I => \U712_CHIP_RAM.N_384\
        );

    \I__1548\ : Odrv4
    port map (
            O => \N__7635\,
            I => \U712_CHIP_RAM.N_384\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__7632\,
            I => \U712_CHIP_RAM.N_384\
        );

    \I__1546\ : Odrv4
    port map (
            O => \N__7629\,
            I => \U712_CHIP_RAM.N_384\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__7626\,
            I => \U712_CHIP_RAM.N_384\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__7621\,
            I => \U712_CHIP_RAM.N_384\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__7616\,
            I => \U712_CHIP_RAM.N_384\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7601\,
            I => \N__7598\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__7598\,
            I => \U712_CHIP_RAM.N_351\
        );

    \I__1540\ : CascadeMux
    port map (
            O => \N__7595\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0_cascade_\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7592\,
            I => \N__7589\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7589\,
            I => \U712_CHIP_RAM.N_117\
        );

    \I__1537\ : InMux
    port map (
            O => \N__7586\,
            I => \N__7582\
        );

    \I__1536\ : InMux
    port map (
            O => \N__7585\,
            I => \N__7570\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__7582\,
            I => \N__7567\
        );

    \I__1534\ : InMux
    port map (
            O => \N__7581\,
            I => \N__7564\
        );

    \I__1533\ : InMux
    port map (
            O => \N__7580\,
            I => \N__7561\
        );

    \I__1532\ : InMux
    port map (
            O => \N__7579\,
            I => \N__7558\
        );

    \I__1531\ : InMux
    port map (
            O => \N__7578\,
            I => \N__7555\
        );

    \I__1530\ : InMux
    port map (
            O => \N__7577\,
            I => \N__7550\
        );

    \I__1529\ : InMux
    port map (
            O => \N__7576\,
            I => \N__7550\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7575\,
            I => \N__7543\
        );

    \I__1527\ : InMux
    port map (
            O => \N__7574\,
            I => \N__7543\
        );

    \I__1526\ : InMux
    port map (
            O => \N__7573\,
            I => \N__7543\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__7570\,
            I => \N__7540\
        );

    \I__1524\ : Odrv12
    port map (
            O => \N__7567\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__7564\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7561\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__7558\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__7555\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__7550\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__7543\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1517\ : Odrv4
    port map (
            O => \N__7540\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__7523\,
            I => \N__7520\
        );

    \I__1515\ : InMux
    port map (
            O => \N__7520\,
            I => \N__7516\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7519\,
            I => \N__7511\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__7516\,
            I => \N__7508\
        );

    \I__1512\ : InMux
    port map (
            O => \N__7515\,
            I => \N__7501\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7514\,
            I => \N__7498\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__7511\,
            I => \N__7495\
        );

    \I__1509\ : Span4Mux_v
    port map (
            O => \N__7508\,
            I => \N__7492\
        );

    \I__1508\ : InMux
    port map (
            O => \N__7507\,
            I => \N__7487\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7506\,
            I => \N__7487\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7505\,
            I => \N__7484\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7504\,
            I => \N__7481\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__7501\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7498\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1502\ : Odrv4
    port map (
            O => \N__7495\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__7492\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__7487\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__7484\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__7481\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__7466\,
            I => \N__7457\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7465\,
            I => \N__7451\
        );

    \I__1495\ : InMux
    port map (
            O => \N__7464\,
            I => \N__7446\
        );

    \I__1494\ : InMux
    port map (
            O => \N__7463\,
            I => \N__7446\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7462\,
            I => \N__7442\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7461\,
            I => \N__7439\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7460\,
            I => \N__7436\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7457\,
            I => \N__7433\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7456\,
            I => \N__7428\
        );

    \I__1488\ : InMux
    port map (
            O => \N__7455\,
            I => \N__7428\
        );

    \I__1487\ : InMux
    port map (
            O => \N__7454\,
            I => \N__7425\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__7451\,
            I => \N__7420\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__7446\,
            I => \N__7420\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7445\,
            I => \N__7417\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7442\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__7439\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__7436\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__7433\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7428\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__7425\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1477\ : Odrv4
    port map (
            O => \N__7420\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__7417\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7400\,
            I => \N__7397\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7397\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_63_i_a2_0_0_a2_0_2\
        );

    \I__1473\ : CascadeMux
    port map (
            O => \N__7394\,
            I => \N__7390\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7393\,
            I => \N__7387\
        );

    \I__1471\ : InMux
    port map (
            O => \N__7390\,
            I => \N__7384\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__7387\,
            I => \N__7381\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__7384\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1468\ : Odrv12
    port map (
            O => \N__7381\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1467\ : CascadeMux
    port map (
            O => \N__7376\,
            I => \U712_CYCLE_TERM.N_274_i_0_0_cascade_\
        );

    \I__1466\ : CascadeMux
    port map (
            O => \N__7373\,
            I => \U712_CYCLE_TERM.N_274_i_0_en_cascade_\
        );

    \I__1465\ : CEMux
    port map (
            O => \N__7370\,
            I => \N__7367\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__7367\,
            I => \N__7364\
        );

    \I__1463\ : Span4Mux_h
    port map (
            O => \N__7364\,
            I => \N__7361\
        );

    \I__1462\ : Span4Mux_h
    port map (
            O => \N__7361\,
            I => \N__7358\
        );

    \I__1461\ : Odrv4
    port map (
            O => \N__7358\,
            I => \U712_CYCLE_TERM.N_274_i_0_en_0\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7355\,
            I => \N__7352\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__7352\,
            I => \N__7349\
        );

    \I__1458\ : Span4Mux_h
    port map (
            O => \N__7349\,
            I => \N__7346\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__7346\,
            I => \U712_CHIP_RAM.N_294\
        );

    \I__1456\ : InMux
    port map (
            O => \N__7343\,
            I => \N__7338\
        );

    \I__1455\ : CascadeMux
    port map (
            O => \N__7342\,
            I => \N__7335\
        );

    \I__1454\ : CascadeMux
    port map (
            O => \N__7341\,
            I => \N__7332\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__7338\,
            I => \N__7327\
        );

    \I__1452\ : InMux
    port map (
            O => \N__7335\,
            I => \N__7324\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7332\,
            I => \N__7320\
        );

    \I__1450\ : InMux
    port map (
            O => \N__7331\,
            I => \N__7317\
        );

    \I__1449\ : InMux
    port map (
            O => \N__7330\,
            I => \N__7314\
        );

    \I__1448\ : Span4Mux_v
    port map (
            O => \N__7327\,
            I => \N__7309\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__7324\,
            I => \N__7309\
        );

    \I__1446\ : InMux
    port map (
            O => \N__7323\,
            I => \N__7306\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__7320\,
            I => \N__7301\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__7317\,
            I => \N__7301\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__7314\,
            I => \N__7298\
        );

    \I__1442\ : Span4Mux_h
    port map (
            O => \N__7309\,
            I => \N__7295\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__7306\,
            I => \N__7292\
        );

    \I__1440\ : Span4Mux_h
    port map (
            O => \N__7301\,
            I => \N__7289\
        );

    \I__1439\ : Odrv4
    port map (
            O => \N__7298\,
            I => \DMA_CYCLE\
        );

    \I__1438\ : Odrv4
    port map (
            O => \N__7295\,
            I => \DMA_CYCLE\
        );

    \I__1437\ : Odrv12
    port map (
            O => \N__7292\,
            I => \DMA_CYCLE\
        );

    \I__1436\ : Odrv4
    port map (
            O => \N__7289\,
            I => \DMA_CYCLE\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__7280\,
            I => \U712_CHIP_RAM.N_305_cascade_\
        );

    \I__1434\ : InMux
    port map (
            O => \N__7277\,
            I => \N__7274\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__7274\,
            I => \N__7267\
        );

    \I__1432\ : InMux
    port map (
            O => \N__7273\,
            I => \N__7262\
        );

    \I__1431\ : InMux
    port map (
            O => \N__7272\,
            I => \N__7262\
        );

    \I__1430\ : InMux
    port map (
            O => \N__7271\,
            I => \N__7259\
        );

    \I__1429\ : InMux
    port map (
            O => \N__7270\,
            I => \N__7256\
        );

    \I__1428\ : Odrv4
    port map (
            O => \N__7267\,
            I => \U712_CHIP_RAM.N_388\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__7262\,
            I => \U712_CHIP_RAM.N_388\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__7259\,
            I => \U712_CHIP_RAM.N_388\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__7256\,
            I => \U712_CHIP_RAM.N_388\
        );

    \I__1424\ : CascadeMux
    port map (
            O => \N__7247\,
            I => \N__7242\
        );

    \I__1423\ : CascadeMux
    port map (
            O => \N__7246\,
            I => \N__7238\
        );

    \I__1422\ : InMux
    port map (
            O => \N__7245\,
            I => \N__7233\
        );

    \I__1421\ : InMux
    port map (
            O => \N__7242\,
            I => \N__7229\
        );

    \I__1420\ : InMux
    port map (
            O => \N__7241\,
            I => \N__7226\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7238\,
            I => \N__7223\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__7237\,
            I => \N__7219\
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__7236\,
            I => \N__7216\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__7233\,
            I => \N__7210\
        );

    \I__1415\ : InMux
    port map (
            O => \N__7232\,
            I => \N__7207\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__7229\,
            I => \N__7202\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__7226\,
            I => \N__7202\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__7223\,
            I => \N__7199\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7222\,
            I => \N__7196\
        );

    \I__1410\ : InMux
    port map (
            O => \N__7219\,
            I => \N__7191\
        );

    \I__1409\ : InMux
    port map (
            O => \N__7216\,
            I => \N__7191\
        );

    \I__1408\ : InMux
    port map (
            O => \N__7215\,
            I => \N__7188\
        );

    \I__1407\ : InMux
    port map (
            O => \N__7214\,
            I => \N__7185\
        );

    \I__1406\ : InMux
    port map (
            O => \N__7213\,
            I => \N__7182\
        );

    \I__1405\ : Span4Mux_h
    port map (
            O => \N__7210\,
            I => \N__7179\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__7207\,
            I => \U712_CHIP_RAM.N_45_i\
        );

    \I__1403\ : Odrv4
    port map (
            O => \N__7202\,
            I => \U712_CHIP_RAM.N_45_i\
        );

    \I__1402\ : Odrv4
    port map (
            O => \N__7199\,
            I => \U712_CHIP_RAM.N_45_i\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__7196\,
            I => \U712_CHIP_RAM.N_45_i\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__7191\,
            I => \U712_CHIP_RAM.N_45_i\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__7188\,
            I => \U712_CHIP_RAM.N_45_i\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__7185\,
            I => \U712_CHIP_RAM.N_45_i\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__7182\,
            I => \U712_CHIP_RAM.N_45_i\
        );

    \I__1396\ : Odrv4
    port map (
            O => \N__7179\,
            I => \U712_CHIP_RAM.N_45_i\
        );

    \I__1395\ : CascadeMux
    port map (
            O => \N__7160\,
            I => \U712_CHIP_RAM.N_346_cascade_\
        );

    \I__1394\ : InMux
    port map (
            O => \N__7157\,
            I => \N__7154\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__7154\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_180_i_2\
        );

    \I__1392\ : CascadeMux
    port map (
            O => \N__7151\,
            I => \N__7147\
        );

    \I__1391\ : InMux
    port map (
            O => \N__7150\,
            I => \N__7144\
        );

    \I__1390\ : InMux
    port map (
            O => \N__7147\,
            I => \N__7140\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__7144\,
            I => \N__7137\
        );

    \I__1388\ : InMux
    port map (
            O => \N__7143\,
            I => \N__7134\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__7140\,
            I => \U712_CHIP_RAM.N_407\
        );

    \I__1386\ : Odrv4
    port map (
            O => \N__7137\,
            I => \U712_CHIP_RAM.N_407\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__7134\,
            I => \U712_CHIP_RAM.N_407\
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__7127\,
            I => \U712_CHIP_RAM.N_407_cascade_\
        );

    \I__1383\ : InMux
    port map (
            O => \N__7124\,
            I => \N__7120\
        );

    \I__1382\ : InMux
    port map (
            O => \N__7123\,
            I => \N__7114\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__7120\,
            I => \N__7111\
        );

    \I__1380\ : InMux
    port map (
            O => \N__7119\,
            I => \N__7108\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7118\,
            I => \N__7103\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7117\,
            I => \N__7103\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__7114\,
            I => \U712_CHIP_RAM.N_400\
        );

    \I__1376\ : Odrv4
    port map (
            O => \N__7111\,
            I => \U712_CHIP_RAM.N_400\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__7108\,
            I => \U712_CHIP_RAM.N_400\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__7103\,
            I => \U712_CHIP_RAM.N_400\
        );

    \I__1373\ : InMux
    port map (
            O => \N__7094\,
            I => \N__7090\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__7093\,
            I => \N__7087\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__7090\,
            I => \N__7084\
        );

    \I__1370\ : InMux
    port map (
            O => \N__7087\,
            I => \N__7081\
        );

    \I__1369\ : Span4Mux_v
    port map (
            O => \N__7084\,
            I => \N__7075\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__7081\,
            I => \N__7072\
        );

    \I__1367\ : InMux
    port map (
            O => \N__7080\,
            I => \N__7067\
        );

    \I__1366\ : InMux
    port map (
            O => \N__7079\,
            I => \N__7067\
        );

    \I__1365\ : CascadeMux
    port map (
            O => \N__7078\,
            I => \N__7063\
        );

    \I__1364\ : Span4Mux_v
    port map (
            O => \N__7075\,
            I => \N__7057\
        );

    \I__1363\ : Span4Mux_h
    port map (
            O => \N__7072\,
            I => \N__7057\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__7067\,
            I => \N__7054\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7066\,
            I => \N__7049\
        );

    \I__1360\ : InMux
    port map (
            O => \N__7063\,
            I => \N__7049\
        );

    \I__1359\ : InMux
    port map (
            O => \N__7062\,
            I => \N__7046\
        );

    \I__1358\ : Odrv4
    port map (
            O => \N__7057\,
            I => \WRITE_CYCLE\
        );

    \I__1357\ : Odrv4
    port map (
            O => \N__7054\,
            I => \WRITE_CYCLE\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__7049\,
            I => \WRITE_CYCLE\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__7046\,
            I => \WRITE_CYCLE\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__7037\,
            I => \U712_CHIP_RAM.N_257_cascade_\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__7034\,
            I => \U712_BYTE_ENABLE.UUBE_cascade_\
        );

    \I__1352\ : IoInMux
    port map (
            O => \N__7031\,
            I => \N__7028\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__7028\,
            I => \N__7025\
        );

    \I__1350\ : Span4Mux_s3_h
    port map (
            O => \N__7025\,
            I => \N__7022\
        );

    \I__1349\ : Span4Mux_v
    port map (
            O => \N__7022\,
            I => \N__7019\
        );

    \I__1348\ : Span4Mux_h
    port map (
            O => \N__7019\,
            I => \N__7016\
        );

    \I__1347\ : Span4Mux_h
    port map (
            O => \N__7016\,
            I => \N__7013\
        );

    \I__1346\ : Span4Mux_h
    port map (
            O => \N__7013\,
            I => \N__7010\
        );

    \I__1345\ : Odrv4
    port map (
            O => \N__7010\,
            I => \N_48_i\
        );

    \I__1344\ : CascadeMux
    port map (
            O => \N__7007\,
            I => \N__7004\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7004\,
            I => \N__7001\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__7001\,
            I => \N__6998\
        );

    \I__1341\ : Odrv12
    port map (
            O => \N__6998\,
            I => \U712_BYTE_ENABLE.N_278\
        );

    \I__1340\ : InMux
    port map (
            O => \N__6995\,
            I => \N__6992\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__6992\,
            I => \N__6989\
        );

    \I__1338\ : Odrv4
    port map (
            O => \N__6989\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0Z0Z_0\
        );

    \I__1337\ : IoInMux
    port map (
            O => \N__6986\,
            I => \N__6983\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__6983\,
            I => \N__6980\
        );

    \I__1335\ : Span12Mux_s4_h
    port map (
            O => \N__6980\,
            I => \N__6977\
        );

    \I__1334\ : Span12Mux_h
    port map (
            O => \N__6977\,
            I => \N__6974\
        );

    \I__1333\ : Span12Mux_v
    port map (
            O => \N__6974\,
            I => \N__6971\
        );

    \I__1332\ : Odrv12
    port map (
            O => \N__6971\,
            I => \N_49_i\
        );

    \I__1331\ : CascadeMux
    port map (
            O => \N__6968\,
            I => \N__6965\
        );

    \I__1330\ : InMux
    port map (
            O => \N__6965\,
            I => \N__6962\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__6962\,
            I => \U712_BYTE_ENABLE.N_277\
        );

    \I__1328\ : IoInMux
    port map (
            O => \N__6959\,
            I => \N__6956\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__6956\,
            I => \N__6953\
        );

    \I__1326\ : Span4Mux_s2_v
    port map (
            O => \N__6953\,
            I => \N__6950\
        );

    \I__1325\ : Sp12to4
    port map (
            O => \N__6950\,
            I => \N__6946\
        );

    \I__1324\ : InMux
    port map (
            O => \N__6949\,
            I => \N__6943\
        );

    \I__1323\ : Span12Mux_h
    port map (
            O => \N__6946\,
            I => \N__6938\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__6943\,
            I => \N__6935\
        );

    \I__1321\ : InMux
    port map (
            O => \N__6942\,
            I => \N__6932\
        );

    \I__1320\ : InMux
    port map (
            O => \N__6941\,
            I => \N__6929\
        );

    \I__1319\ : Odrv12
    port map (
            O => \N__6938\,
            I => \DBENn_c\
        );

    \I__1318\ : Odrv4
    port map (
            O => \N__6935\,
            I => \DBENn_c\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__6932\,
            I => \DBENn_c\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__6929\,
            I => \DBENn_c\
        );

    \I__1315\ : InMux
    port map (
            O => \N__6920\,
            I => \N__6914\
        );

    \I__1314\ : InMux
    port map (
            O => \N__6919\,
            I => \N__6914\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__6914\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0Z0Z_0\
        );

    \I__1312\ : InMux
    port map (
            O => \N__6911\,
            I => \N__6908\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__6908\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_2_0\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__6905\,
            I => \U712_CHIP_RAM.N_325_0_cascade_\
        );

    \I__1309\ : InMux
    port map (
            O => \N__6902\,
            I => \N__6899\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__6899\,
            I => \N__6896\
        );

    \I__1307\ : Odrv4
    port map (
            O => \N__6896\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0\
        );

    \I__1306\ : CascadeMux
    port map (
            O => \N__6893\,
            I => \N__6890\
        );

    \I__1305\ : InMux
    port map (
            O => \N__6890\,
            I => \N__6887\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__6887\,
            I => \N__6884\
        );

    \I__1303\ : Span4Mux_h
    port map (
            O => \N__6884\,
            I => \N__6881\
        );

    \I__1302\ : Odrv4
    port map (
            O => \N__6881\,
            I => \U712_CHIP_RAM.N_365_1\
        );

    \I__1301\ : IoInMux
    port map (
            O => \N__6878\,
            I => \N__6875\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__6875\,
            I => \N__6872\
        );

    \I__1299\ : Span4Mux_s2_v
    port map (
            O => \N__6872\,
            I => \N__6869\
        );

    \I__1298\ : Span4Mux_v
    port map (
            O => \N__6869\,
            I => \N__6866\
        );

    \I__1297\ : Odrv4
    port map (
            O => \N__6866\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1296\ : InMux
    port map (
            O => \N__6863\,
            I => \N__6860\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__6860\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__1294\ : IoInMux
    port map (
            O => \N__6857\,
            I => \N__6854\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__6854\,
            I => \N__6851\
        );

    \I__1292\ : Span4Mux_s3_h
    port map (
            O => \N__6851\,
            I => \N__6848\
        );

    \I__1291\ : Span4Mux_v
    port map (
            O => \N__6848\,
            I => \N__6845\
        );

    \I__1290\ : Sp12to4
    port map (
            O => \N__6845\,
            I => \N__6842\
        );

    \I__1289\ : Span12Mux_h
    port map (
            O => \N__6842\,
            I => \N__6839\
        );

    \I__1288\ : Odrv12
    port map (
            O => \N__6839\,
            I => \CMA_c_7\
        );

    \I__1287\ : InMux
    port map (
            O => \N__6836\,
            I => \N__6833\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__6833\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__1285\ : IoInMux
    port map (
            O => \N__6830\,
            I => \N__6827\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__6827\,
            I => \N__6824\
        );

    \I__1283\ : IoSpan4Mux
    port map (
            O => \N__6824\,
            I => \N__6821\
        );

    \I__1282\ : Sp12to4
    port map (
            O => \N__6821\,
            I => \N__6818\
        );

    \I__1281\ : Span12Mux_s9_h
    port map (
            O => \N__6818\,
            I => \N__6815\
        );

    \I__1280\ : Span12Mux_v
    port map (
            O => \N__6815\,
            I => \N__6812\
        );

    \I__1279\ : Odrv12
    port map (
            O => \N__6812\,
            I => \CMA_c_4\
        );

    \I__1278\ : InMux
    port map (
            O => \N__6809\,
            I => \N__6806\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6806\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1276\ : IoInMux
    port map (
            O => \N__6803\,
            I => \N__6800\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__6800\,
            I => \N__6797\
        );

    \I__1274\ : IoSpan4Mux
    port map (
            O => \N__6797\,
            I => \N__6794\
        );

    \I__1273\ : Span4Mux_s2_h
    port map (
            O => \N__6794\,
            I => \N__6791\
        );

    \I__1272\ : Sp12to4
    port map (
            O => \N__6791\,
            I => \N__6788\
        );

    \I__1271\ : Span12Mux_h
    port map (
            O => \N__6788\,
            I => \N__6785\
        );

    \I__1270\ : Odrv12
    port map (
            O => \N__6785\,
            I => \CMA_c_3\
        );

    \I__1269\ : InMux
    port map (
            O => \N__6782\,
            I => \N__6779\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__6779\,
            I => \N__6776\
        );

    \I__1267\ : Odrv4
    port map (
            O => \N__6776\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__1266\ : IoInMux
    port map (
            O => \N__6773\,
            I => \N__6770\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6770\,
            I => \N__6767\
        );

    \I__1264\ : IoSpan4Mux
    port map (
            O => \N__6767\,
            I => \N__6764\
        );

    \I__1263\ : Span4Mux_s3_h
    port map (
            O => \N__6764\,
            I => \N__6761\
        );

    \I__1262\ : Span4Mux_v
    port map (
            O => \N__6761\,
            I => \N__6758\
        );

    \I__1261\ : Span4Mux_v
    port map (
            O => \N__6758\,
            I => \N__6755\
        );

    \I__1260\ : Sp12to4
    port map (
            O => \N__6755\,
            I => \N__6752\
        );

    \I__1259\ : Odrv12
    port map (
            O => \N__6752\,
            I => \CMA_c_6\
        );

    \I__1258\ : InMux
    port map (
            O => \N__6749\,
            I => \N__6746\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__6746\,
            I => \N__6743\
        );

    \I__1256\ : Span12Mux_v
    port map (
            O => \N__6743\,
            I => \N__6740\
        );

    \I__1255\ : Span12Mux_h
    port map (
            O => \N__6740\,
            I => \N__6737\
        );

    \I__1254\ : Odrv12
    port map (
            O => \N__6737\,
            I => \A_c_19\
        );

    \I__1253\ : IoInMux
    port map (
            O => \N__6734\,
            I => \N__6731\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__6731\,
            I => \N__6728\
        );

    \I__1251\ : Span12Mux_s4_h
    port map (
            O => \N__6728\,
            I => \N__6725\
        );

    \I__1250\ : Span12Mux_h
    port map (
            O => \N__6725\,
            I => \N__6722\
        );

    \I__1249\ : Odrv12
    port map (
            O => \N__6722\,
            I => \CMA_c_9\
        );

    \I__1248\ : InMux
    port map (
            O => \N__6719\,
            I => \N__6716\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__6716\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__1246\ : IoInMux
    port map (
            O => \N__6713\,
            I => \N__6710\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__6710\,
            I => \N__6707\
        );

    \I__1244\ : Span4Mux_s1_v
    port map (
            O => \N__6707\,
            I => \N__6704\
        );

    \I__1243\ : Span4Mux_v
    port map (
            O => \N__6704\,
            I => \N__6701\
        );

    \I__1242\ : Span4Mux_v
    port map (
            O => \N__6701\,
            I => \N__6698\
        );

    \I__1241\ : Span4Mux_v
    port map (
            O => \N__6698\,
            I => \N__6695\
        );

    \I__1240\ : Odrv4
    port map (
            O => \N__6695\,
            I => \CMA_c_2\
        );

    \I__1239\ : IoInMux
    port map (
            O => \N__6692\,
            I => \N__6689\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6689\,
            I => \N__6686\
        );

    \I__1237\ : Span4Mux_s0_h
    port map (
            O => \N__6686\,
            I => \N__6683\
        );

    \I__1236\ : Span4Mux_h
    port map (
            O => \N__6683\,
            I => \N__6680\
        );

    \I__1235\ : Sp12to4
    port map (
            O => \N__6680\,
            I => \N__6677\
        );

    \I__1234\ : Span12Mux_s10_v
    port map (
            O => \N__6677\,
            I => \N__6674\
        );

    \I__1233\ : Span12Mux_h
    port map (
            O => \N__6674\,
            I => \N__6671\
        );

    \I__1232\ : Odrv12
    port map (
            O => \N__6671\,
            I => \N_46_i\
        );

    \I__1231\ : InMux
    port map (
            O => \N__6668\,
            I => \N__6665\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__6665\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0_0\
        );

    \I__1229\ : CascadeMux
    port map (
            O => \N__6662\,
            I => \N__6657\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__6661\,
            I => \N__6650\
        );

    \I__1227\ : InMux
    port map (
            O => \N__6660\,
            I => \N__6645\
        );

    \I__1226\ : InMux
    port map (
            O => \N__6657\,
            I => \N__6642\
        );

    \I__1225\ : InMux
    port map (
            O => \N__6656\,
            I => \N__6635\
        );

    \I__1224\ : InMux
    port map (
            O => \N__6655\,
            I => \N__6635\
        );

    \I__1223\ : InMux
    port map (
            O => \N__6654\,
            I => \N__6635\
        );

    \I__1222\ : InMux
    port map (
            O => \N__6653\,
            I => \N__6632\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6650\,
            I => \N__6627\
        );

    \I__1220\ : InMux
    port map (
            O => \N__6649\,
            I => \N__6627\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6648\,
            I => \N__6624\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__6645\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__6642\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__6635\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__6632\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__6627\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__6624\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1212\ : CascadeMux
    port map (
            O => \N__6611\,
            I => \N__6608\
        );

    \I__1211\ : InMux
    port map (
            O => \N__6608\,
            I => \N__6605\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__6605\,
            I => \N__6602\
        );

    \I__1209\ : Odrv4
    port map (
            O => \N__6602\,
            I => \U712_CHIP_RAM.N_444\
        );

    \I__1208\ : CascadeMux
    port map (
            O => \N__6599\,
            I => \N__6596\
        );

    \I__1207\ : InMux
    port map (
            O => \N__6596\,
            I => \N__6592\
        );

    \I__1206\ : InMux
    port map (
            O => \N__6595\,
            I => \N__6589\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__6592\,
            I => \N__6586\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__6589\,
            I => \N__6583\
        );

    \I__1203\ : Span4Mux_h
    port map (
            O => \N__6586\,
            I => \N__6579\
        );

    \I__1202\ : Span4Mux_h
    port map (
            O => \N__6583\,
            I => \N__6576\
        );

    \I__1201\ : InMux
    port map (
            O => \N__6582\,
            I => \N__6573\
        );

    \I__1200\ : Odrv4
    port map (
            O => \N__6579\,
            I => \U712_CHIP_RAM.N_392\
        );

    \I__1199\ : Odrv4
    port map (
            O => \N__6576\,
            I => \U712_CHIP_RAM.N_392\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__6573\,
            I => \U712_CHIP_RAM.N_392\
        );

    \I__1197\ : CascadeMux
    port map (
            O => \N__6566\,
            I => \U712_CHIP_RAM.N_444_cascade_\
        );

    \I__1196\ : InMux
    port map (
            O => \N__6563\,
            I => \N__6560\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__6560\,
            I => \N__6556\
        );

    \I__1194\ : InMux
    port map (
            O => \N__6559\,
            I => \N__6553\
        );

    \I__1193\ : Odrv12
    port map (
            O => \N__6556\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__6553\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6548\,
            I => \N__6545\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__6545\,
            I => \N__6542\
        );

    \I__1189\ : Odrv4
    port map (
            O => \N__6542\,
            I => \U712_CHIP_RAM.N_334\
        );

    \I__1188\ : CascadeMux
    port map (
            O => \N__6539\,
            I => \U712_CHIP_RAM.N_334_cascade_\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6536\,
            I => \N__6533\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__6533\,
            I => \N__6530\
        );

    \I__1185\ : Odrv12
    port map (
            O => \N__6530\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0\
        );

    \I__1184\ : CascadeMux
    port map (
            O => \N__6527\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_cascade_\
        );

    \I__1183\ : CEMux
    port map (
            O => \N__6524\,
            I => \N__6521\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__6521\,
            I => \N__6518\
        );

    \I__1181\ : Span4Mux_h
    port map (
            O => \N__6518\,
            I => \N__6515\
        );

    \I__1180\ : Odrv4
    port map (
            O => \N__6515\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_0\
        );

    \I__1179\ : CascadeMux
    port map (
            O => \N__6512\,
            I => \N__6508\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__6511\,
            I => \N__6505\
        );

    \I__1177\ : InMux
    port map (
            O => \N__6508\,
            I => \N__6502\
        );

    \I__1176\ : InMux
    port map (
            O => \N__6505\,
            I => \N__6499\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6502\,
            I => \U712_CHIP_RAM.N_448\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__6499\,
            I => \U712_CHIP_RAM.N_448\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6494\,
            I => \N__6491\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__6491\,
            I => \U712_CHIP_RAM.N_323\
        );

    \I__1171\ : CascadeMux
    port map (
            O => \N__6488\,
            I => \U712_CHIP_RAM.N_323_cascade_\
        );

    \I__1170\ : InMux
    port map (
            O => \N__6485\,
            I => \N__6482\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__6482\,
            I => \N__6479\
        );

    \I__1168\ : Odrv4
    port map (
            O => \N__6479\,
            I => \U712_CHIP_RAM.un3_DMA_CYCLE_START\
        );

    \I__1167\ : InMux
    port map (
            O => \N__6476\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__1166\ : InMux
    port map (
            O => \N__6473\,
            I => \N__6470\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6470\,
            I => \N__6467\
        );

    \I__1164\ : Odrv4
    port map (
            O => \N__6467\,
            I => \U712_CHIP_RAM.N_363\
        );

    \I__1163\ : InMux
    port map (
            O => \N__6464\,
            I => \N__6460\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6463\,
            I => \N__6457\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__6460\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__6457\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6452\,
            I => \N__6448\
        );

    \I__1158\ : InMux
    port map (
            O => \N__6451\,
            I => \N__6445\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__6448\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__6445\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6440\,
            I => \N__6436\
        );

    \I__1154\ : InMux
    port map (
            O => \N__6439\,
            I => \N__6433\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__6436\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__6433\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1151\ : CascadeMux
    port map (
            O => \N__6428\,
            I => \U712_CHIP_RAM.N_384_cascade_\
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__6425\,
            I => \U712_CHIP_RAM.N_448_cascade_\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6422\,
            I => \N__6419\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__6419\,
            I => \U712_CHIP_RAM.N_255\
        );

    \I__1147\ : CascadeMux
    port map (
            O => \N__6416\,
            I => \U712_CHIP_RAM.N_255_cascade_\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6413\,
            I => \N__6410\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__6410\,
            I => \U712_CHIP_RAM.N_269\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__6407\,
            I => \N__6404\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6404\,
            I => \N__6401\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__6401\,
            I => \N__6394\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6400\,
            I => \N__6391\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6399\,
            I => \N__6386\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6398\,
            I => \N__6386\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6397\,
            I => \N__6383\
        );

    \I__1137\ : Odrv4
    port map (
            O => \N__6394\,
            I => \U712_CHIP_RAM.N_324\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6391\,
            I => \U712_CHIP_RAM.N_324\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__6386\,
            I => \U712_CHIP_RAM.N_324\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__6383\,
            I => \U712_CHIP_RAM.N_324\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__6374\,
            I => \U712_CHIP_RAM.N_456_cascade_\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6371\,
            I => \N__6365\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6370\,
            I => \N__6362\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6369\,
            I => \N__6357\
        );

    \I__1129\ : InMux
    port map (
            O => \N__6368\,
            I => \N__6357\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__6365\,
            I => \N__6352\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__6362\,
            I => \N__6352\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__6357\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1\
        );

    \I__1125\ : Odrv4
    port map (
            O => \N__6352\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1\
        );

    \I__1124\ : InMux
    port map (
            O => \N__6347\,
            I => \bfn_11_11_0_\
        );

    \I__1123\ : InMux
    port map (
            O => \N__6344\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__1122\ : InMux
    port map (
            O => \N__6341\,
            I => \N__6338\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__6338\,
            I => \N__6334\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6337\,
            I => \N__6331\
        );

    \I__1119\ : Odrv4
    port map (
            O => \N__6334\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6331\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6326\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6323\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6320\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__1114\ : InMux
    port map (
            O => \N__6317\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__1113\ : InMux
    port map (
            O => \N__6314\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__1112\ : CascadeMux
    port map (
            O => \N__6311\,
            I => \N__6308\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6308\,
            I => \N__6305\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6305\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__6302\,
            I => \U712_CHIP_RAM.CMA_5_0_8_cascade_\
        );

    \I__1108\ : InMux
    port map (
            O => \N__6299\,
            I => \N__6296\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__6296\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__1106\ : InMux
    port map (
            O => \N__6293\,
            I => \N__6290\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__6290\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\
        );

    \I__1104\ : InMux
    port map (
            O => \N__6287\,
            I => \N__6281\
        );

    \I__1103\ : InMux
    port map (
            O => \N__6286\,
            I => \N__6281\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__6281\,
            I => \N__6278\
        );

    \I__1101\ : Span4Mux_v
    port map (
            O => \N__6278\,
            I => \N__6275\
        );

    \I__1100\ : Sp12to4
    port map (
            O => \N__6275\,
            I => \N__6272\
        );

    \I__1099\ : Span12Mux_h
    port map (
            O => \N__6272\,
            I => \N__6269\
        );

    \I__1098\ : Odrv12
    port map (
            O => \N__6269\,
            I => \A_c_10\
        );

    \I__1097\ : InMux
    port map (
            O => \N__6266\,
            I => \N__6263\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__6263\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6260\,
            I => \N__6257\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6257\,
            I => \N__6253\
        );

    \I__1093\ : InMux
    port map (
            O => \N__6256\,
            I => \N__6250\
        );

    \I__1092\ : Span4Mux_v
    port map (
            O => \N__6253\,
            I => \N__6245\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__6250\,
            I => \N__6245\
        );

    \I__1090\ : Span4Mux_v
    port map (
            O => \N__6245\,
            I => \N__6242\
        );

    \I__1089\ : Sp12to4
    port map (
            O => \N__6242\,
            I => \N__6239\
        );

    \I__1088\ : Span12Mux_h
    port map (
            O => \N__6239\,
            I => \N__6236\
        );

    \I__1087\ : Odrv12
    port map (
            O => \N__6236\,
            I => \AWEn_c\
        );

    \I__1086\ : IoInMux
    port map (
            O => \N__6233\,
            I => \N__6230\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__6230\,
            I => \N__6227\
        );

    \I__1084\ : Span4Mux_s2_v
    port map (
            O => \N__6227\,
            I => \N__6224\
        );

    \I__1083\ : Span4Mux_h
    port map (
            O => \N__6224\,
            I => \N__6220\
        );

    \I__1082\ : CascadeMux
    port map (
            O => \N__6223\,
            I => \N__6217\
        );

    \I__1081\ : Sp12to4
    port map (
            O => \N__6220\,
            I => \N__6214\
        );

    \I__1080\ : InMux
    port map (
            O => \N__6217\,
            I => \N__6211\
        );

    \I__1079\ : Odrv12
    port map (
            O => \N__6214\,
            I => \DBDIR_c\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__6211\,
            I => \DBDIR_c\
        );

    \I__1077\ : InMux
    port map (
            O => \N__6206\,
            I => \N__6202\
        );

    \I__1076\ : InMux
    port map (
            O => \N__6205\,
            I => \N__6199\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__6202\,
            I => \N__6196\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__6199\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1073\ : Odrv12
    port map (
            O => \N__6196\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6191\,
            I => \N__6187\
        );

    \I__1071\ : InMux
    port map (
            O => \N__6190\,
            I => \N__6184\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__6187\,
            I => \N__6181\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__6184\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1068\ : Odrv4
    port map (
            O => \N__6181\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1067\ : CascadeMux
    port map (
            O => \N__6176\,
            I => \N__6173\
        );

    \I__1066\ : InMux
    port map (
            O => \N__6173\,
            I => \N__6169\
        );

    \I__1065\ : InMux
    port map (
            O => \N__6172\,
            I => \N__6166\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__6169\,
            I => \N__6163\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__6166\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1062\ : Odrv12
    port map (
            O => \N__6163\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1061\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6155\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__6155\,
            I => \N__6152\
        );

    \I__1059\ : Odrv4
    port map (
            O => \N__6152\,
            I => \U712_CHIP_RAM.REFRESH5lt7\
        );

    \I__1058\ : CascadeMux
    port map (
            O => \N__6149\,
            I => \N__6144\
        );

    \I__1057\ : InMux
    port map (
            O => \N__6148\,
            I => \N__6140\
        );

    \I__1056\ : InMux
    port map (
            O => \N__6147\,
            I => \N__6137\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6144\,
            I => \N__6134\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6143\,
            I => \N__6130\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__6140\,
            I => \N__6127\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6137\,
            I => \N__6123\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__6134\,
            I => \N__6120\
        );

    \I__1050\ : InMux
    port map (
            O => \N__6133\,
            I => \N__6117\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__6130\,
            I => \N__6112\
        );

    \I__1048\ : Span4Mux_v
    port map (
            O => \N__6127\,
            I => \N__6112\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6126\,
            I => \N__6109\
        );

    \I__1046\ : Span4Mux_h
    port map (
            O => \N__6123\,
            I => \N__6106\
        );

    \I__1045\ : Span4Mux_h
    port map (
            O => \N__6120\,
            I => \N__6101\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__6117\,
            I => \N__6101\
        );

    \I__1043\ : Odrv4
    port map (
            O => \N__6112\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__6109\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1041\ : Odrv4
    port map (
            O => \N__6106\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1040\ : Odrv4
    port map (
            O => \N__6101\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6092\,
            I => \N__6089\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__6089\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\
        );

    \I__1037\ : InMux
    port map (
            O => \N__6086\,
            I => \N__6083\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__6083\,
            I => \N__6079\
        );

    \I__1035\ : InMux
    port map (
            O => \N__6082\,
            I => \N__6076\
        );

    \I__1034\ : Odrv4
    port map (
            O => \N__6079\,
            I => \LATCH_RAM\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__6076\,
            I => \LATCH_RAM\
        );

    \I__1032\ : InMux
    port map (
            O => \N__6071\,
            I => \N__6068\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__6068\,
            I => \N__6064\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6067\,
            I => \N__6061\
        );

    \I__1029\ : Odrv12
    port map (
            O => \N__6064\,
            I => \U712_REG_SM.N_265\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__6061\,
            I => \U712_REG_SM.N_265\
        );

    \I__1027\ : InMux
    port map (
            O => \N__6056\,
            I => \N__6053\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__6053\,
            I => \N__6050\
        );

    \I__1025\ : Span4Mux_h
    port map (
            O => \N__6050\,
            I => \N__6044\
        );

    \I__1024\ : InMux
    port map (
            O => \N__6049\,
            I => \N__6041\
        );

    \I__1023\ : InMux
    port map (
            O => \N__6048\,
            I => \N__6038\
        );

    \I__1022\ : InMux
    port map (
            O => \N__6047\,
            I => \N__6035\
        );

    \I__1021\ : Odrv4
    port map (
            O => \N__6044\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_1\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__6041\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_1\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__6038\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_1\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__6035\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_1\
        );

    \I__1017\ : InMux
    port map (
            O => \N__6026\,
            I => \N__6019\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6025\,
            I => \N__6016\
        );

    \I__1015\ : CascadeMux
    port map (
            O => \N__6024\,
            I => \N__6013\
        );

    \I__1014\ : InMux
    port map (
            O => \N__6023\,
            I => \N__6008\
        );

    \I__1013\ : InMux
    port map (
            O => \N__6022\,
            I => \N__6005\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__6019\,
            I => \N__6000\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__6016\,
            I => \N__6000\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6013\,
            I => \N__5994\
        );

    \I__1009\ : InMux
    port map (
            O => \N__6012\,
            I => \N__5991\
        );

    \I__1008\ : InMux
    port map (
            O => \N__6011\,
            I => \N__5988\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__6008\,
            I => \N__5983\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__6005\,
            I => \N__5983\
        );

    \I__1005\ : Span4Mux_h
    port map (
            O => \N__6000\,
            I => \N__5980\
        );

    \I__1004\ : InMux
    port map (
            O => \N__5999\,
            I => \N__5973\
        );

    \I__1003\ : InMux
    port map (
            O => \N__5998\,
            I => \N__5973\
        );

    \I__1002\ : InMux
    port map (
            O => \N__5997\,
            I => \N__5973\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__5994\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__5991\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__5988\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__998\ : Odrv4
    port map (
            O => \N__5983\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__997\ : Odrv4
    port map (
            O => \N__5980\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5973\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__995\ : InMux
    port map (
            O => \N__5960\,
            I => \N__5955\
        );

    \I__994\ : InMux
    port map (
            O => \N__5959\,
            I => \N__5952\
        );

    \I__993\ : InMux
    port map (
            O => \N__5958\,
            I => \N__5949\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__5955\,
            I => \U712_REG_SM.DBR_SYNCZ0Z_1\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__5952\,
            I => \U712_REG_SM.DBR_SYNCZ0Z_1\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__5949\,
            I => \U712_REG_SM.DBR_SYNCZ0Z_1\
        );

    \I__989\ : InMux
    port map (
            O => \N__5942\,
            I => \N__5939\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__5939\,
            I => \N__5935\
        );

    \I__987\ : InMux
    port map (
            O => \N__5938\,
            I => \N__5932\
        );

    \I__986\ : Span4Mux_v
    port map (
            O => \N__5935\,
            I => \N__5926\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__5932\,
            I => \N__5926\
        );

    \I__984\ : InMux
    port map (
            O => \N__5931\,
            I => \N__5923\
        );

    \I__983\ : Span4Mux_h
    port map (
            O => \N__5926\,
            I => \N__5918\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__5923\,
            I => \N__5918\
        );

    \I__981\ : Span4Mux_v
    port map (
            O => \N__5918\,
            I => \N__5915\
        );

    \I__980\ : Sp12to4
    port map (
            O => \N__5915\,
            I => \N__5912\
        );

    \I__979\ : Span12Mux_h
    port map (
            O => \N__5912\,
            I => \N__5909\
        );

    \I__978\ : Odrv12
    port map (
            O => \N__5909\,
            I => \DBRn_c\
        );

    \I__977\ : InMux
    port map (
            O => \N__5906\,
            I => \N__5903\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__5903\,
            I => \U712_REG_SM.DBR_SYNCZ0Z_0\
        );

    \I__975\ : InMux
    port map (
            O => \N__5900\,
            I => \N__5897\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__5897\,
            I => \N__5894\
        );

    \I__973\ : Span4Mux_v
    port map (
            O => \N__5894\,
            I => \N__5886\
        );

    \I__972\ : InMux
    port map (
            O => \N__5893\,
            I => \N__5881\
        );

    \I__971\ : InMux
    port map (
            O => \N__5892\,
            I => \N__5881\
        );

    \I__970\ : InMux
    port map (
            O => \N__5891\,
            I => \N__5874\
        );

    \I__969\ : InMux
    port map (
            O => \N__5890\,
            I => \N__5874\
        );

    \I__968\ : InMux
    port map (
            O => \N__5889\,
            I => \N__5874\
        );

    \I__967\ : Odrv4
    port map (
            O => \N__5886\,
            I => \REG_WRITE_CYCLE\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5881\,
            I => \REG_WRITE_CYCLE\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__5874\,
            I => \REG_WRITE_CYCLE\
        );

    \I__964\ : IoInMux
    port map (
            O => \N__5867\,
            I => \N__5864\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__5864\,
            I => \N__5860\
        );

    \I__962\ : IoInMux
    port map (
            O => \N__5863\,
            I => \N__5857\
        );

    \I__961\ : IoSpan4Mux
    port map (
            O => \N__5860\,
            I => \N__5854\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__5857\,
            I => \N__5851\
        );

    \I__959\ : Span4Mux_s3_h
    port map (
            O => \N__5854\,
            I => \N__5848\
        );

    \I__958\ : IoSpan4Mux
    port map (
            O => \N__5851\,
            I => \N__5845\
        );

    \I__957\ : Span4Mux_h
    port map (
            O => \N__5848\,
            I => \N__5842\
        );

    \I__956\ : Span4Mux_s2_v
    port map (
            O => \N__5845\,
            I => \N__5839\
        );

    \I__955\ : Sp12to4
    port map (
            O => \N__5842\,
            I => \N__5836\
        );

    \I__954\ : Sp12to4
    port map (
            O => \N__5839\,
            I => \N__5833\
        );

    \I__953\ : Span12Mux_h
    port map (
            O => \N__5836\,
            I => \N__5830\
        );

    \I__952\ : Span12Mux_s10_v
    port map (
            O => \N__5833\,
            I => \N__5827\
        );

    \I__951\ : Odrv12
    port map (
            O => \N__5830\,
            I => \N_289\
        );

    \I__950\ : Odrv12
    port map (
            O => \N__5827\,
            I => \N_289\
        );

    \I__949\ : InMux
    port map (
            O => \N__5822\,
            I => \N__5819\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__5819\,
            I => \N__5816\
        );

    \I__947\ : Sp12to4
    port map (
            O => \N__5816\,
            I => \N__5813\
        );

    \I__946\ : Span12Mux_v
    port map (
            O => \N__5813\,
            I => \N__5810\
        );

    \I__945\ : Span12Mux_h
    port map (
            O => \N__5810\,
            I => \N__5807\
        );

    \I__944\ : Odrv12
    port map (
            O => \N__5807\,
            I => \A_c_5\
        );

    \I__943\ : InMux
    port map (
            O => \N__5804\,
            I => \N__5801\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__5801\,
            I => \N__5798\
        );

    \I__941\ : Span4Mux_v
    port map (
            O => \N__5798\,
            I => \N__5795\
        );

    \I__940\ : Sp12to4
    port map (
            O => \N__5795\,
            I => \N__5792\
        );

    \I__939\ : Span12Mux_h
    port map (
            O => \N__5792\,
            I => \N__5789\
        );

    \I__938\ : Odrv12
    port map (
            O => \N__5789\,
            I => \A_c_12\
        );

    \I__937\ : CascadeMux
    port map (
            O => \N__5786\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\
        );

    \I__936\ : InMux
    port map (
            O => \N__5783\,
            I => \N__5780\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__5780\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\
        );

    \I__934\ : CascadeMux
    port map (
            O => \N__5777\,
            I => \U712_CHIP_RAM.N_365_1_cascade_\
        );

    \I__933\ : CascadeMux
    port map (
            O => \N__5774\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_\
        );

    \I__932\ : CEMux
    port map (
            O => \N__5771\,
            I => \N__5768\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__5768\,
            I => \N__5765\
        );

    \I__930\ : Span4Mux_h
    port map (
            O => \N__5765\,
            I => \N__5762\
        );

    \I__929\ : Odrv4
    port map (
            O => \N__5762\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0\
        );

    \I__928\ : InMux
    port map (
            O => \N__5759\,
            I => \N__5753\
        );

    \I__927\ : CascadeMux
    port map (
            O => \N__5758\,
            I => \N__5750\
        );

    \I__926\ : InMux
    port map (
            O => \N__5757\,
            I => \N__5747\
        );

    \I__925\ : InMux
    port map (
            O => \N__5756\,
            I => \N__5744\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__5753\,
            I => \N__5741\
        );

    \I__923\ : InMux
    port map (
            O => \N__5750\,
            I => \N__5738\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__5747\,
            I => \N__5735\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__5744\,
            I => \N__5732\
        );

    \I__920\ : Span4Mux_h
    port map (
            O => \N__5741\,
            I => \N__5727\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__5738\,
            I => \N__5727\
        );

    \I__918\ : Sp12to4
    port map (
            O => \N__5735\,
            I => \N__5724\
        );

    \I__917\ : Span4Mux_v
    port map (
            O => \N__5732\,
            I => \N__5719\
        );

    \I__916\ : Span4Mux_v
    port map (
            O => \N__5727\,
            I => \N__5719\
        );

    \I__915\ : Span12Mux_v
    port map (
            O => \N__5724\,
            I => \N__5716\
        );

    \I__914\ : Sp12to4
    port map (
            O => \N__5719\,
            I => \N__5713\
        );

    \I__913\ : Span12Mux_h
    port map (
            O => \N__5716\,
            I => \N__5710\
        );

    \I__912\ : Span12Mux_h
    port map (
            O => \N__5713\,
            I => \N__5707\
        );

    \I__911\ : Odrv12
    port map (
            O => \N__5710\,
            I => \RnW_c\
        );

    \I__910\ : Odrv12
    port map (
            O => \N__5707\,
            I => \RnW_c\
        );

    \I__909\ : IoInMux
    port map (
            O => \N__5702\,
            I => \N__5699\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__5699\,
            I => \N__5696\
        );

    \I__907\ : IoSpan4Mux
    port map (
            O => \N__5696\,
            I => \N__5693\
        );

    \I__906\ : Span4Mux_s3_h
    port map (
            O => \N__5693\,
            I => \N__5690\
        );

    \I__905\ : Span4Mux_h
    port map (
            O => \N__5690\,
            I => \N__5687\
        );

    \I__904\ : Sp12to4
    port map (
            O => \N__5687\,
            I => \N__5684\
        );

    \I__903\ : Span12Mux_h
    port map (
            O => \N__5684\,
            I => \N__5680\
        );

    \I__902\ : InMux
    port map (
            O => \N__5683\,
            I => \N__5677\
        );

    \I__901\ : Odrv12
    port map (
            O => \N__5680\,
            I => \CLK_EN_c\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__5677\,
            I => \CLK_EN_c\
        );

    \I__899\ : InMux
    port map (
            O => \N__5672\,
            I => \N__5669\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__5669\,
            I => \N__5666\
        );

    \I__897\ : Span12Mux_h
    port map (
            O => \N__5666\,
            I => \N__5663\
        );

    \I__896\ : Span12Mux_v
    port map (
            O => \N__5663\,
            I => \N__5660\
        );

    \I__895\ : Odrv12
    port map (
            O => \N__5660\,
            I => \RAMSPACEn_c\
        );

    \I__894\ : CascadeMux
    port map (
            O => \N__5657\,
            I => \N__5654\
        );

    \I__893\ : InMux
    port map (
            O => \N__5654\,
            I => \N__5650\
        );

    \I__892\ : CascadeMux
    port map (
            O => \N__5653\,
            I => \N__5647\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__5650\,
            I => \N__5644\
        );

    \I__890\ : InMux
    port map (
            O => \N__5647\,
            I => \N__5641\
        );

    \I__889\ : Span4Mux_h
    port map (
            O => \N__5644\,
            I => \N__5636\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__5641\,
            I => \N__5636\
        );

    \I__887\ : Span4Mux_v
    port map (
            O => \N__5636\,
            I => \N__5633\
        );

    \I__886\ : Sp12to4
    port map (
            O => \N__5633\,
            I => \N__5630\
        );

    \I__885\ : Span12Mux_h
    port map (
            O => \N__5630\,
            I => \N__5627\
        );

    \I__884\ : Odrv12
    port map (
            O => \N__5627\,
            I => \TSn_c\
        );

    \I__883\ : InMux
    port map (
            O => \N__5624\,
            I => \N__5617\
        );

    \I__882\ : CascadeMux
    port map (
            O => \N__5623\,
            I => \N__5614\
        );

    \I__881\ : InMux
    port map (
            O => \N__5622\,
            I => \N__5611\
        );

    \I__880\ : InMux
    port map (
            O => \N__5621\,
            I => \N__5608\
        );

    \I__879\ : InMux
    port map (
            O => \N__5620\,
            I => \N__5605\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__5617\,
            I => \N__5602\
        );

    \I__877\ : InMux
    port map (
            O => \N__5614\,
            I => \N__5599\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__5611\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5608\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__5605\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__873\ : Odrv4
    port map (
            O => \N__5602\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__5599\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__871\ : InMux
    port map (
            O => \N__5588\,
            I => \N__5584\
        );

    \I__870\ : InMux
    port map (
            O => \N__5587\,
            I => \N__5579\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__5584\,
            I => \N__5576\
        );

    \I__868\ : InMux
    port map (
            O => \N__5583\,
            I => \N__5573\
        );

    \I__867\ : InMux
    port map (
            O => \N__5582\,
            I => \N__5570\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5579\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__865\ : Odrv4
    port map (
            O => \N__5576\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__5573\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__5570\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__862\ : InMux
    port map (
            O => \N__5561\,
            I => \N__5558\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__5558\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__5555\,
            I => \U712_CHIP_RAM.N_376_cascade_\
        );

    \I__859\ : CascadeMux
    port map (
            O => \N__5552\,
            I => \U712_CHIP_RAM.N_45_i_cascade_\
        );

    \I__858\ : InMux
    port map (
            O => \N__5549\,
            I => \N__5546\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__5546\,
            I => \U712_CHIP_RAM.N_324_2\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__5543\,
            I => \U712_CHIP_RAM.N_324_2_cascade_\
        );

    \I__855\ : CascadeMux
    port map (
            O => \N__5540\,
            I => \N__5537\
        );

    \I__854\ : InMux
    port map (
            O => \N__5537\,
            I => \N__5532\
        );

    \I__853\ : InMux
    port map (
            O => \N__5536\,
            I => \N__5529\
        );

    \I__852\ : InMux
    port map (
            O => \N__5535\,
            I => \N__5526\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__5532\,
            I => \U712_CHIP_RAM.N_450\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__5529\,
            I => \U712_CHIP_RAM.N_450\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__5526\,
            I => \U712_CHIP_RAM.N_450\
        );

    \I__848\ : InMux
    port map (
            O => \N__5519\,
            I => \N__5515\
        );

    \I__847\ : InMux
    port map (
            O => \N__5518\,
            I => \N__5512\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__5515\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIVIFVCZ0Z_4\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__5512\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIVIFVCZ0Z_4\
        );

    \I__844\ : InMux
    port map (
            O => \N__5507\,
            I => \N__5504\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__5504\,
            I => \U712_CHIP_RAM.N_252\
        );

    \I__842\ : CascadeMux
    port map (
            O => \N__5501\,
            I => \U712_CHIP_RAM.N_252_cascade_\
        );

    \I__841\ : CascadeMux
    port map (
            O => \N__5498\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\
        );

    \I__840\ : InMux
    port map (
            O => \N__5495\,
            I => \N__5492\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__5492\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\
        );

    \I__838\ : InMux
    port map (
            O => \N__5489\,
            I => \N__5486\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__5486\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_1\
        );

    \I__836\ : CascadeMux
    port map (
            O => \N__5483\,
            I => \U712_CHIP_RAM.N_325_cascade_\
        );

    \I__835\ : InMux
    port map (
            O => \N__5480\,
            I => \N__5477\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__5477\,
            I => \N__5474\
        );

    \I__833\ : Span4Mux_v
    port map (
            O => \N__5474\,
            I => \N__5471\
        );

    \I__832\ : Odrv4
    port map (
            O => \N__5471\,
            I => \U712_CHIP_RAM.N_301\
        );

    \I__831\ : CascadeMux
    port map (
            O => \N__5468\,
            I => \U712_CHIP_RAM.N_392_cascade_\
        );

    \I__830\ : InMux
    port map (
            O => \N__5465\,
            I => \N__5462\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__5462\,
            I => \U712_CHIP_RAM.N_449\
        );

    \I__828\ : InMux
    port map (
            O => \N__5459\,
            I => \N__5456\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__5456\,
            I => \N__5453\
        );

    \I__826\ : Span4Mux_h
    port map (
            O => \N__5453\,
            I => \N__5450\
        );

    \I__825\ : Span4Mux_v
    port map (
            O => \N__5450\,
            I => \N__5447\
        );

    \I__824\ : Sp12to4
    port map (
            O => \N__5447\,
            I => \N__5444\
        );

    \I__823\ : Odrv12
    port map (
            O => \N__5444\,
            I => \A_c_8\
        );

    \I__822\ : InMux
    port map (
            O => \N__5441\,
            I => \N__5438\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5438\,
            I => \N__5435\
        );

    \I__820\ : Span4Mux_v
    port map (
            O => \N__5435\,
            I => \N__5432\
        );

    \I__819\ : Span4Mux_v
    port map (
            O => \N__5432\,
            I => \N__5429\
        );

    \I__818\ : Sp12to4
    port map (
            O => \N__5429\,
            I => \N__5426\
        );

    \I__817\ : Span12Mux_h
    port map (
            O => \N__5426\,
            I => \N__5423\
        );

    \I__816\ : Odrv12
    port map (
            O => \N__5423\,
            I => \A_c_15\
        );

    \I__815\ : CascadeMux
    port map (
            O => \N__5420\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\
        );

    \I__814\ : InMux
    port map (
            O => \N__5417\,
            I => \N__5414\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5414\,
            I => \N__5411\
        );

    \I__812\ : Span4Mux_v
    port map (
            O => \N__5411\,
            I => \N__5408\
        );

    \I__811\ : Sp12to4
    port map (
            O => \N__5408\,
            I => \N__5405\
        );

    \I__810\ : Span12Mux_h
    port map (
            O => \N__5405\,
            I => \N__5402\
        );

    \I__809\ : Odrv12
    port map (
            O => \N__5402\,
            I => \A_c_13\
        );

    \I__808\ : InMux
    port map (
            O => \N__5399\,
            I => \N__5396\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__5396\,
            I => \N__5393\
        );

    \I__806\ : Span12Mux_v
    port map (
            O => \N__5393\,
            I => \N__5390\
        );

    \I__805\ : Span12Mux_h
    port map (
            O => \N__5390\,
            I => \N__5387\
        );

    \I__804\ : Odrv12
    port map (
            O => \N__5387\,
            I => \A_c_6\
        );

    \I__803\ : InMux
    port map (
            O => \N__5384\,
            I => \N__5381\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__5381\,
            I => \N__5378\
        );

    \I__801\ : Span12Mux_v
    port map (
            O => \N__5378\,
            I => \N__5375\
        );

    \I__800\ : Span12Mux_h
    port map (
            O => \N__5375\,
            I => \N__5372\
        );

    \I__799\ : Odrv12
    port map (
            O => \N__5372\,
            I => \A_c_16\
        );

    \I__798\ : InMux
    port map (
            O => \N__5369\,
            I => \N__5366\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5366\,
            I => \N__5363\
        );

    \I__796\ : Span12Mux_v
    port map (
            O => \N__5363\,
            I => \N__5360\
        );

    \I__795\ : Span12Mux_h
    port map (
            O => \N__5360\,
            I => \N__5357\
        );

    \I__794\ : Odrv12
    port map (
            O => \N__5357\,
            I => \A_c_18\
        );

    \I__793\ : CascadeMux
    port map (
            O => \N__5354\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5_cascade_\
        );

    \I__792\ : InMux
    port map (
            O => \N__5351\,
            I => \N__5348\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__5348\,
            I => \N__5345\
        );

    \I__790\ : Odrv4
    port map (
            O => \N__5345\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\
        );

    \I__789\ : IoInMux
    port map (
            O => \N__5342\,
            I => \N__5339\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__5339\,
            I => \N__5336\
        );

    \I__787\ : IoSpan4Mux
    port map (
            O => \N__5336\,
            I => \N__5333\
        );

    \I__786\ : Sp12to4
    port map (
            O => \N__5333\,
            I => \N__5330\
        );

    \I__785\ : Span12Mux_s7_h
    port map (
            O => \N__5330\,
            I => \N__5327\
        );

    \I__784\ : Span12Mux_v
    port map (
            O => \N__5327\,
            I => \N__5324\
        );

    \I__783\ : Odrv12
    port map (
            O => \N__5324\,
            I => \CMA_c_5\
        );

    \I__782\ : InMux
    port map (
            O => \N__5321\,
            I => \N__5318\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__5318\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\
        );

    \I__780\ : IoInMux
    port map (
            O => \N__5315\,
            I => \N__5312\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5312\,
            I => \N__5309\
        );

    \I__778\ : Span4Mux_s1_v
    port map (
            O => \N__5309\,
            I => \N__5306\
        );

    \I__777\ : Span4Mux_v
    port map (
            O => \N__5306\,
            I => \N__5303\
        );

    \I__776\ : Span4Mux_v
    port map (
            O => \N__5303\,
            I => \N__5300\
        );

    \I__775\ : Span4Mux_v
    port map (
            O => \N__5300\,
            I => \N__5297\
        );

    \I__774\ : Odrv4
    port map (
            O => \N__5297\,
            I => \CMA_c_1\
        );

    \I__773\ : InMux
    port map (
            O => \N__5294\,
            I => \N__5291\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__5291\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i\
        );

    \I__771\ : InMux
    port map (
            O => \N__5288\,
            I => \N__5285\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__5285\,
            I => \N__5282\
        );

    \I__769\ : Span4Mux_v
    port map (
            O => \N__5282\,
            I => \N__5279\
        );

    \I__768\ : Sp12to4
    port map (
            O => \N__5279\,
            I => \N__5276\
        );

    \I__767\ : Span12Mux_h
    port map (
            O => \N__5276\,
            I => \N__5273\
        );

    \I__766\ : Odrv12
    port map (
            O => \N__5273\,
            I => \A_c_11\
        );

    \I__765\ : InMux
    port map (
            O => \N__5270\,
            I => \N__5267\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5267\,
            I => \N__5264\
        );

    \I__763\ : Span12Mux_v
    port map (
            O => \N__5264\,
            I => \N__5261\
        );

    \I__762\ : Span12Mux_h
    port map (
            O => \N__5261\,
            I => \N__5258\
        );

    \I__761\ : Odrv12
    port map (
            O => \N__5258\,
            I => \A_c_4\
        );

    \I__760\ : InMux
    port map (
            O => \N__5255\,
            I => \N__5250\
        );

    \I__759\ : InMux
    port map (
            O => \N__5254\,
            I => \N__5247\
        );

    \I__758\ : InMux
    port map (
            O => \N__5253\,
            I => \N__5244\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__5250\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_7\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__5247\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_7\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__5244\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_7\
        );

    \I__754\ : CascadeMux
    port map (
            O => \N__5237\,
            I => \N__5234\
        );

    \I__753\ : InMux
    port map (
            O => \N__5234\,
            I => \N__5228\
        );

    \I__752\ : InMux
    port map (
            O => \N__5233\,
            I => \N__5221\
        );

    \I__751\ : InMux
    port map (
            O => \N__5232\,
            I => \N__5221\
        );

    \I__750\ : InMux
    port map (
            O => \N__5231\,
            I => \N__5221\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__5228\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_3\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__5221\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_3\
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__5216\,
            I => \U712_REG_SM.un18_0_i_0_0_1_cascade_\
        );

    \I__746\ : CascadeMux
    port map (
            O => \N__5213\,
            I => \N__5209\
        );

    \I__745\ : CascadeMux
    port map (
            O => \N__5212\,
            I => \N__5203\
        );

    \I__744\ : InMux
    port map (
            O => \N__5209\,
            I => \N__5198\
        );

    \I__743\ : InMux
    port map (
            O => \N__5208\,
            I => \N__5195\
        );

    \I__742\ : InMux
    port map (
            O => \N__5207\,
            I => \N__5188\
        );

    \I__741\ : InMux
    port map (
            O => \N__5206\,
            I => \N__5188\
        );

    \I__740\ : InMux
    port map (
            O => \N__5203\,
            I => \N__5188\
        );

    \I__739\ : InMux
    port map (
            O => \N__5202\,
            I => \N__5185\
        );

    \I__738\ : InMux
    port map (
            O => \N__5201\,
            I => \N__5182\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__5198\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_8\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__5195\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_8\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__5188\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_8\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__5185\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_8\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__5182\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_8\
        );

    \I__732\ : InMux
    port map (
            O => \N__5171\,
            I => \N__5167\
        );

    \I__731\ : InMux
    port map (
            O => \N__5170\,
            I => \N__5162\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__5167\,
            I => \N__5159\
        );

    \I__729\ : InMux
    port map (
            O => \N__5166\,
            I => \N__5154\
        );

    \I__728\ : InMux
    port map (
            O => \N__5165\,
            I => \N__5154\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__5162\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_4\
        );

    \I__726\ : Odrv4
    port map (
            O => \N__5159\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_4\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__5154\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_4\
        );

    \I__724\ : CascadeMux
    port map (
            O => \N__5147\,
            I => \U712_REG_SM.N_442_cascade_\
        );

    \I__723\ : CascadeMux
    port map (
            O => \N__5144\,
            I => \N__5141\
        );

    \I__722\ : InMux
    port map (
            O => \N__5141\,
            I => \N__5138\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__5138\,
            I => \N__5135\
        );

    \I__720\ : Odrv4
    port map (
            O => \N__5135\,
            I => \U712_REG_SM.REG_CPU_CYCLE_e_1\
        );

    \I__719\ : InMux
    port map (
            O => \N__5132\,
            I => \N__5129\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__5129\,
            I => \U712_REG_SM.N_84\
        );

    \I__717\ : CascadeMux
    port map (
            O => \N__5126\,
            I => \N__5120\
        );

    \I__716\ : CascadeMux
    port map (
            O => \N__5125\,
            I => \N__5115\
        );

    \I__715\ : CascadeMux
    port map (
            O => \N__5124\,
            I => \N__5109\
        );

    \I__714\ : InMux
    port map (
            O => \N__5123\,
            I => \N__5105\
        );

    \I__713\ : InMux
    port map (
            O => \N__5120\,
            I => \N__5102\
        );

    \I__712\ : InMux
    port map (
            O => \N__5119\,
            I => \N__5099\
        );

    \I__711\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5094\
        );

    \I__710\ : InMux
    port map (
            O => \N__5115\,
            I => \N__5094\
        );

    \I__709\ : InMux
    port map (
            O => \N__5114\,
            I => \N__5091\
        );

    \I__708\ : InMux
    port map (
            O => \N__5113\,
            I => \N__5084\
        );

    \I__707\ : InMux
    port map (
            O => \N__5112\,
            I => \N__5084\
        );

    \I__706\ : InMux
    port map (
            O => \N__5109\,
            I => \N__5084\
        );

    \I__705\ : InMux
    port map (
            O => \N__5108\,
            I => \N__5081\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__5105\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__5102\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5099\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__5094\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__5091\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__5084\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__5081\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__697\ : CascadeMux
    port map (
            O => \N__5066\,
            I => \N__5059\
        );

    \I__696\ : CascadeMux
    port map (
            O => \N__5065\,
            I => \N__5055\
        );

    \I__695\ : CascadeMux
    port map (
            O => \N__5064\,
            I => \N__5050\
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__5063\,
            I => \N__5047\
        );

    \I__693\ : InMux
    port map (
            O => \N__5062\,
            I => \N__5042\
        );

    \I__692\ : InMux
    port map (
            O => \N__5059\,
            I => \N__5039\
        );

    \I__691\ : InMux
    port map (
            O => \N__5058\,
            I => \N__5036\
        );

    \I__690\ : InMux
    port map (
            O => \N__5055\,
            I => \N__5031\
        );

    \I__689\ : InMux
    port map (
            O => \N__5054\,
            I => \N__5031\
        );

    \I__688\ : InMux
    port map (
            O => \N__5053\,
            I => \N__5028\
        );

    \I__687\ : InMux
    port map (
            O => \N__5050\,
            I => \N__5025\
        );

    \I__686\ : InMux
    port map (
            O => \N__5047\,
            I => \N__5020\
        );

    \I__685\ : InMux
    port map (
            O => \N__5046\,
            I => \N__5020\
        );

    \I__684\ : InMux
    port map (
            O => \N__5045\,
            I => \N__5017\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__5042\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__5039\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__5036\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__5031\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__5028\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__5025\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__5020\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__5017\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__675\ : InMux
    port map (
            O => \N__5000\,
            I => \N__4995\
        );

    \I__674\ : InMux
    port map (
            O => \N__4999\,
            I => \N__4992\
        );

    \I__673\ : InMux
    port map (
            O => \N__4998\,
            I => \N__4989\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__4995\,
            I => \U712_REG_SM.N_447\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__4992\,
            I => \U712_REG_SM.N_447\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__4989\,
            I => \U712_REG_SM.N_447\
        );

    \I__669\ : InMux
    port map (
            O => \N__4982\,
            I => \N__4976\
        );

    \I__668\ : InMux
    port map (
            O => \N__4981\,
            I => \N__4973\
        );

    \I__667\ : InMux
    port map (
            O => \N__4980\,
            I => \N__4968\
        );

    \I__666\ : InMux
    port map (
            O => \N__4979\,
            I => \N__4968\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__4976\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_6\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__4973\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_6\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__4968\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_6\
        );

    \I__662\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4958\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__4958\,
            I => \U712_REG_SM.N_288\
        );

    \I__660\ : InMux
    port map (
            O => \N__4955\,
            I => \N__4951\
        );

    \I__659\ : InMux
    port map (
            O => \N__4954\,
            I => \N__4948\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__4951\,
            I => \LATCH_REG\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__4948\,
            I => \LATCH_REG\
        );

    \I__656\ : IoInMux
    port map (
            O => \N__4943\,
            I => \N__4940\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__4940\,
            I => \N__4937\
        );

    \I__654\ : Span4Mux_s3_v
    port map (
            O => \N__4937\,
            I => \N__4934\
        );

    \I__653\ : Span4Mux_h
    port map (
            O => \N__4934\,
            I => \N__4931\
        );

    \I__652\ : Span4Mux_v
    port map (
            O => \N__4931\,
            I => \N__4928\
        );

    \I__651\ : Span4Mux_v
    port map (
            O => \N__4928\,
            I => \N__4925\
        );

    \I__650\ : Odrv4
    port map (
            O => \N__4925\,
            I => \LATCH_CLK_0_i\
        );

    \I__649\ : CascadeMux
    port map (
            O => \N__4922\,
            I => \U712_CHIP_RAM.N_452_cascade_\
        );

    \I__648\ : CascadeMux
    port map (
            O => \N__4919\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_cascade_\
        );

    \I__647\ : CEMux
    port map (
            O => \N__4916\,
            I => \N__4913\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__4913\,
            I => \N__4910\
        );

    \I__645\ : Odrv12
    port map (
            O => \N__4910\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0\
        );

    \I__644\ : IoInMux
    port map (
            O => \N__4907\,
            I => \N__4904\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__4904\,
            I => \N__4901\
        );

    \I__642\ : IoSpan4Mux
    port map (
            O => \N__4901\,
            I => \N__4898\
        );

    \I__641\ : IoSpan4Mux
    port map (
            O => \N__4898\,
            I => \N__4895\
        );

    \I__640\ : Span4Mux_s1_v
    port map (
            O => \N__4895\,
            I => \N__4892\
        );

    \I__639\ : Sp12to4
    port map (
            O => \N__4892\,
            I => \N__4889\
        );

    \I__638\ : Span12Mux_v
    port map (
            O => \N__4889\,
            I => \N__4883\
        );

    \I__637\ : InMux
    port map (
            O => \N__4888\,
            I => \N__4880\
        );

    \I__636\ : InMux
    port map (
            O => \N__4887\,
            I => \N__4877\
        );

    \I__635\ : InMux
    port map (
            O => \N__4886\,
            I => \N__4874\
        );

    \I__634\ : Odrv12
    port map (
            O => \N__4883\,
            I => \LDSn_c\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__4880\,
            I => \LDSn_c\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__4877\,
            I => \LDSn_c\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__4874\,
            I => \LDSn_c\
        );

    \I__630\ : InMux
    port map (
            O => \N__4865\,
            I => \N__4856\
        );

    \I__629\ : InMux
    port map (
            O => \N__4864\,
            I => \N__4856\
        );

    \I__628\ : InMux
    port map (
            O => \N__4863\,
            I => \N__4853\
        );

    \I__627\ : InMux
    port map (
            O => \N__4862\,
            I => \N__4850\
        );

    \I__626\ : InMux
    port map (
            O => \N__4861\,
            I => \N__4847\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__4856\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__4853\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__4850\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__4847\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__621\ : InMux
    port map (
            O => \N__4838\,
            I => \N__4835\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__4835\,
            I => \U712_REG_SM.N_309\
        );

    \I__619\ : InMux
    port map (
            O => \N__4832\,
            I => \N__4829\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__4829\,
            I => \U712_REG_SM.STATE_COUNTER_srsts_i_i_i_a3_2_0\
        );

    \I__617\ : CascadeMux
    port map (
            O => \N__4826\,
            I => \N__4822\
        );

    \I__616\ : InMux
    port map (
            O => \N__4825\,
            I => \N__4817\
        );

    \I__615\ : InMux
    port map (
            O => \N__4822\,
            I => \N__4817\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__4817\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_5\
        );

    \I__613\ : SRMux
    port map (
            O => \N__4814\,
            I => \N__4811\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__4811\,
            I => \N__4808\
        );

    \I__611\ : Odrv4
    port map (
            O => \N__4808\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__610\ : InMux
    port map (
            O => \N__4805\,
            I => \N__4802\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__4802\,
            I => \N__4799\
        );

    \I__608\ : Span4Mux_v
    port map (
            O => \N__4799\,
            I => \N__4796\
        );

    \I__607\ : Span4Mux_h
    port map (
            O => \N__4796\,
            I => \N__4793\
        );

    \I__606\ : Sp12to4
    port map (
            O => \N__4793\,
            I => \N__4790\
        );

    \I__605\ : Span12Mux_v
    port map (
            O => \N__4790\,
            I => \N__4787\
        );

    \I__604\ : Odrv12
    port map (
            O => \N__4787\,
            I => \A_c_14\
        );

    \I__603\ : InMux
    port map (
            O => \N__4784\,
            I => \N__4781\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__4781\,
            I => \N__4778\
        );

    \I__601\ : Span4Mux_v
    port map (
            O => \N__4778\,
            I => \N__4775\
        );

    \I__600\ : Sp12to4
    port map (
            O => \N__4775\,
            I => \N__4772\
        );

    \I__599\ : Odrv12
    port map (
            O => \N__4772\,
            I => \A_c_7\
        );

    \I__598\ : CascadeMux
    port map (
            O => \N__4769\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5_cascade_\
        );

    \I__597\ : IoInMux
    port map (
            O => \N__4766\,
            I => \N__4763\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__4763\,
            I => \N__4760\
        );

    \I__595\ : Span12Mux_s1_h
    port map (
            O => \N__4760\,
            I => \N__4757\
        );

    \I__594\ : Odrv12
    port map (
            O => \N__4757\,
            I => \DBRn_c_i_0\
        );

    \I__593\ : InMux
    port map (
            O => \N__4754\,
            I => \N__4751\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__4751\,
            I => \N__4748\
        );

    \I__591\ : Span4Mux_h
    port map (
            O => \N__4748\,
            I => \N__4745\
        );

    \I__590\ : Span4Mux_v
    port map (
            O => \N__4745\,
            I => \N__4742\
        );

    \I__589\ : Sp12to4
    port map (
            O => \N__4742\,
            I => \N__4739\
        );

    \I__588\ : Odrv12
    port map (
            O => \N__4739\,
            I => \A_c_20\
        );

    \I__587\ : CascadeMux
    port map (
            O => \N__4736\,
            I => \U712_CHIP_RAM.N_361_cascade_\
        );

    \I__586\ : IoInMux
    port map (
            O => \N__4733\,
            I => \N__4730\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__4730\,
            I => \N__4727\
        );

    \I__584\ : Span4Mux_s3_v
    port map (
            O => \N__4727\,
            I => \N__4724\
        );

    \I__583\ : Span4Mux_h
    port map (
            O => \N__4724\,
            I => \N__4721\
        );

    \I__582\ : Sp12to4
    port map (
            O => \N__4721\,
            I => \N__4718\
        );

    \I__581\ : Span12Mux_v
    port map (
            O => \N__4718\,
            I => \N__4715\
        );

    \I__580\ : Odrv12
    port map (
            O => \N__4715\,
            I => \BANK0_c\
        );

    \I__579\ : InMux
    port map (
            O => \N__4712\,
            I => \N__4709\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__4709\,
            I => \U712_CHIP_RAM.N_452\
        );

    \I__577\ : InMux
    port map (
            O => \N__4706\,
            I => \N__4703\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__4703\,
            I => \N__4700\
        );

    \I__575\ : Odrv4
    port map (
            O => \N__4700\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__574\ : InMux
    port map (
            O => \N__4697\,
            I => \N__4693\
        );

    \I__573\ : IoInMux
    port map (
            O => \N__4696\,
            I => \N__4690\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__4693\,
            I => \N__4687\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__4690\,
            I => \N__4684\
        );

    \I__570\ : Span4Mux_v
    port map (
            O => \N__4687\,
            I => \N__4681\
        );

    \I__569\ : IoSpan4Mux
    port map (
            O => \N__4684\,
            I => \N__4678\
        );

    \I__568\ : Sp12to4
    port map (
            O => \N__4681\,
            I => \N__4675\
        );

    \I__567\ : IoSpan4Mux
    port map (
            O => \N__4678\,
            I => \N__4672\
        );

    \I__566\ : Span12Mux_h
    port map (
            O => \N__4675\,
            I => \N__4669\
        );

    \I__565\ : IoSpan4Mux
    port map (
            O => \N__4672\,
            I => \N__4666\
        );

    \I__564\ : Odrv12
    port map (
            O => \N__4669\,
            I => \C1_c\
        );

    \I__563\ : Odrv4
    port map (
            O => \N__4666\,
            I => \C1_c\
        );

    \I__562\ : InMux
    port map (
            O => \N__4661\,
            I => \N__4658\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__4658\,
            I => \N__4655\
        );

    \I__560\ : Odrv4
    port map (
            O => \N__4655\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__559\ : InMux
    port map (
            O => \N__4652\,
            I => \N__4649\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__4649\,
            I => \N__4646\
        );

    \I__557\ : Sp12to4
    port map (
            O => \N__4646\,
            I => \N__4643\
        );

    \I__556\ : Span12Mux_v
    port map (
            O => \N__4643\,
            I => \N__4640\
        );

    \I__555\ : Span12Mux_h
    port map (
            O => \N__4640\,
            I => \N__4637\
        );

    \I__554\ : Odrv12
    port map (
            O => \N__4637\,
            I => \A_c_3\
        );

    \I__553\ : CascadeMux
    port map (
            O => \N__4634\,
            I => \U712_CHIP_RAM.N_241_cascade_\
        );

    \I__552\ : InMux
    port map (
            O => \N__4631\,
            I => \N__4628\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__4628\,
            I => \U712_BYTE_ENABLE.N_276\
        );

    \I__550\ : CascadeMux
    port map (
            O => \N__4625\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0Z0Z_0_cascade_\
        );

    \I__549\ : IoInMux
    port map (
            O => \N__4622\,
            I => \N__4619\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__4619\,
            I => \N__4616\
        );

    \I__547\ : Span4Mux_s2_v
    port map (
            O => \N__4616\,
            I => \N__4613\
        );

    \I__546\ : Span4Mux_v
    port map (
            O => \N__4613\,
            I => \N__4610\
        );

    \I__545\ : Span4Mux_v
    port map (
            O => \N__4610\,
            I => \N__4607\
        );

    \I__544\ : Span4Mux_v
    port map (
            O => \N__4607\,
            I => \N__4604\
        );

    \I__543\ : Odrv4
    port map (
            O => \N__4604\,
            I => \N_47_i\
        );

    \I__542\ : InMux
    port map (
            O => \N__4601\,
            I => \N__4597\
        );

    \I__541\ : InMux
    port map (
            O => \N__4600\,
            I => \N__4594\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__4597\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__4594\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__538\ : InMux
    port map (
            O => \N__4589\,
            I => \N__4585\
        );

    \I__537\ : InMux
    port map (
            O => \N__4588\,
            I => \N__4582\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4585\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4582\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__534\ : CascadeMux
    port map (
            O => \N__4577\,
            I => \N__4573\
        );

    \I__533\ : InMux
    port map (
            O => \N__4576\,
            I => \N__4570\
        );

    \I__532\ : InMux
    port map (
            O => \N__4573\,
            I => \N__4567\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__4570\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__4567\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__529\ : InMux
    port map (
            O => \N__4562\,
            I => \N__4558\
        );

    \I__528\ : InMux
    port map (
            O => \N__4561\,
            I => \N__4555\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__4558\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__4555\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__525\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4547\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__4547\,
            I => \U712_REG_SM.N_266\
        );

    \I__523\ : CascadeMux
    port map (
            O => \N__4544\,
            I => \U712_REG_SM.STATE_COUNTER_srsts_i_i_i_a3_3_0_cascade_\
        );

    \I__522\ : InMux
    port map (
            O => \N__4541\,
            I => \N__4538\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4538\,
            I => \N__4535\
        );

    \I__520\ : Span4Mux_v
    port map (
            O => \N__4535\,
            I => \N__4532\
        );

    \I__519\ : Sp12to4
    port map (
            O => \N__4532\,
            I => \N__4529\
        );

    \I__518\ : Span12Mux_h
    port map (
            O => \N__4529\,
            I => \N__4526\
        );

    \I__517\ : Span12Mux_v
    port map (
            O => \N__4526\,
            I => \N__4523\
        );

    \I__516\ : Odrv12
    port map (
            O => \N__4523\,
            I => \REGSPACEn_c\
        );

    \I__515\ : InMux
    port map (
            O => \N__4520\,
            I => \N__4516\
        );

    \I__514\ : InMux
    port map (
            O => \N__4519\,
            I => \N__4513\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4516\,
            I => \U712_REG_SM.CYCLE_RUNZ0\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__4513\,
            I => \U712_REG_SM.CYCLE_RUNZ0\
        );

    \I__511\ : InMux
    port map (
            O => \N__4508\,
            I => \N__4502\
        );

    \I__510\ : InMux
    port map (
            O => \N__4507\,
            I => \N__4497\
        );

    \I__509\ : InMux
    port map (
            O => \N__4506\,
            I => \N__4497\
        );

    \I__508\ : InMux
    port map (
            O => \N__4505\,
            I => \N__4494\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__4502\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__4497\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4494\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__504\ : InMux
    port map (
            O => \N__4487\,
            I => \N__4478\
        );

    \I__503\ : InMux
    port map (
            O => \N__4486\,
            I => \N__4475\
        );

    \I__502\ : InMux
    port map (
            O => \N__4485\,
            I => \N__4472\
        );

    \I__501\ : InMux
    port map (
            O => \N__4484\,
            I => \N__4469\
        );

    \I__500\ : InMux
    port map (
            O => \N__4483\,
            I => \N__4462\
        );

    \I__499\ : InMux
    port map (
            O => \N__4482\,
            I => \N__4462\
        );

    \I__498\ : InMux
    port map (
            O => \N__4481\,
            I => \N__4462\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__4478\,
            I => \N__4457\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__4475\,
            I => \N__4457\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__4472\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_9\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4469\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_9\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__4462\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_9\
        );

    \I__492\ : Odrv4
    port map (
            O => \N__4457\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_9\
        );

    \I__491\ : InMux
    port map (
            O => \N__4448\,
            I => \N__4443\
        );

    \I__490\ : InMux
    port map (
            O => \N__4447\,
            I => \N__4438\
        );

    \I__489\ : InMux
    port map (
            O => \N__4446\,
            I => \N__4438\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__4443\,
            I => \N__4433\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__4438\,
            I => \N__4433\
        );

    \I__486\ : Odrv4
    port map (
            O => \N__4433\,
            I => \U712_REG_SM.N_71_i\
        );

    \I__485\ : InMux
    port map (
            O => \N__4430\,
            I => \N__4427\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4427\,
            I => \N__4423\
        );

    \I__483\ : InMux
    port map (
            O => \N__4426\,
            I => \N__4420\
        );

    \I__482\ : Odrv12
    port map (
            O => \N__4423\,
            I => \REG_CPU_CYCLE\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__4420\,
            I => \REG_CPU_CYCLE\
        );

    \I__480\ : IoInMux
    port map (
            O => \N__4415\,
            I => \N__4412\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4412\,
            I => \N__4409\
        );

    \I__478\ : IoSpan4Mux
    port map (
            O => \N__4409\,
            I => \N__4406\
        );

    \I__477\ : Span4Mux_s0_h
    port map (
            O => \N__4406\,
            I => \N__4403\
        );

    \I__476\ : Span4Mux_h
    port map (
            O => \N__4403\,
            I => \N__4399\
        );

    \I__475\ : InMux
    port map (
            O => \N__4402\,
            I => \N__4396\
        );

    \I__474\ : Sp12to4
    port map (
            O => \N__4399\,
            I => \N__4393\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__4396\,
            I => \N__4390\
        );

    \I__472\ : Span12Mux_v
    port map (
            O => \N__4393\,
            I => \N__4387\
        );

    \I__471\ : Span4Mux_v
    port map (
            O => \N__4390\,
            I => \N__4384\
        );

    \I__470\ : Span12Mux_h
    port map (
            O => \N__4387\,
            I => \N__4381\
        );

    \I__469\ : Sp12to4
    port map (
            O => \N__4384\,
            I => \N__4378\
        );

    \I__468\ : Span12Mux_h
    port map (
            O => \N__4381\,
            I => \N__4375\
        );

    \I__467\ : Span12Mux_h
    port map (
            O => \N__4378\,
            I => \N__4372\
        );

    \I__466\ : Odrv12
    port map (
            O => \N__4375\,
            I => \C3_c\
        );

    \I__465\ : Odrv12
    port map (
            O => \N__4372\,
            I => \C3_c\
        );

    \I__464\ : InMux
    port map (
            O => \N__4367\,
            I => \N__4364\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__4364\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0\
        );

    \I__462\ : IoInMux
    port map (
            O => \N__4361\,
            I => \N__4358\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__4358\,
            I => \N__4355\
        );

    \I__460\ : Span4Mux_s3_h
    port map (
            O => \N__4355\,
            I => \N__4352\
        );

    \I__459\ : Span4Mux_h
    port map (
            O => \N__4352\,
            I => \N__4349\
        );

    \I__458\ : Span4Mux_h
    port map (
            O => \N__4349\,
            I => \N__4346\
        );

    \I__457\ : Sp12to4
    port map (
            O => \N__4346\,
            I => \N__4342\
        );

    \I__456\ : InMux
    port map (
            O => \N__4345\,
            I => \N__4339\
        );

    \I__455\ : Odrv12
    port map (
            O => \N__4342\,
            I => \TACK_OUTn\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__4339\,
            I => \TACK_OUTn\
        );

    \I__453\ : CascadeMux
    port map (
            O => \N__4334\,
            I => \U712_REG_SM.N_295_cascade_\
        );

    \I__452\ : InMux
    port map (
            O => \N__4331\,
            I => \N__4328\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__4328\,
            I => \U712_REG_SM.LDSn_6_iv_i_0_0\
        );

    \I__450\ : InMux
    port map (
            O => \N__4325\,
            I => \N__4318\
        );

    \I__449\ : InMux
    port map (
            O => \N__4324\,
            I => \N__4318\
        );

    \I__448\ : InMux
    port map (
            O => \N__4323\,
            I => \N__4315\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__4318\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__4315\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__445\ : InMux
    port map (
            O => \N__4310\,
            I => \N__4307\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__4307\,
            I => \U712_REG_SM.N_332\
        );

    \I__443\ : CascadeMux
    port map (
            O => \N__4304\,
            I => \N__4301\
        );

    \I__442\ : InMux
    port map (
            O => \N__4301\,
            I => \N__4298\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__4298\,
            I => \U712_REG_SM.UDSn_6_iv_i_0_0\
        );

    \I__440\ : InMux
    port map (
            O => \N__4295\,
            I => \N__4291\
        );

    \I__439\ : InMux
    port map (
            O => \N__4294\,
            I => \N__4288\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__4291\,
            I => \U712_REG_SM.STATE_COUNTER_RNI7KTS1Z0Z_9\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__4288\,
            I => \U712_REG_SM.STATE_COUNTER_RNI7KTS1Z0Z_9\
        );

    \I__436\ : IoInMux
    port map (
            O => \N__4283\,
            I => \N__4280\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__4280\,
            I => \N__4277\
        );

    \I__434\ : Span4Mux_s2_v
    port map (
            O => \N__4277\,
            I => \N__4274\
        );

    \I__433\ : Span4Mux_h
    port map (
            O => \N__4274\,
            I => \N__4271\
        );

    \I__432\ : Sp12to4
    port map (
            O => \N__4271\,
            I => \N__4268\
        );

    \I__431\ : Span12Mux_h
    port map (
            O => \N__4268\,
            I => \N__4263\
        );

    \I__430\ : InMux
    port map (
            O => \N__4267\,
            I => \N__4260\
        );

    \I__429\ : InMux
    port map (
            O => \N__4266\,
            I => \N__4257\
        );

    \I__428\ : Odrv12
    port map (
            O => \N__4263\,
            I => \UDSn_c\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__4260\,
            I => \UDSn_c\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__4257\,
            I => \UDSn_c\
        );

    \I__425\ : InMux
    port map (
            O => \N__4250\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__424\ : InMux
    port map (
            O => \N__4247\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__423\ : InMux
    port map (
            O => \N__4244\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__422\ : InMux
    port map (
            O => \N__4241\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__421\ : InMux
    port map (
            O => \N__4238\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__420\ : InMux
    port map (
            O => \N__4235\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__419\ : ClkMux
    port map (
            O => \N__4232\,
            I => \N__4205\
        );

    \I__418\ : ClkMux
    port map (
            O => \N__4231\,
            I => \N__4205\
        );

    \I__417\ : ClkMux
    port map (
            O => \N__4230\,
            I => \N__4205\
        );

    \I__416\ : ClkMux
    port map (
            O => \N__4229\,
            I => \N__4205\
        );

    \I__415\ : ClkMux
    port map (
            O => \N__4228\,
            I => \N__4205\
        );

    \I__414\ : ClkMux
    port map (
            O => \N__4227\,
            I => \N__4205\
        );

    \I__413\ : ClkMux
    port map (
            O => \N__4226\,
            I => \N__4205\
        );

    \I__412\ : ClkMux
    port map (
            O => \N__4225\,
            I => \N__4205\
        );

    \I__411\ : ClkMux
    port map (
            O => \N__4224\,
            I => \N__4205\
        );

    \I__410\ : GlobalMux
    port map (
            O => \N__4205\,
            I => \N__4202\
        );

    \I__409\ : gio2CtrlBuf
    port map (
            O => \N__4202\,
            I => \C1_c_g\
        );

    \I__408\ : CascadeMux
    port map (
            O => \N__4199\,
            I => \U712_REG_SM.N_330_cascade_\
        );

    \I__407\ : IoInMux
    port map (
            O => \N__4196\,
            I => \N__4193\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__4193\,
            I => \N__4190\
        );

    \I__405\ : Span4Mux_s3_v
    port map (
            O => \N__4190\,
            I => \N__4187\
        );

    \I__404\ : Span4Mux_h
    port map (
            O => \N__4187\,
            I => \N__4184\
        );

    \I__403\ : Span4Mux_h
    port map (
            O => \N__4184\,
            I => \N__4181\
        );

    \I__402\ : Sp12to4
    port map (
            O => \N__4181\,
            I => \N__4178\
        );

    \I__401\ : Span12Mux_s11_v
    port map (
            O => \N__4178\,
            I => \N__4174\
        );

    \I__400\ : InMux
    port map (
            O => \N__4177\,
            I => \N__4171\
        );

    \I__399\ : Odrv12
    port map (
            O => \N__4174\,
            I => \ASn_c\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__4171\,
            I => \ASn_c\
        );

    \I__397\ : IoInMux
    port map (
            O => \N__4166\,
            I => \N__4163\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__4163\,
            I => \N__4160\
        );

    \I__395\ : IoSpan4Mux
    port map (
            O => \N__4160\,
            I => \N__4157\
        );

    \I__394\ : Span4Mux_s2_v
    port map (
            O => \N__4157\,
            I => \N__4154\
        );

    \I__393\ : Span4Mux_v
    port map (
            O => \N__4154\,
            I => \N__4151\
        );

    \I__392\ : Span4Mux_v
    port map (
            O => \N__4151\,
            I => \N__4147\
        );

    \I__391\ : InMux
    port map (
            O => \N__4150\,
            I => \N__4144\
        );

    \I__390\ : Odrv4
    port map (
            O => \N__4147\,
            I => \REGENn_c\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__4144\,
            I => \REGENn_c\
        );

    \I__388\ : IoInMux
    port map (
            O => \N__4139\,
            I => \N__4136\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__4136\,
            I => \N__4133\
        );

    \I__386\ : Span12Mux_s7_v
    port map (
            O => \N__4133\,
            I => \N__4130\
        );

    \I__385\ : Odrv12
    port map (
            O => \N__4130\,
            I => \VBENn_c\
        );

    \I__384\ : InMux
    port map (
            O => \N__4127\,
            I => \N__4124\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__4124\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__382\ : InMux
    port map (
            O => \N__4121\,
            I => \bfn_8_10_0_\
        );

    \I__381\ : InMux
    port map (
            O => \N__4118\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__380\ : IoInMux
    port map (
            O => \N__4115\,
            I => \N__4112\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__4112\,
            I => \N__4109\
        );

    \I__378\ : Span4Mux_s2_v
    port map (
            O => \N__4109\,
            I => \N__4106\
        );

    \I__377\ : Span4Mux_v
    port map (
            O => \N__4106\,
            I => \N__4103\
        );

    \I__376\ : Odrv4
    port map (
            O => \N__4103\,
            I => \CLK80_PLL_i_i\
        );

    \I__375\ : IoInMux
    port map (
            O => \N__4100\,
            I => \N__4097\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__4097\,
            I => \N__4094\
        );

    \I__373\ : IoSpan4Mux
    port map (
            O => \N__4094\,
            I => \N__4091\
        );

    \I__372\ : IoSpan4Mux
    port map (
            O => \N__4091\,
            I => \N__4088\
        );

    \I__371\ : Span4Mux_s2_h
    port map (
            O => \N__4088\,
            I => \N__4085\
        );

    \I__370\ : Span4Mux_h
    port map (
            O => \N__4085\,
            I => \N__4082\
        );

    \I__369\ : Odrv4
    port map (
            O => \N__4082\,
            I => \N_882_i\
        );

    \I__368\ : CascadeMux
    port map (
            O => \N__4079\,
            I => \U712_REG_SM.N_71_i_cascade_\
        );

    \I__367\ : InMux
    port map (
            O => \N__4076\,
            I => \N__4073\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__4073\,
            I => \N__4070\
        );

    \I__365\ : Span4Mux_v
    port map (
            O => \N__4070\,
            I => \N__4067\
        );

    \I__364\ : Odrv4
    port map (
            O => \N__4067\,
            I => \TACK_EN_i_ess\
        );

    \I__363\ : CascadeMux
    port map (
            O => \N__4064\,
            I => \U712_REG_SM.N_265_cascade_\
        );

    \I__362\ : IoInMux
    port map (
            O => \N__4061\,
            I => \N__4058\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__4058\,
            I => \N__4055\
        );

    \I__360\ : IoSpan4Mux
    port map (
            O => \N__4055\,
            I => \N__4052\
        );

    \I__359\ : Span4Mux_s2_v
    port map (
            O => \N__4052\,
            I => \N__4049\
        );

    \I__358\ : Sp12to4
    port map (
            O => \N__4049\,
            I => \N__4046\
        );

    \I__357\ : Span12Mux_v
    port map (
            O => \N__4046\,
            I => \N__4043\
        );

    \I__356\ : Odrv12
    port map (
            O => \N__4043\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__4229\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            I => \N__4230\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__4231\
        );

    \INVU712_CHIP_RAM.DMA_A20C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A20C_net\,
            I => \N__4225\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            I => \N__4227\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            I => \N__4224\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            I => \N__4226\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            I => \N__4228\
        );

    \INVU712_REG_SM.STATE_COUNTER_2C\ : INV
    port map (
            O => \INVU712_REG_SM.STATE_COUNTER_2C_net\,
            I => \N__8862\
        );

    \INVU712_REG_SM.STATE_COUNTER_5C\ : INV
    port map (
            O => \INVU712_REG_SM.STATE_COUNTER_5C_net\,
            I => \N__8863\
        );

    \INVU712_REG_SM.C3_SYNC_0C\ : INV
    port map (
            O => \INVU712_REG_SM.C3_SYNC_0C_net\,
            I => \N__8870\
        );

    \INVU712_REG_SM.LATCH_REGC\ : INV
    port map (
            O => \INVU712_REG_SM.LATCH_REGC_net\,
            I => \N__8865\
        );

    \INVU712_REG_SM.UDSnC\ : INV
    port map (
            O => \INVU712_REG_SM.UDSnC_net\,
            I => \N__8864\
        );

    \INVU712_REG_SM.LDSnC\ : INV
    port map (
            O => \INVU712_REG_SM.LDSnC_net\,
            I => \N__8861\
        );

    \INVU712_REG_SM.REGENnC\ : INV
    port map (
            O => \INVU712_REG_SM.REGENnC_net\,
            I => \N__8871\
        );

    \INVU712_REG_SM.STATE_COUNTER_9C\ : INV
    port map (
            O => \INVU712_REG_SM.STATE_COUNTER_9C_net\,
            I => \N__8869\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_10_0_\
        );

    \CLK40_PLL_derived_clock_RNIIOT\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8335\,
            GLOBALBUFFEROUTPUT => \CLK40_PLL_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8381\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4696\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4766\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4415\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9926\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_obuft_RNO_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4076\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_882_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8284\,
            in1 => \N__8169\,
            in2 => \N__8212\,
            in3 => \N__4323\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNIQANC1_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__4505\,
            in1 => \N__5114\,
            in2 => \N__5064\,
            in3 => \N__4861\,
            lcout => \U712_REG_SM.N_71_i\,
            ltout => \U712_REG_SM.N_71_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNTER_RNI7KTS1_9_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4487\,
            in2 => \N__4079\,
            in3 => \N__6026\,
            lcout => \U712_REG_SM.STATE_COUNTER_RNI7KTS1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001111111111111"
        )
    port map (
            in0 => \N__8216\,
            in1 => \N__8256\,
            in2 => \N__8362\,
            in3 => \N__8498\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9922\,
            ce => \N__7370\,
            sr => \N__10819\
        );

    \U712_REG_SM.C1_SYNC_RNI6FIN_1_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5045\,
            in2 => \_gnd_net_\,
            in3 => \N__5108\,
            lcout => \U712_REG_SM.N_265\,
            ltout => \U712_REG_SM.N_265_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDSn_RNO_0_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__9261\,
            in1 => \N__4266\,
            in2 => \N__4064\,
            in3 => \N__6022\,
            lcout => \U712_REG_SM.N_332\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNTER_RNO_0_0_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__4506\,
            in1 => \N__5054\,
            in2 => \N__5125\,
            in3 => \N__4481\,
            lcout => \U712_REG_SM.N_266\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNTER_9_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5119\,
            in1 => \N__5208\,
            in2 => \_gnd_net_\,
            in3 => \N__5062\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_9C_net\,
            ce => 'H',
            sr => \N__10811\
        );

    \U712_REG_SM.UDSn_RNO_1_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111001100"
        )
    port map (
            in0 => \N__9260\,
            in1 => \N__4482\,
            in2 => \N__5758\,
            in3 => \N__4864\,
            lcout => \U712_REG_SM.UDSn_6_iv_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNTER_1_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4865\,
            in1 => \N__4507\,
            in2 => \N__5065\,
            in3 => \N__5118\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_9C_net\,
            ce => 'H',
            sr => \N__10811\
        );

    \U712_REG_SM.ASn_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__4447\,
            in1 => \N__4177\,
            in2 => \_gnd_net_\,
            in3 => \N__4483\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_9C_net\,
            ce => 'H',
            sr => \N__10811\
        );

    \U712_REG_SM.CYCLE_RUN_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__6049\,
            in1 => \N__4519\,
            in2 => \_gnd_net_\,
            in3 => \N__4446\,
            lcout => \U712_REG_SM.CYCLE_RUNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_9C_net\,
            ce => 'H',
            sr => \N__10811\
        );

    \U712_REG_SM.REGENn_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110011101110"
        )
    port map (
            in0 => \N__4150\,
            in1 => \N__4485\,
            in2 => \N__5213\,
            in3 => \N__6047\,
            lcout => \REGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REGENnC_net\,
            ce => 'H',
            sr => \N__10807\
        );

    \U712_BUFFERS.un1_VBENn_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4430\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9592\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_0_i_o3_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010110011"
        )
    port map (
            in0 => \N__9246\,
            in1 => \N__9180\,
            in2 => \N__9094\,
            in3 => \N__9021\,
            lcout => \U712_BYTE_ENABLE.N_276\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4127\,
            in2 => \_gnd_net_\,
            in3 => \N__4121\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__4232\,
            ce => 'H',
            sr => \N__4814\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4562\,
            in2 => \_gnd_net_\,
            in3 => \N__4118\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__4232\,
            ce => 'H',
            sr => \N__4814\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4589\,
            in2 => \_gnd_net_\,
            in3 => \N__4250\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__4232\,
            ce => 'H',
            sr => \N__4814\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4601\,
            in2 => \_gnd_net_\,
            in3 => \N__4247\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__4232\,
            ce => 'H',
            sr => \N__4814\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4576\,
            in2 => \_gnd_net_\,
            in3 => \N__4244\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__4232\,
            ce => 'H',
            sr => \N__4814\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6190\,
            in2 => \_gnd_net_\,
            in3 => \N__4241\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__4232\,
            ce => 'H',
            sr => \N__4814\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6205\,
            in2 => \_gnd_net_\,
            in3 => \N__4238\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__4232\,
            ce => 'H',
            sr => \N__4814\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6172\,
            in2 => \_gnd_net_\,
            in3 => \N__4235\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4232\,
            ce => 'H',
            sr => \N__4814\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__7586\,
            in1 => \N__8582\,
            in2 => \N__6599\,
            in3 => \N__7664\,
            lcout => \DMA_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9917\,
            ce => \N__6524\,
            sr => \N__10837\
        );

    \U712_REG_SM.LDSn_RNO_0_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__8997\,
            in1 => \N__9245\,
            in2 => \N__9167\,
            in3 => \N__4838\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_330_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101011001100"
        )
    port map (
            in0 => \N__4331\,
            in1 => \N__4888\,
            in2 => \N__4199\,
            in3 => \N__4295\,
            lcout => \LDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.LDSnC_net\,
            ce => 'H',
            sr => \N__10829\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__8170\,
            in1 => \N__4367\,
            in2 => \N__7394\,
            in3 => \N__8248\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9921\,
            ce => 'H',
            sr => \N__10820\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110110011101110"
        )
    port map (
            in0 => \N__4345\,
            in1 => \N__4324\,
            in2 => \N__8339\,
            in3 => \N__8171\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9921\,
            ce => 'H',
            sr => \N__10820\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4325\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9921\,
            ce => 'H',
            sr => \N__10820\
        );

    \U712_REG_SM.LDSn_RNO_3_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__5759\,
            in1 => \N__4486\,
            in2 => \_gnd_net_\,
            in3 => \N__4863\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_295_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_RNO_1_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__6067\,
            in1 => \N__4887\,
            in2 => \N__4334\,
            in3 => \N__6025\,
            lcout => \U712_REG_SM.LDSn_6_iv_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8288\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9921\,
            ce => 'H',
            sr => \N__10820\
        );

    \U712_REG_SM.UDSn_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110010101010"
        )
    port map (
            in0 => \N__4267\,
            in1 => \N__4310\,
            in2 => \N__4304\,
            in3 => \N__4294\,
            lcout => \UDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.UDSnC_net\,
            ce => 'H',
            sr => \N__10812\
        );

    \U712_REG_SM.C1_SYNC_1_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4661\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.UDSnC_net\,
            ce => 'H',
            sr => \N__10812\
        );

    \U712_REG_SM.C3_SYNC_1_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4706\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.UDSnC_net\,
            ce => 'H',
            sr => \N__10812\
        );

    \U712_REG_SM.STATE_COUNTER_RNO_1_0_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5253\,
            in1 => \N__4832\,
            in2 => \_gnd_net_\,
            in3 => \N__5202\,
            lcout => OPEN,
            ltout => \U712_REG_SM.STATE_COUNTER_srsts_i_i_i_a3_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNTER_0_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6048\,
            in1 => \N__4550\,
            in2 => \N__4544\,
            in3 => \N__6023\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.UDSnC_net\,
            ce => 'H',
            sr => \N__10812\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011100000101"
        )
    port map (
            in0 => \N__4541\,
            in1 => \N__4520\,
            in2 => \N__5653\,
            in3 => \N__4508\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.UDSnC_net\,
            ce => 'H',
            sr => \N__10812\
        );

    \U712_REG_SM.LATCH_REG_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110100000"
        )
    port map (
            in0 => \N__5892\,
            in1 => \N__4484\,
            in2 => \N__5237\,
            in3 => \N__4954\,
            lcout => \LATCH_REG\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.LATCH_REGC_net\,
            ce => 'H',
            sr => \N__10808\
        );

    \U712_REG_SM.REG_WRITE_CYCLE_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__5756\,
            in1 => \N__4448\,
            in2 => \_gnd_net_\,
            in3 => \N__5893\,
            lcout => \REG_WRITE_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.LATCH_REGC_net\,
            ce => 'H',
            sr => \N__10808\
        );

    \U712_REG_SM.REG_CPU_CYCLE_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000011100101"
        )
    port map (
            in0 => \N__5170\,
            in1 => \N__4426\,
            in2 => \N__5144\,
            in3 => \N__5206\,
            lcout => \REG_CPU_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.LATCH_REGC_net\,
            ce => 'H',
            sr => \N__10808\
        );

    \U712_REG_SM.REG_CYCLE_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100111010"
        )
    port map (
            in0 => \N__7992\,
            in1 => \N__5132\,
            in2 => \N__5212\,
            in3 => \N__5000\,
            lcout => \REG_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.LATCH_REGC_net\,
            ce => 'H',
            sr => \N__10808\
        );

    \U712_REG_SM.STATE_COUNTER_8_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__5255\,
            in1 => \N__5058\,
            in2 => \N__5126\,
            in3 => \N__5207\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.LATCH_REGC_net\,
            ce => 'H',
            sr => \N__10808\
        );

    \U712_REG_SM.STATE_COUNTER_7_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4982\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.LATCH_REGC_net\,
            ce => 'H',
            sr => \N__10808\
        );

    \U712_REG_SM.C3_SYNC_0_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4402\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C3_SYNC_0C_net\,
            ce => 'H',
            sr => \N__10801\
        );

    \U712_REG_SM.C1_SYNC_0_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4697\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C3_SYNC_0C_net\,
            ce => 'H',
            sr => \N__10801\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4652\,
            in1 => \N__9519\,
            in2 => \_gnd_net_\,
            in3 => \N__9326\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_241_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10024\,
            in2 => \N__4634\,
            in3 => \N__9727\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LMBE_0_a3_i_o3_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010001001111"
        )
    port map (
            in0 => \N__9273\,
            in1 => \N__9110\,
            in2 => \N__9185\,
            in3 => \N__9022\,
            lcout => \U712_BYTE_ENABLE.N_278\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__7330\,
            in1 => \N__6949\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0Z0Z_0\,
            ltout => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_47_i_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001110101111"
        )
    port map (
            in0 => \N__8111\,
            in1 => \N__4631\,
            in2 => \N__4625\,
            in3 => \N__9591\,
            lcout => \N_47_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100111"
        )
    port map (
            in0 => \N__10295\,
            in1 => \N__9665\,
            in2 => \N__10216\,
            in3 => \N__10248\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__4600\,
            in1 => \N__4588\,
            in2 => \N__4577\,
            in3 => \N__4561\,
            lcout => \U712_CHIP_RAM.REFRESH5lt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__10294\,
            in1 => \N__9664\,
            in2 => \N__10215\,
            in3 => \N__10247\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4805\,
            in1 => \N__4784\,
            in2 => \_gnd_net_\,
            in3 => \N__9709\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9710\,
            in1 => \N__9495\,
            in2 => \N__4769\,
            in3 => \N__10658\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011010101"
        )
    port map (
            in0 => \N__5489\,
            in1 => \N__5535\,
            in2 => \N__7093\,
            in3 => \N__8581\,
            lcout => \U712_CHIP_RAM.N_301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6147\,
            in1 => \N__8459\,
            in2 => \N__6662\,
            in3 => \N__7215\,
            lcout => \U712_CHIP_RAM.N_359\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10639\,
            in2 => \_gnd_net_\,
            in3 => \N__10873\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6655\,
            in1 => \N__4754\,
            in2 => \N__11192\,
            in3 => \N__4712\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_361_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__7232\,
            in1 => \N__6656\,
            in2 => \N__4736\,
            in3 => \N__10628\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9918\,
            ce => \N__5771\,
            sr => \N__10821\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIH3Q74_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5620\,
            in1 => \N__5583\,
            in2 => \N__6149\,
            in3 => \N__7214\,
            lcout => \U712_CHIP_RAM.N_452\,
            ltout => \U712_CHIP_RAM.N_452_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__6654\,
            in1 => \N__7727\,
            in2 => \N__4922\,
            in3 => \N__7882\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10872\,
            in1 => \_gnd_net_\,
            in2 => \N__4919\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5621\,
            in1 => \N__5587\,
            in2 => \N__7246\,
            in3 => \N__6148\,
            lcout => \CPU_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9920\,
            ce => \N__4916\,
            sr => \N__10813\
        );

    \U712_CHIP_RAM.LATCH_RAM_RNO_0_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__7754\,
            in1 => \N__6548\,
            in2 => \_gnd_net_\,
            in3 => \N__7784\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_RNO_2_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__4886\,
            in1 => \N__4862\,
            in2 => \_gnd_net_\,
            in3 => \N__6011\,
            lcout => \U712_REG_SM.N_309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNTER_RNO_2_0_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4979\,
            in1 => \N__5165\,
            in2 => \N__4826\,
            in3 => \N__5231\,
            lcout => \U712_REG_SM.STATE_COUNTER_srsts_i_i_i_a3_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNTER_5_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5166\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__10809\
        );

    \U712_REG_SM.STATE_COUNTER_4_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5233\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__10809\
        );

    \U712_REG_SM.STATE_COUNTER_6_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4825\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__10809\
        );

    \U712_REG_SM.STATE_COUNTER_3_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6012\,
            in1 => \N__5123\,
            in2 => \N__5066\,
            in3 => \N__5960\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__10809\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4980\,
            in1 => \N__5254\,
            in2 => \_gnd_net_\,
            in3 => \N__5232\,
            lcout => OPEN,
            ltout => \U712_REG_SM.un18_0_i_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__4961\,
            in1 => \N__4999\,
            in2 => \N__5216\,
            in3 => \N__8249\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__10809\
        );

    \U712_REG_SM.STATE_COUNTER_RNIFMLV_8_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__5201\,
            in1 => \N__5053\,
            in2 => \_gnd_net_\,
            in3 => \N__5112\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_442_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CPU_CYCLE_RNO_0_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000111"
        )
    port map (
            in0 => \N__5891\,
            in1 => \N__5171\,
            in2 => \N__5147\,
            in3 => \N__4998\,
            lcout => \U712_REG_SM.REG_CPU_CYCLE_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_0_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100011111"
        )
    port map (
            in0 => \N__5999\,
            in1 => \N__5889\,
            in2 => \N__5063\,
            in3 => \N__5113\,
            lcout => \U712_REG_SM.N_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DBR_SYNC_RNIVIGC1_1_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5958\,
            in1 => \N__5997\,
            in2 => \N__5124\,
            in3 => \N__5046\,
            lcout => \U712_REG_SM.N_447\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__5890\,
            in1 => \N__4981\,
            in2 => \_gnd_net_\,
            in3 => \N__5998\,
            lcout => \U712_REG_SM.N_288\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.LATCH_CLK_0_i_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__6086\,
            in1 => \N__4955\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \LATCH_CLK_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5459\,
            in1 => \N__5441\,
            in2 => \_gnd_net_\,
            in3 => \N__9725\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9726\,
            in1 => \N__9588\,
            in2 => \N__5420\,
            in3 => \N__10442\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5417\,
            in1 => \N__5399\,
            in2 => \_gnd_net_\,
            in3 => \N__9724\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9723\,
            in1 => \N__5384\,
            in2 => \_gnd_net_\,
            in3 => \N__5369\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101001111"
        )
    port map (
            in0 => \N__10036\,
            in1 => \N__10102\,
            in2 => \N__9741\,
            in3 => \N__9589\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5495\,
            in2 => \N__5354\,
            in3 => \N__5351\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9901\,
            ce => \N__9792\,
            sr => \N__10844\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6266\,
            in1 => \N__6299\,
            in2 => \_gnd_net_\,
            in3 => \N__5321\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9901\,
            ce => \N__9792\,
            sr => \N__10844\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10874\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5294\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5288\,
            in1 => \N__5270\,
            in2 => \_gnd_net_\,
            in3 => \N__9702\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10301\,
            in2 => \_gnd_net_\,
            in3 => \N__10211\,
            lcout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\,
            ltout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011110000"
        )
    port map (
            in0 => \N__9590\,
            in1 => \N__10103\,
            in2 => \N__5498\,
            in3 => \N__9703\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011111111111"
        )
    port map (
            in0 => \N__8497\,
            in1 => \N__5465\,
            in2 => \N__7712\,
            in3 => \N__7660\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100011"
        )
    port map (
            in0 => \N__10302\,
            in1 => \N__5519\,
            in2 => \N__6407\,
            in3 => \N__6369\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__5549\,
            in1 => \N__6143\,
            in2 => \N__5540\,
            in3 => \N__6473\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_325_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100000001"
        )
    port map (
            in0 => \N__6398\,
            in1 => \N__6371\,
            in2 => \N__5483\,
            in3 => \N__9714\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011010001"
        )
    port map (
            in0 => \N__5480\,
            in1 => \N__6399\,
            in2 => \N__10224\,
            in3 => \N__6368\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7445\,
            in2 => \_gnd_net_\,
            in3 => \N__7505\,
            lcout => \U712_CHIP_RAM.N_392\,
            ltout => \U712_CHIP_RAM.N_392_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110000"
        )
    port map (
            in0 => \N__7579\,
            in1 => \N__7942\,
            in2 => \N__5468\,
            in3 => \N__7876\,
            lcout => \U712_CHIP_RAM.N_449\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__5536\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5518\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_376_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100000001"
        )
    port map (
            in0 => \N__6370\,
            in1 => \N__6400\,
            in2 => \N__5555\,
            in3 => \N__10260\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9913\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_0_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__7578\,
            in1 => \N__8579\,
            in2 => \N__7658\,
            in3 => \N__6582\,
            lcout => \U712_CHIP_RAM.N_45_i\,
            ltout => \U712_CHIP_RAM.N_45_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNI15FJ4_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8455\,
            in1 => \N__6653\,
            in2 => \N__5552\,
            in3 => \N__7867\,
            lcout => \U712_CHIP_RAM.N_324_2\,
            ltout => \U712_CHIP_RAM.N_324_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__6126\,
            in1 => \N__5624\,
            in2 => \N__5543\,
            in3 => \N__5588\,
            lcout => \U712_CHIP_RAM.N_324\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIFMOI5_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8456\,
            in1 => \N__5507\,
            in2 => \N__7237\,
            in3 => \N__7869\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNILDP34_4_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__7868\,
            in1 => \N__8457\,
            in2 => \N__7954\,
            in3 => \N__7119\,
            lcout => \U712_CHIP_RAM.N_450\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVIFVC_4_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010100000"
        )
    port map (
            in0 => \N__8458\,
            in1 => \N__7946\,
            in2 => \N__7236\,
            in3 => \N__6413\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_RNIVIFVCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__6649\,
            in1 => \N__6133\,
            in2 => \N__5623\,
            in3 => \N__5582\,
            lcout => \U712_CHIP_RAM.N_252\,
            ltout => \U712_CHIP_RAM.N_252_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIURFN4_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5501\,
            in3 => \N__7213\,
            lcout => \U712_CHIP_RAM.N_365_1\,
            ltout => \U712_CHIP_RAM.N_365_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__6668\,
            in1 => \N__7947\,
            in2 => \N__5777\,
            in3 => \N__7881\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10871\,
            in1 => \_gnd_net_\,
            in2 => \N__5774\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110001000"
        )
    port map (
            in0 => \N__8488\,
            in1 => \N__6485\,
            in2 => \N__7342\,
            in3 => \N__6660\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBRn_ibuf_RNIBAB_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5942\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001011111"
        )
    port map (
            in0 => \N__6256\,
            in1 => \_gnd_net_\,
            in2 => \N__6661\,
            in3 => \N__5757\,
            lcout => \U712_CHIP_RAM.N_294\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111111101000000"
        )
    port map (
            in0 => \N__6494\,
            in1 => \N__7711\,
            in2 => \N__6512\,
            in3 => \N__5683\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9919\,
            ce => 'H',
            sr => \N__10810\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011100000101"
        )
    port map (
            in0 => \N__5672\,
            in1 => \N__9483\,
            in2 => \N__5657\,
            in3 => \N__5622\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9919\,
            ce => 'H',
            sr => \N__10810\
        );

    \DBR_SYNC_1_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5561\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9919\,
            ce => 'H',
            sr => \N__10810\
        );

    \DBR_SYNC_0_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5938\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9919\,
            ce => 'H',
            sr => \N__10810\
        );

    \U712_CHIP_RAM.LATCH_RAM_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__6092\,
            in1 => \N__8578\,
            in2 => \N__7341\,
            in3 => \N__6082\,
            lcout => \LATCH_RAM\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9919\,
            ce => 'H',
            sr => \N__10810\
        );

    \U712_REG_SM.STATE_COUNTER_2_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110110000"
        )
    port map (
            in0 => \N__6071\,
            in1 => \N__5959\,
            in2 => \N__6024\,
            in3 => \N__6056\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__10802\
        );

    \U712_REG_SM.DBR_SYNC_1_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5906\,
            lcout => \U712_REG_SM.DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__10802\
        );

    \U712_REG_SM.DBR_SYNC_0_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5931\,
            lcout => \U712_REG_SM.DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__10802\
        );

    \U712_BUFFERS.DMA_LATCH_EN_1_i_m2_i_m2_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__7094\,
            in1 => \N__8005\,
            in2 => \_gnd_net_\,
            in3 => \N__5900\,
            lcout => \N_289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5822\,
            in1 => \N__5804\,
            in2 => \_gnd_net_\,
            in3 => \N__9717\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9718\,
            in1 => \N__9583\,
            in2 => \N__5786\,
            in3 => \N__8690\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9582\,
            in1 => \N__5783\,
            in2 => \N__9740\,
            in3 => \N__8678\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9719\,
            in1 => \N__9584\,
            in2 => \N__6311\,
            in3 => \N__10541\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__10311\,
            in1 => \N__9715\,
            in2 => \_gnd_net_\,
            in3 => \N__10217\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => \U712_CHIP_RAM.CMA_5_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__6286\,
            in1 => \N__9581\,
            in2 => \N__6302\,
            in3 => \N__10354\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9716\,
            in1 => \N__6293\,
            in2 => \N__9598\,
            in3 => \N__9380\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011111111"
        )
    port map (
            in0 => \N__10355\,
            in1 => \N__6287\,
            in2 => \N__9597\,
            in3 => \N__8754\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100111011101110"
        )
    port map (
            in0 => \N__6536\,
            in1 => \N__6941\,
            in2 => \N__7247\,
            in3 => \N__10427\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9902\,
            ce => 'H',
            sr => \N__10830\
        );

    \U712_CHIP_RAM.DBDIR_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111001011110000"
        )
    port map (
            in0 => \N__7241\,
            in1 => \N__6260\,
            in2 => \N__6223\,
            in3 => \N__6563\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9902\,
            ce => 'H',
            sr => \N__10830\
        );

    \U712_CHIP_RAM.REFRESH_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6206\,
            in1 => \N__6191\,
            in2 => \N__6176\,
            in3 => \N__6158\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9907\,
            ce => 'H',
            sr => \N__10822\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKCP34_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__8492\,
            in1 => \N__7877\,
            in2 => \_gnd_net_\,
            in3 => \N__7222\,
            lcout => \U712_CHIP_RAM.N_456\,
            ltout => \U712_CHIP_RAM.N_456_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6397\,
            in2 => \N__6374\,
            in3 => \N__7952\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI8SVVB_3_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__8493\,
            in1 => \N__6902\,
            in2 => \N__7151\,
            in3 => \N__7124\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8580\,
            in2 => \_gnd_net_\,
            in3 => \N__6347\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__6337\,
            in1 => \N__7581\,
            in2 => \N__8634\,
            in3 => \N__6344\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__9911\,
            ce => \N__8509\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__6341\,
            in1 => \N__7462\,
            in2 => \N__8635\,
            in3 => \N__6326\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \N__9911\,
            ce => \N__8509\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__8623\,
            in1 => \N__7515\,
            in2 => \_gnd_net_\,
            in3 => \N__6323\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__9911\,
            ce => \N__8509\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__8629\,
            in1 => \N__7953\,
            in2 => \_gnd_net_\,
            in3 => \N__6320\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__9911\,
            ce => \N__8509\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__8624\,
            in1 => \N__6440\,
            in2 => \_gnd_net_\,
            in3 => \N__6317\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__9911\,
            ce => \N__8509\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__8630\,
            in1 => \N__6452\,
            in2 => \_gnd_net_\,
            in3 => \N__6314\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__9911\,
            ce => \N__8509\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__6464\,
            in1 => \N__8628\,
            in2 => \_gnd_net_\,
            in3 => \N__6476\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9911\,
            ce => \N__8509\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_0_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7641\,
            in1 => \N__7574\,
            in2 => \_gnd_net_\,
            in3 => \N__8557\,
            lcout => \U712_CHIP_RAM.N_388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__6422\,
            in1 => \N__8479\,
            in2 => \N__7886\,
            in3 => \N__7948\,
            lcout => \U712_CHIP_RAM.N_363\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__7856\,
            in1 => \N__7514\,
            in2 => \N__7955\,
            in3 => \N__7123\,
            lcout => \U712_CHIP_RAM.N_351\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6463\,
            in1 => \N__6451\,
            in2 => \_gnd_net_\,
            in3 => \N__6439\,
            lcout => \U712_CHIP_RAM.N_384\,
            ltout => \U712_CHIP_RAM.N_384_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI3PIP2_0_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7455\,
            in1 => \N__7575\,
            in2 => \N__6428\,
            in3 => \N__8558\,
            lcout => \U712_CHIP_RAM.N_400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_0_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7573\,
            in1 => \N__8562\,
            in2 => \_gnd_net_\,
            in3 => \N__7642\,
            lcout => \U712_CHIP_RAM.N_448\,
            ltout => \U712_CHIP_RAM.N_448_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6B326_2_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__7456\,
            in1 => \N__7651\,
            in2 => \N__6425\,
            in3 => \N__7400\,
            lcout => \U712_CHIP_RAM.N_255\,
            ltout => \U712_CHIP_RAM.N_255_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5T4O8_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7855\,
            in2 => \N__6416\,
            in3 => \N__7271\,
            lcout => \U712_CHIP_RAM.N_269\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_3_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__7273\,
            in1 => \N__7776\,
            in2 => \N__6611\,
            in3 => \N__7746\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNI892R_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7857\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6648\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI4LVP1_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7331\,
            in1 => \N__7684\,
            in2 => \_gnd_net_\,
            in3 => \N__7463\,
            lcout => \U712_CHIP_RAM.N_444\,
            ltout => \U712_CHIP_RAM.N_444_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNIFGIT5_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__6595\,
            in1 => \N__7272\,
            in2 => \N__6566\,
            in3 => \N__6559\,
            lcout => \U712_CHIP_RAM.N_334\,
            ltout => \U712_CHIP_RAM.N_334_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNI7SS3A_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__7079\,
            in1 => \N__7464\,
            in2 => \N__6539\,
            in3 => \N__7777\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6527\,
            in3 => \N__10870\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNISH5V3_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__9566\,
            in1 => \N__7747\,
            in2 => \N__6511\,
            in3 => \N__7150\,
            lcout => \U712_CHIP_RAM.N_323\,
            ltout => \U712_CHIP_RAM.N_323_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__7519\,
            in1 => \N__9567\,
            in2 => \N__6488\,
            in3 => \N__7080\,
            lcout => \U712_CHIP_RAM.N_117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8129\,
            in2 => \_gnd_net_\,
            in3 => \N__8122\,
            lcout => \U712_CHIP_RAM.un3_DMA_CYCLE_START\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__10054\,
            in1 => \N__9988\,
            in2 => \N__10151\,
            in3 => \N__6863\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9896\,
            ce => \N__9839\,
            sr => \N__10836\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__10053\,
            in1 => \N__8702\,
            in2 => \N__9996\,
            in3 => \N__6836\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9896\,
            ce => \N__9839\,
            sr => \N__10836\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__10052\,
            in1 => \N__8696\,
            in2 => \N__9995\,
            in3 => \N__6809\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9896\,
            ce => \N__9839\,
            sr => \N__10836\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__9431\,
            in1 => \N__9987\,
            in2 => \N__10058\,
            in3 => \N__6782\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9896\,
            ce => \N__9839\,
            sr => \N__10836\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__6749\,
            in1 => \N__9593\,
            in2 => \N__8764\,
            in3 => \N__10070\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9896\,
            ce => \N__9839\,
            sr => \N__10836\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__10051\,
            in1 => \N__8666\,
            in2 => \N__9997\,
            in3 => \N__6719\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9899\,
            ce => \N__9829\,
            sr => \N__10828\
        );

    \U712_BYTE_ENABLE.N_46_i_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111011101"
        )
    port map (
            in0 => \N__6919\,
            in1 => \N__8107\,
            in2 => \N__6968\,
            in3 => \N__9575\,
            lcout => \N_46_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UUBE_0_a2_0_a2_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__9272\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9093\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.UUBE_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_48_i_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111011101"
        )
    port map (
            in0 => \N__6920\,
            in1 => \N__8056\,
            in2 => \N__7034\,
            in3 => \N__9576\,
            lcout => \N_48_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_49_i_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001011111"
        )
    port map (
            in0 => \N__9577\,
            in1 => \N__8057\,
            in2 => \N__7007\,
            in3 => \N__6995\,
            lcout => \N_49_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UMBE_0_i_o3_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011111010011"
        )
    port map (
            in0 => \N__9092\,
            in1 => \N__9184\,
            in2 => \N__9026\,
            in3 => \N__9271\,
            lcout => \U712_BYTE_ENABLE.N_277\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6942\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7343\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIHC4P1_2_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8460\,
            in1 => \N__7941\,
            in2 => \N__7466\,
            in3 => \N__7839\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__9731\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9520\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIPORK3_1_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8461\,
            in1 => \N__7580\,
            in2 => \N__7707\,
            in3 => \N__7659\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_325_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIE6LO7_1_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6911\,
            in2 => \N__6905\,
            in3 => \N__7277\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__7066\,
            in1 => \N__7854\,
            in2 => \N__6893\,
            in3 => \N__7355\,
            lcout => \WRITE_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9903\,
            ce => 'H',
            sr => \N__10806\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8ALV_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111111"
        )
    port map (
            in0 => \N__7323\,
            in1 => \N__7460\,
            in2 => \_gnd_net_\,
            in3 => \N__7507\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_305_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI8MK44_4_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7940\,
            in1 => \N__7852\,
            in2 => \N__7280\,
            in3 => \N__7270\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_346_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIUHSBF_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__7245\,
            in1 => \N__8432\,
            in2 => \N__7160\,
            in3 => \N__7157\,
            lcout => \U712_CHIP_RAM.N_202\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNITVQE7_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__7143\,
            in1 => \N__7775\,
            in2 => \N__7078\,
            in3 => \N__7117\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_180_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_3_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7939\,
            in2 => \_gnd_net_\,
            in3 => \N__7506\,
            lcout => \U712_CHIP_RAM.N_407\,
            ltout => \U712_CHIP_RAM.N_407_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7853\,
            in2 => \N__7127\,
            in3 => \N__7118\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9903\,
            ce => 'H',
            sr => \N__10806\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7062\,
            in2 => \_gnd_net_\,
            in3 => \N__7454\,
            lcout => \U712_CHIP_RAM.N_257\,
            ltout => \U712_CHIP_RAM.N_257_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100010001"
        )
    port map (
            in0 => \N__8560\,
            in1 => \N__7461\,
            in2 => \N__7037\,
            in3 => \N__7577\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIS3891_3_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__7938\,
            in1 => \N__7504\,
            in2 => \_gnd_net_\,
            in3 => \N__7828\,
            lcout => \U712_CHIP_RAM.N_396\,
            ltout => \U712_CHIP_RAM.N_396_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7576\,
            in1 => \N__8559\,
            in2 => \N__7787\,
            in3 => \N__7643\,
            lcout => \U712_CHIP_RAM.N_436\,
            ltout => \U712_CHIP_RAM.N_436_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7757\,
            in3 => \N__7745\,
            lcout => \U712_CHIP_RAM.N_357\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7718\,
            in1 => \N__7703\,
            in2 => \_gnd_net_\,
            in3 => \N__7644\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__8204\,
            in1 => \N__7601\,
            in2 => \N__7595\,
            in3 => \N__7592\,
            lcout => \CPU_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9909\,
            ce => 'H',
            sr => \N__10800\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__7585\,
            in1 => \N__8561\,
            in2 => \N__7523\,
            in3 => \N__7465\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_63_i_a2_0_0_a2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_2_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__8463\,
            in1 => \N__8358\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_274_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__8194\,
            in1 => \N__7393\,
            in2 => \N__7376\,
            in3 => \N__8257\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_274_i_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7373\,
            in3 => \N__8374\,
            lcout => \U712_CYCLE_TERM.N_274_i_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010101100"
        )
    port map (
            in0 => \N__8660\,
            in1 => \N__8648\,
            in2 => \N__8639\,
            in3 => \N__8594\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9912\,
            ce => \N__8513\,
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8462\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001111"
        )
    port map (
            in0 => \N__8147\,
            in1 => \_gnd_net_\,
            in2 => \N__8363\,
            in3 => \N__8878\,
            lcout => \U712_CYCLE_TERM.N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__8328\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8153\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9914\,
            ce => 'H',
            sr => \N__10799\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__8264\,
            in1 => \N__8154\,
            in2 => \N__8258\,
            in3 => \N__8211\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9914\,
            ce => 'H',
            sr => \N__10799\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8123\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9916\,
            ce => 'H',
            sr => \N__10798\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8094\,
            in2 => \_gnd_net_\,
            in3 => \N__8049\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9916\,
            ce => 'H',
            sr => \N__10798\
        );

    \U712_BUFFERS.un1_DRDENn_0_a2_0_a3_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__8093\,
            in1 => \N__8039\,
            in2 => \_gnd_net_\,
            in3 => \N__8006\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK40_PLL_derived_clock_RNIIOT_0_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8879\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_PLL_iso_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UUBE_i_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9274\,
            in2 => \_gnd_net_\,
            in3 => \N__9084\,
            lcout => \U712_BYTE_ENABLE_UUBE_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__8765\,
            in1 => \N__8738\,
            in2 => \N__9602\,
            in3 => \N__10613\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9897\,
            ce => \N__9833\,
            sr => \N__10848\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__10136\,
            in1 => \_gnd_net_\,
            in2 => \N__11188\,
            in3 => \N__9422\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10943\,
            ce => \N__10914\,
            sr => \N__10845\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9368\,
            in1 => \N__9421\,
            in2 => \_gnd_net_\,
            in3 => \N__11177\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10943\,
            ce => \N__10914\,
            sr => \N__10845\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11183\,
            in1 => \N__9414\,
            in2 => \_gnd_net_\,
            in3 => \N__10134\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            ce => \N__10912\,
            sr => \N__10838\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__10135\,
            in1 => \_gnd_net_\,
            in2 => \N__10697\,
            in3 => \N__11184\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            ce => \N__10912\,
            sr => \N__10838\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9367\,
            in1 => \N__10411\,
            in2 => \_gnd_net_\,
            in3 => \N__11181\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10940\,
            ce => \N__10911\,
            sr => \N__10831\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11182\,
            in1 => \N__10693\,
            in2 => \_gnd_net_\,
            in3 => \N__10529\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10940\,
            ce => \N__10911\,
            sr => \N__10831\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11113\,
            in1 => \N__9360\,
            in2 => \_gnd_net_\,
            in3 => \N__9413\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__10909\,
            sr => \N__10823\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11163\,
            in1 => \N__10410\,
            in2 => \_gnd_net_\,
            in3 => \N__9359\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__10907\,
            sr => \N__10814\
        );

    \U712_BYTE_ENABLE.N_276_i_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101001100"
        )
    port map (
            in0 => \N__9282\,
            in1 => \N__9177\,
            in2 => \N__9108\,
            in3 => \N__9006\,
            lcout => \N_276_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_278_i_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100001011010"
        )
    port map (
            in0 => \N__9179\,
            in1 => \N__9284\,
            in2 => \N__9020\,
            in3 => \N__9104\,
            lcout => \N_278_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_277_i_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011000100"
        )
    port map (
            in0 => \N__9283\,
            in1 => \N__9178\,
            in2 => \N__9109\,
            in3 => \N__9007\,
            lcout => \N_277_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CRCSn_LC_14_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10267\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9895\,
            ce => 'H',
            sr => \N__10854\
        );

    \U712_CHIP_RAM.RASn_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10322\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9895\,
            ce => 'H',
            sr => \N__10854\
        );

    \U712_CHIP_RAM.CASn_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9743\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9898\,
            ce => 'H',
            sr => \N__10853\
        );

    \U712_CHIP_RAM.WEn_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10231\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9898\,
            ce => 'H',
            sr => \N__10853\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__10321\,
            in1 => \N__9742\,
            in2 => \N__10271\,
            in3 => \N__10232\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9900\,
            ce => \N__9837\,
            sr => \N__10849\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10527\,
            in1 => \N__10477\,
            in2 => \_gnd_net_\,
            in3 => \N__11155\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10941\,
            ce => \N__10915\,
            sr => \N__10846\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10125\,
            in1 => \N__10686\,
            in2 => \_gnd_net_\,
            in3 => \N__11154\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10941\,
            ce => \N__10915\,
            sr => \N__10846\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10082\,
            in1 => \N__10600\,
            in2 => \_gnd_net_\,
            in3 => \N__11156\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10941\,
            ce => \N__10915\,
            sr => \N__10846\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__10050\,
            in1 => \N__10952\,
            in2 => \N__9998\,
            in3 => \N__9437\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9908\,
            ce => \N__9838\,
            sr => \N__10839\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9776\,
            in1 => \N__9764\,
            in2 => \_gnd_net_\,
            in3 => \N__9735\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9736\,
            in1 => \N__9568\,
            in2 => \N__9440\,
            in3 => \N__10418\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10685\,
            in1 => \N__10528\,
            in2 => \_gnd_net_\,
            in3 => \N__11099\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__10908\,
            sr => \N__10824\
        );

    \U712_CHIP_RAM.DMA_A20_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__11083\,
            in1 => \N__10646\,
            in2 => \N__10586\,
            in3 => \N__10627\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A20C_net\,
            ce => 'H',
            sr => \N__10815\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10601\,
            in1 => \N__10478\,
            in2 => \_gnd_net_\,
            in3 => \N__11112\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10942\,
            ce => \N__10919\,
            sr => \N__10852\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10599\,
            in1 => \N__10476\,
            in2 => \_gnd_net_\,
            in3 => \N__11153\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__10917\,
            sr => \N__10850\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11152\,
            in1 => \N__10526\,
            in2 => \_gnd_net_\,
            in3 => \N__10459\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__10916\,
            sr => \N__10847\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10996\,
            in1 => \N__11151\,
            in2 => \_gnd_net_\,
            in3 => \N__11021\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__10916\,
            sr => \N__10847\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10412\,
            in1 => \N__10997\,
            in2 => \_gnd_net_\,
            in3 => \N__11150\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__10913\,
            sr => \N__10840\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10991\,
            in1 => \N__10400\,
            in2 => \_gnd_net_\,
            in3 => \N__11087\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10939\,
            ce => \N__10910\,
            sr => \N__10832\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11157\,
            in1 => \N__11020\,
            in2 => \_gnd_net_\,
            in3 => \N__10995\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10938\,
            ce => \N__10918\,
            sr => \N__10851\
        );
end \INTERFACE\;

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jul 1 2025 18:43:57

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U409_TOP" view "INTERFACE"

module U409_TOP (
    ROM_DELAY,
    F_BANK,
    PCIAT,
    TM,
    TT,
    A,
    D,
    PCS0,
    F_ENn,
    TSn,
    SPIO_J,
    SPIO,
    RTC_ENn,
    RESETn,
    OVL,
    F_RDY,
    CONFIGENn,
    PPIO,
    PORTSIZE,
    F_RSTn,
    TICK60,
    PCS1,
    CIACS0n,
    SCS0,
    CPUCONFn,
    CLK6,
    AGNUS_CLK,
    CLK_CIA,
    BUFENn,
    AUTOBOOT,
    RnW,
    XCLK,
    F_WRITEn,
    F_READn,
    CIACS1n,
    PPIO_J,
    TICK50,
    TCIn,
    TBIn,
    RAMSPACEn,
    BPRO_ENn,
    CLK40_IN,
    CLK28_IN,
    XCLK_ENn,
    SCS1,
    REGSPACEn,
    F_WPn,
    ATA_ENn,
    TACKn,
    BREG_ENn,
    ROMENn);

    input [1:0] ROM_DELAY;
    output [1:0] F_BANK;
    output [1:0] PCIAT;
    input [2:0] TM;
    input [1:0] TT;
    input [31:1] A;
    inout [7:4] D;
    output PCS0;
    output F_ENn;
    input TSn;
    input SPIO_J;
    output SPIO;
    output RTC_ENn;
    input RESETn;
    input OVL;
    input F_RDY;
    output CONFIGENn;
    output PPIO;
    output PORTSIZE;
    output F_RSTn;
    output TICK60;
    output PCS1;
    output CIACS0n;
    output SCS0;
    input CPUCONFn;
    input CLK6;
    output AGNUS_CLK;
    output CLK_CIA;
    output BUFENn;
    input AUTOBOOT;
    input RnW;
    input XCLK;
    output F_WRITEn;
    output F_READn;
    output CIACS1n;
    input PPIO_J;
    output TICK50;
    output TCIn;
    output TBIn;
    output RAMSPACEn;
    output BPRO_ENn;
    input CLK40_IN;
    input CLK28_IN;
    input XCLK_ENn;
    output SCS1;
    output REGSPACEn;
    output F_WPn;
    output ATA_ENn;
    inout TACKn;
    output BREG_ENn;
    output ROMENn;

    wire N__13653;
    wire N__13652;
    wire N__13651;
    wire N__13643;
    wire N__13642;
    wire N__13641;
    wire N__13633;
    wire N__13632;
    wire N__13631;
    wire N__13622;
    wire N__13621;
    wire N__13620;
    wire N__13613;
    wire N__13612;
    wire N__13611;
    wire N__13604;
    wire N__13603;
    wire N__13602;
    wire N__13595;
    wire N__13594;
    wire N__13593;
    wire N__13586;
    wire N__13585;
    wire N__13584;
    wire N__13577;
    wire N__13576;
    wire N__13575;
    wire N__13568;
    wire N__13567;
    wire N__13566;
    wire N__13559;
    wire N__13558;
    wire N__13557;
    wire N__13550;
    wire N__13549;
    wire N__13548;
    wire N__13541;
    wire N__13540;
    wire N__13539;
    wire N__13532;
    wire N__13531;
    wire N__13530;
    wire N__13523;
    wire N__13522;
    wire N__13521;
    wire N__13514;
    wire N__13513;
    wire N__13512;
    wire N__13505;
    wire N__13504;
    wire N__13503;
    wire N__13496;
    wire N__13495;
    wire N__13494;
    wire N__13487;
    wire N__13486;
    wire N__13485;
    wire N__13478;
    wire N__13477;
    wire N__13476;
    wire N__13469;
    wire N__13468;
    wire N__13467;
    wire N__13460;
    wire N__13459;
    wire N__13458;
    wire N__13451;
    wire N__13450;
    wire N__13449;
    wire N__13442;
    wire N__13441;
    wire N__13440;
    wire N__13433;
    wire N__13432;
    wire N__13431;
    wire N__13424;
    wire N__13423;
    wire N__13422;
    wire N__13415;
    wire N__13414;
    wire N__13413;
    wire N__13406;
    wire N__13405;
    wire N__13404;
    wire N__13397;
    wire N__13396;
    wire N__13395;
    wire N__13388;
    wire N__13387;
    wire N__13386;
    wire N__13379;
    wire N__13378;
    wire N__13377;
    wire N__13370;
    wire N__13369;
    wire N__13368;
    wire N__13361;
    wire N__13360;
    wire N__13359;
    wire N__13352;
    wire N__13351;
    wire N__13350;
    wire N__13343;
    wire N__13342;
    wire N__13341;
    wire N__13334;
    wire N__13333;
    wire N__13332;
    wire N__13325;
    wire N__13324;
    wire N__13323;
    wire N__13316;
    wire N__13315;
    wire N__13314;
    wire N__13307;
    wire N__13306;
    wire N__13305;
    wire N__13298;
    wire N__13297;
    wire N__13296;
    wire N__13289;
    wire N__13288;
    wire N__13287;
    wire N__13280;
    wire N__13279;
    wire N__13278;
    wire N__13271;
    wire N__13270;
    wire N__13269;
    wire N__13262;
    wire N__13261;
    wire N__13260;
    wire N__13253;
    wire N__13252;
    wire N__13251;
    wire N__13244;
    wire N__13243;
    wire N__13242;
    wire N__13235;
    wire N__13234;
    wire N__13233;
    wire N__13226;
    wire N__13225;
    wire N__13224;
    wire N__13217;
    wire N__13216;
    wire N__13215;
    wire N__13208;
    wire N__13207;
    wire N__13206;
    wire N__13199;
    wire N__13198;
    wire N__13197;
    wire N__13190;
    wire N__13189;
    wire N__13188;
    wire N__13181;
    wire N__13180;
    wire N__13179;
    wire N__13172;
    wire N__13171;
    wire N__13170;
    wire N__13163;
    wire N__13162;
    wire N__13161;
    wire N__13154;
    wire N__13153;
    wire N__13152;
    wire N__13145;
    wire N__13144;
    wire N__13143;
    wire N__13136;
    wire N__13135;
    wire N__13134;
    wire N__13127;
    wire N__13126;
    wire N__13125;
    wire N__13118;
    wire N__13117;
    wire N__13116;
    wire N__13109;
    wire N__13108;
    wire N__13107;
    wire N__13100;
    wire N__13099;
    wire N__13098;
    wire N__13091;
    wire N__13090;
    wire N__13089;
    wire N__13082;
    wire N__13081;
    wire N__13080;
    wire N__13073;
    wire N__13072;
    wire N__13071;
    wire N__13064;
    wire N__13063;
    wire N__13062;
    wire N__13055;
    wire N__13054;
    wire N__13053;
    wire N__13046;
    wire N__13045;
    wire N__13044;
    wire N__13037;
    wire N__13036;
    wire N__13035;
    wire N__13028;
    wire N__13027;
    wire N__13026;
    wire N__13019;
    wire N__13018;
    wire N__13017;
    wire N__13010;
    wire N__13009;
    wire N__13008;
    wire N__13001;
    wire N__13000;
    wire N__12999;
    wire N__12992;
    wire N__12991;
    wire N__12990;
    wire N__12983;
    wire N__12982;
    wire N__12981;
    wire N__12974;
    wire N__12973;
    wire N__12972;
    wire N__12965;
    wire N__12964;
    wire N__12963;
    wire N__12956;
    wire N__12955;
    wire N__12954;
    wire N__12947;
    wire N__12946;
    wire N__12945;
    wire N__12938;
    wire N__12937;
    wire N__12936;
    wire N__12929;
    wire N__12928;
    wire N__12927;
    wire N__12920;
    wire N__12919;
    wire N__12918;
    wire N__12911;
    wire N__12910;
    wire N__12909;
    wire N__12902;
    wire N__12901;
    wire N__12900;
    wire N__12893;
    wire N__12892;
    wire N__12891;
    wire N__12874;
    wire N__12871;
    wire N__12868;
    wire N__12865;
    wire N__12862;
    wire N__12859;
    wire N__12856;
    wire N__12853;
    wire N__12850;
    wire N__12847;
    wire N__12846;
    wire N__12845;
    wire N__12844;
    wire N__12843;
    wire N__12840;
    wire N__12829;
    wire N__12826;
    wire N__12823;
    wire N__12820;
    wire N__12817;
    wire N__12814;
    wire N__12811;
    wire N__12810;
    wire N__12807;
    wire N__12804;
    wire N__12801;
    wire N__12796;
    wire N__12793;
    wire N__12790;
    wire N__12787;
    wire N__12786;
    wire N__12783;
    wire N__12780;
    wire N__12775;
    wire N__12772;
    wire N__12769;
    wire N__12766;
    wire N__12763;
    wire N__12760;
    wire N__12757;
    wire N__12756;
    wire N__12753;
    wire N__12750;
    wire N__12747;
    wire N__12742;
    wire N__12739;
    wire N__12738;
    wire N__12737;
    wire N__12736;
    wire N__12735;
    wire N__12734;
    wire N__12733;
    wire N__12732;
    wire N__12725;
    wire N__12716;
    wire N__12713;
    wire N__12706;
    wire N__12705;
    wire N__12704;
    wire N__12703;
    wire N__12702;
    wire N__12701;
    wire N__12698;
    wire N__12697;
    wire N__12696;
    wire N__12687;
    wire N__12684;
    wire N__12677;
    wire N__12670;
    wire N__12669;
    wire N__12668;
    wire N__12665;
    wire N__12664;
    wire N__12663;
    wire N__12662;
    wire N__12661;
    wire N__12660;
    wire N__12657;
    wire N__12654;
    wire N__12651;
    wire N__12642;
    wire N__12635;
    wire N__12632;
    wire N__12625;
    wire N__12622;
    wire N__12619;
    wire N__12618;
    wire N__12615;
    wire N__12612;
    wire N__12607;
    wire N__12606;
    wire N__12605;
    wire N__12604;
    wire N__12603;
    wire N__12602;
    wire N__12601;
    wire N__12600;
    wire N__12599;
    wire N__12598;
    wire N__12577;
    wire N__12574;
    wire N__12571;
    wire N__12568;
    wire N__12565;
    wire N__12562;
    wire N__12559;
    wire N__12556;
    wire N__12553;
    wire N__12550;
    wire N__12547;
    wire N__12544;
    wire N__12541;
    wire N__12538;
    wire N__12535;
    wire N__12532;
    wire N__12529;
    wire N__12528;
    wire N__12525;
    wire N__12522;
    wire N__12519;
    wire N__12516;
    wire N__12513;
    wire N__12510;
    wire N__12505;
    wire N__12502;
    wire N__12499;
    wire N__12496;
    wire N__12493;
    wire N__12490;
    wire N__12487;
    wire N__12486;
    wire N__12483;
    wire N__12480;
    wire N__12475;
    wire N__12472;
    wire N__12471;
    wire N__12470;
    wire N__12469;
    wire N__12466;
    wire N__12463;
    wire N__12460;
    wire N__12457;
    wire N__12452;
    wire N__12447;
    wire N__12444;
    wire N__12439;
    wire N__12436;
    wire N__12433;
    wire N__12430;
    wire N__12427;
    wire N__12424;
    wire N__12421;
    wire N__12418;
    wire N__12415;
    wire N__12414;
    wire N__12411;
    wire N__12408;
    wire N__12405;
    wire N__12402;
    wire N__12397;
    wire N__12394;
    wire N__12391;
    wire N__12388;
    wire N__12387;
    wire N__12384;
    wire N__12381;
    wire N__12376;
    wire N__12373;
    wire N__12372;
    wire N__12369;
    wire N__12366;
    wire N__12361;
    wire N__12358;
    wire N__12357;
    wire N__12354;
    wire N__12351;
    wire N__12346;
    wire N__12343;
    wire N__12340;
    wire N__12337;
    wire N__12334;
    wire N__12333;
    wire N__12330;
    wire N__12327;
    wire N__12322;
    wire N__12319;
    wire N__12316;
    wire N__12313;
    wire N__12312;
    wire N__12309;
    wire N__12306;
    wire N__12301;
    wire N__12298;
    wire N__12297;
    wire N__12294;
    wire N__12291;
    wire N__12286;
    wire N__12283;
    wire N__12280;
    wire N__12277;
    wire N__12274;
    wire N__12271;
    wire N__12268;
    wire N__12265;
    wire N__12262;
    wire N__12261;
    wire N__12258;
    wire N__12255;
    wire N__12250;
    wire N__12247;
    wire N__12246;
    wire N__12243;
    wire N__12242;
    wire N__12239;
    wire N__12236;
    wire N__12233;
    wire N__12226;
    wire N__12225;
    wire N__12222;
    wire N__12221;
    wire N__12220;
    wire N__12217;
    wire N__12214;
    wire N__12209;
    wire N__12206;
    wire N__12199;
    wire N__12196;
    wire N__12195;
    wire N__12192;
    wire N__12189;
    wire N__12184;
    wire N__12181;
    wire N__12180;
    wire N__12177;
    wire N__12174;
    wire N__12169;
    wire N__12166;
    wire N__12163;
    wire N__12162;
    wire N__12159;
    wire N__12156;
    wire N__12151;
    wire N__12148;
    wire N__12147;
    wire N__12144;
    wire N__12141;
    wire N__12136;
    wire N__12133;
    wire N__12130;
    wire N__12127;
    wire N__12124;
    wire N__12123;
    wire N__12122;
    wire N__12121;
    wire N__12120;
    wire N__12117;
    wire N__12116;
    wire N__12115;
    wire N__12112;
    wire N__12103;
    wire N__12098;
    wire N__12091;
    wire N__12090;
    wire N__12087;
    wire N__12086;
    wire N__12083;
    wire N__12082;
    wire N__12081;
    wire N__12080;
    wire N__12079;
    wire N__12076;
    wire N__12069;
    wire N__12062;
    wire N__12055;
    wire N__12054;
    wire N__12053;
    wire N__12052;
    wire N__12051;
    wire N__12050;
    wire N__12049;
    wire N__12046;
    wire N__12041;
    wire N__12032;
    wire N__12025;
    wire N__12022;
    wire N__12019;
    wire N__12016;
    wire N__12013;
    wire N__12012;
    wire N__12009;
    wire N__12006;
    wire N__12001;
    wire N__12000;
    wire N__11997;
    wire N__11994;
    wire N__11993;
    wire N__11988;
    wire N__11985;
    wire N__11982;
    wire N__11981;
    wire N__11978;
    wire N__11977;
    wire N__11974;
    wire N__11971;
    wire N__11968;
    wire N__11965;
    wire N__11962;
    wire N__11959;
    wire N__11956;
    wire N__11953;
    wire N__11948;
    wire N__11945;
    wire N__11942;
    wire N__11935;
    wire N__11932;
    wire N__11929;
    wire N__11926;
    wire N__11923;
    wire N__11922;
    wire N__11921;
    wire N__11914;
    wire N__11911;
    wire N__11910;
    wire N__11909;
    wire N__11908;
    wire N__11905;
    wire N__11898;
    wire N__11893;
    wire N__11890;
    wire N__11887;
    wire N__11884;
    wire N__11883;
    wire N__11880;
    wire N__11877;
    wire N__11876;
    wire N__11875;
    wire N__11870;
    wire N__11867;
    wire N__11864;
    wire N__11859;
    wire N__11856;
    wire N__11855;
    wire N__11854;
    wire N__11853;
    wire N__11852;
    wire N__11851;
    wire N__11850;
    wire N__11849;
    wire N__11848;
    wire N__11847;
    wire N__11846;
    wire N__11843;
    wire N__11842;
    wire N__11839;
    wire N__11838;
    wire N__11837;
    wire N__11836;
    wire N__11829;
    wire N__11826;
    wire N__11821;
    wire N__11816;
    wire N__11815;
    wire N__11810;
    wire N__11809;
    wire N__11806;
    wire N__11803;
    wire N__11800;
    wire N__11797;
    wire N__11796;
    wire N__11795;
    wire N__11792;
    wire N__11789;
    wire N__11788;
    wire N__11779;
    wire N__11776;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11764;
    wire N__11759;
    wire N__11756;
    wire N__11753;
    wire N__11750;
    wire N__11745;
    wire N__11740;
    wire N__11739;
    wire N__11738;
    wire N__11735;
    wire N__11732;
    wire N__11731;
    wire N__11728;
    wire N__11725;
    wire N__11722;
    wire N__11719;
    wire N__11716;
    wire N__11711;
    wire N__11708;
    wire N__11701;
    wire N__11698;
    wire N__11695;
    wire N__11692;
    wire N__11687;
    wire N__11672;
    wire N__11669;
    wire N__11666;
    wire N__11663;
    wire N__11660;
    wire N__11655;
    wire N__11650;
    wire N__11649;
    wire N__11648;
    wire N__11645;
    wire N__11640;
    wire N__11637;
    wire N__11632;
    wire N__11629;
    wire N__11628;
    wire N__11627;
    wire N__11626;
    wire N__11625;
    wire N__11622;
    wire N__11619;
    wire N__11616;
    wire N__11607;
    wire N__11602;
    wire N__11601;
    wire N__11596;
    wire N__11593;
    wire N__11590;
    wire N__11587;
    wire N__11586;
    wire N__11583;
    wire N__11580;
    wire N__11577;
    wire N__11574;
    wire N__11573;
    wire N__11570;
    wire N__11567;
    wire N__11566;
    wire N__11563;
    wire N__11560;
    wire N__11557;
    wire N__11554;
    wire N__11551;
    wire N__11542;
    wire N__11541;
    wire N__11540;
    wire N__11537;
    wire N__11532;
    wire N__11527;
    wire N__11524;
    wire N__11521;
    wire N__11518;
    wire N__11515;
    wire N__11512;
    wire N__11509;
    wire N__11506;
    wire N__11505;
    wire N__11502;
    wire N__11499;
    wire N__11498;
    wire N__11497;
    wire N__11494;
    wire N__11491;
    wire N__11488;
    wire N__11485;
    wire N__11482;
    wire N__11479;
    wire N__11476;
    wire N__11473;
    wire N__11464;
    wire N__11463;
    wire N__11460;
    wire N__11459;
    wire N__11458;
    wire N__11455;
    wire N__11452;
    wire N__11447;
    wire N__11440;
    wire N__11437;
    wire N__11436;
    wire N__11435;
    wire N__11434;
    wire N__11431;
    wire N__11430;
    wire N__11429;
    wire N__11426;
    wire N__11421;
    wire N__11420;
    wire N__11417;
    wire N__11412;
    wire N__11407;
    wire N__11404;
    wire N__11395;
    wire N__11394;
    wire N__11393;
    wire N__11392;
    wire N__11391;
    wire N__11390;
    wire N__11389;
    wire N__11388;
    wire N__11387;
    wire N__11386;
    wire N__11385;
    wire N__11384;
    wire N__11383;
    wire N__11382;
    wire N__11353;
    wire N__11350;
    wire N__11347;
    wire N__11346;
    wire N__11343;
    wire N__11340;
    wire N__11335;
    wire N__11334;
    wire N__11331;
    wire N__11328;
    wire N__11323;
    wire N__11320;
    wire N__11319;
    wire N__11316;
    wire N__11315;
    wire N__11312;
    wire N__11309;
    wire N__11306;
    wire N__11299;
    wire N__11298;
    wire N__11295;
    wire N__11292;
    wire N__11287;
    wire N__11284;
    wire N__11281;
    wire N__11280;
    wire N__11277;
    wire N__11274;
    wire N__11269;
    wire N__11266;
    wire N__11265;
    wire N__11262;
    wire N__11259;
    wire N__11254;
    wire N__11251;
    wire N__11248;
    wire N__11245;
    wire N__11244;
    wire N__11241;
    wire N__11238;
    wire N__11233;
    wire N__11230;
    wire N__11227;
    wire N__11224;
    wire N__11221;
    wire N__11220;
    wire N__11217;
    wire N__11214;
    wire N__11209;
    wire N__11206;
    wire N__11205;
    wire N__11204;
    wire N__11203;
    wire N__11202;
    wire N__11199;
    wire N__11196;
    wire N__11191;
    wire N__11188;
    wire N__11187;
    wire N__11184;
    wire N__11183;
    wire N__11182;
    wire N__11181;
    wire N__11180;
    wire N__11179;
    wire N__11176;
    wire N__11175;
    wire N__11174;
    wire N__11173;
    wire N__11172;
    wire N__11171;
    wire N__11170;
    wire N__11169;
    wire N__11166;
    wire N__11165;
    wire N__11162;
    wire N__11161;
    wire N__11122;
    wire N__11119;
    wire N__11116;
    wire N__11115;
    wire N__11112;
    wire N__11109;
    wire N__11104;
    wire N__11101;
    wire N__11098;
    wire N__11095;
    wire N__11092;
    wire N__11089;
    wire N__11086;
    wire N__11085;
    wire N__11082;
    wire N__11079;
    wire N__11074;
    wire N__11071;
    wire N__11068;
    wire N__11067;
    wire N__11064;
    wire N__11061;
    wire N__11056;
    wire N__11055;
    wire N__11052;
    wire N__11049;
    wire N__11044;
    wire N__11043;
    wire N__11040;
    wire N__11037;
    wire N__11034;
    wire N__11029;
    wire N__11026;
    wire N__11023;
    wire N__11020;
    wire N__11017;
    wire N__11016;
    wire N__11013;
    wire N__11010;
    wire N__11005;
    wire N__11004;
    wire N__11001;
    wire N__10998;
    wire N__10993;
    wire N__10992;
    wire N__10989;
    wire N__10986;
    wire N__10981;
    wire N__10978;
    wire N__10977;
    wire N__10974;
    wire N__10971;
    wire N__10966;
    wire N__10963;
    wire N__10962;
    wire N__10961;
    wire N__10960;
    wire N__10957;
    wire N__10954;
    wire N__10949;
    wire N__10946;
    wire N__10939;
    wire N__10938;
    wire N__10935;
    wire N__10932;
    wire N__10929;
    wire N__10924;
    wire N__10923;
    wire N__10920;
    wire N__10917;
    wire N__10914;
    wire N__10911;
    wire N__10908;
    wire N__10905;
    wire N__10904;
    wire N__10901;
    wire N__10898;
    wire N__10895;
    wire N__10888;
    wire N__10887;
    wire N__10884;
    wire N__10881;
    wire N__10878;
    wire N__10875;
    wire N__10870;
    wire N__10867;
    wire N__10864;
    wire N__10861;
    wire N__10860;
    wire N__10859;
    wire N__10858;
    wire N__10855;
    wire N__10852;
    wire N__10851;
    wire N__10850;
    wire N__10849;
    wire N__10848;
    wire N__10845;
    wire N__10842;
    wire N__10839;
    wire N__10834;
    wire N__10829;
    wire N__10826;
    wire N__10813;
    wire N__10812;
    wire N__10809;
    wire N__10808;
    wire N__10807;
    wire N__10806;
    wire N__10805;
    wire N__10802;
    wire N__10799;
    wire N__10796;
    wire N__10795;
    wire N__10792;
    wire N__10789;
    wire N__10786;
    wire N__10783;
    wire N__10780;
    wire N__10777;
    wire N__10774;
    wire N__10759;
    wire N__10758;
    wire N__10757;
    wire N__10756;
    wire N__10755;
    wire N__10754;
    wire N__10751;
    wire N__10748;
    wire N__10745;
    wire N__10742;
    wire N__10737;
    wire N__10726;
    wire N__10723;
    wire N__10720;
    wire N__10717;
    wire N__10716;
    wire N__10715;
    wire N__10712;
    wire N__10709;
    wire N__10708;
    wire N__10707;
    wire N__10704;
    wire N__10701;
    wire N__10698;
    wire N__10695;
    wire N__10692;
    wire N__10687;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10668;
    wire N__10665;
    wire N__10662;
    wire N__10659;
    wire N__10656;
    wire N__10653;
    wire N__10648;
    wire N__10647;
    wire N__10646;
    wire N__10641;
    wire N__10638;
    wire N__10637;
    wire N__10632;
    wire N__10629;
    wire N__10628;
    wire N__10623;
    wire N__10620;
    wire N__10615;
    wire N__10612;
    wire N__10609;
    wire N__10606;
    wire N__10603;
    wire N__10602;
    wire N__10599;
    wire N__10596;
    wire N__10593;
    wire N__10588;
    wire N__10585;
    wire N__10582;
    wire N__10579;
    wire N__10576;
    wire N__10573;
    wire N__10570;
    wire N__10567;
    wire N__10564;
    wire N__10561;
    wire N__10558;
    wire N__10555;
    wire N__10552;
    wire N__10549;
    wire N__10546;
    wire N__10543;
    wire N__10540;
    wire N__10537;
    wire N__10534;
    wire N__10533;
    wire N__10530;
    wire N__10527;
    wire N__10522;
    wire N__10519;
    wire N__10516;
    wire N__10513;
    wire N__10510;
    wire N__10509;
    wire N__10506;
    wire N__10503;
    wire N__10498;
    wire N__10495;
    wire N__10492;
    wire N__10489;
    wire N__10486;
    wire N__10483;
    wire N__10482;
    wire N__10479;
    wire N__10476;
    wire N__10471;
    wire N__10468;
    wire N__10465;
    wire N__10462;
    wire N__10459;
    wire N__10456;
    wire N__10453;
    wire N__10450;
    wire N__10447;
    wire N__10444;
    wire N__10441;
    wire N__10438;
    wire N__10435;
    wire N__10432;
    wire N__10429;
    wire N__10426;
    wire N__10425;
    wire N__10420;
    wire N__10417;
    wire N__10414;
    wire N__10411;
    wire N__10408;
    wire N__10407;
    wire N__10404;
    wire N__10401;
    wire N__10396;
    wire N__10395;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10376;
    wire N__10373;
    wire N__10370;
    wire N__10367;
    wire N__10362;
    wire N__10359;
    wire N__10354;
    wire N__10351;
    wire N__10348;
    wire N__10347;
    wire N__10344;
    wire N__10341;
    wire N__10336;
    wire N__10333;
    wire N__10332;
    wire N__10329;
    wire N__10326;
    wire N__10321;
    wire N__10318;
    wire N__10315;
    wire N__10314;
    wire N__10311;
    wire N__10308;
    wire N__10303;
    wire N__10300;
    wire N__10297;
    wire N__10294;
    wire N__10291;
    wire N__10288;
    wire N__10285;
    wire N__10282;
    wire N__10279;
    wire N__10276;
    wire N__10275;
    wire N__10272;
    wire N__10269;
    wire N__10264;
    wire N__10261;
    wire N__10258;
    wire N__10255;
    wire N__10252;
    wire N__10249;
    wire N__10246;
    wire N__10245;
    wire N__10242;
    wire N__10239;
    wire N__10234;
    wire N__10231;
    wire N__10228;
    wire N__10225;
    wire N__10222;
    wire N__10219;
    wire N__10218;
    wire N__10215;
    wire N__10214;
    wire N__10213;
    wire N__10210;
    wire N__10209;
    wire N__10206;
    wire N__10203;
    wire N__10198;
    wire N__10195;
    wire N__10194;
    wire N__10191;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10181;
    wire N__10178;
    wire N__10175;
    wire N__10174;
    wire N__10171;
    wire N__10168;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10143;
    wire N__10138;
    wire N__10135;
    wire N__10132;
    wire N__10129;
    wire N__10126;
    wire N__10123;
    wire N__10116;
    wire N__10111;
    wire N__10110;
    wire N__10109;
    wire N__10108;
    wire N__10107;
    wire N__10104;
    wire N__10101;
    wire N__10100;
    wire N__10097;
    wire N__10094;
    wire N__10091;
    wire N__10090;
    wire N__10085;
    wire N__10082;
    wire N__10079;
    wire N__10074;
    wire N__10071;
    wire N__10068;
    wire N__10065;
    wire N__10062;
    wire N__10057;
    wire N__10054;
    wire N__10051;
    wire N__10046;
    wire N__10045;
    wire N__10042;
    wire N__10037;
    wire N__10034;
    wire N__10027;
    wire N__10024;
    wire N__10021;
    wire N__10018;
    wire N__10017;
    wire N__10016;
    wire N__10013;
    wire N__10012;
    wire N__10011;
    wire N__10010;
    wire N__10009;
    wire N__10006;
    wire N__10005;
    wire N__10002;
    wire N__9999;
    wire N__9996;
    wire N__9993;
    wire N__9990;
    wire N__9987;
    wire N__9984;
    wire N__9981;
    wire N__9978;
    wire N__9975;
    wire N__9974;
    wire N__9969;
    wire N__9966;
    wire N__9963;
    wire N__9960;
    wire N__9957;
    wire N__9954;
    wire N__9951;
    wire N__9948;
    wire N__9943;
    wire N__9930;
    wire N__9927;
    wire N__9924;
    wire N__9919;
    wire N__9916;
    wire N__9915;
    wire N__9914;
    wire N__9913;
    wire N__9912;
    wire N__9909;
    wire N__9906;
    wire N__9903;
    wire N__9900;
    wire N__9899;
    wire N__9896;
    wire N__9895;
    wire N__9892;
    wire N__9889;
    wire N__9886;
    wire N__9883;
    wire N__9880;
    wire N__9877;
    wire N__9874;
    wire N__9871;
    wire N__9868;
    wire N__9867;
    wire N__9864;
    wire N__9861;
    wire N__9854;
    wire N__9851;
    wire N__9848;
    wire N__9845;
    wire N__9840;
    wire N__9837;
    wire N__9834;
    wire N__9831;
    wire N__9828;
    wire N__9825;
    wire N__9822;
    wire N__9819;
    wire N__9816;
    wire N__9813;
    wire N__9808;
    wire N__9801;
    wire N__9796;
    wire N__9795;
    wire N__9792;
    wire N__9789;
    wire N__9786;
    wire N__9785;
    wire N__9782;
    wire N__9779;
    wire N__9776;
    wire N__9769;
    wire N__9766;
    wire N__9763;
    wire N__9760;
    wire N__9759;
    wire N__9758;
    wire N__9755;
    wire N__9754;
    wire N__9751;
    wire N__9748;
    wire N__9745;
    wire N__9744;
    wire N__9741;
    wire N__9740;
    wire N__9733;
    wire N__9730;
    wire N__9729;
    wire N__9728;
    wire N__9725;
    wire N__9724;
    wire N__9723;
    wire N__9720;
    wire N__9715;
    wire N__9712;
    wire N__9709;
    wire N__9708;
    wire N__9705;
    wire N__9702;
    wire N__9699;
    wire N__9698;
    wire N__9695;
    wire N__9690;
    wire N__9687;
    wire N__9684;
    wire N__9683;
    wire N__9676;
    wire N__9673;
    wire N__9668;
    wire N__9665;
    wire N__9662;
    wire N__9659;
    wire N__9656;
    wire N__9653;
    wire N__9646;
    wire N__9643;
    wire N__9640;
    wire N__9637;
    wire N__9632;
    wire N__9625;
    wire N__9622;
    wire N__9619;
    wire N__9616;
    wire N__9613;
    wire N__9610;
    wire N__9607;
    wire N__9604;
    wire N__9603;
    wire N__9600;
    wire N__9597;
    wire N__9594;
    wire N__9591;
    wire N__9590;
    wire N__9589;
    wire N__9586;
    wire N__9583;
    wire N__9580;
    wire N__9577;
    wire N__9574;
    wire N__9569;
    wire N__9566;
    wire N__9559;
    wire N__9556;
    wire N__9553;
    wire N__9550;
    wire N__9547;
    wire N__9544;
    wire N__9541;
    wire N__9538;
    wire N__9535;
    wire N__9532;
    wire N__9529;
    wire N__9526;
    wire N__9523;
    wire N__9522;
    wire N__9519;
    wire N__9516;
    wire N__9513;
    wire N__9508;
    wire N__9505;
    wire N__9502;
    wire N__9499;
    wire N__9498;
    wire N__9495;
    wire N__9492;
    wire N__9491;
    wire N__9486;
    wire N__9483;
    wire N__9480;
    wire N__9477;
    wire N__9474;
    wire N__9471;
    wire N__9470;
    wire N__9469;
    wire N__9466;
    wire N__9463;
    wire N__9458;
    wire N__9451;
    wire N__9450;
    wire N__9449;
    wire N__9448;
    wire N__9445;
    wire N__9438;
    wire N__9433;
    wire N__9432;
    wire N__9431;
    wire N__9430;
    wire N__9427;
    wire N__9420;
    wire N__9415;
    wire N__9414;
    wire N__9411;
    wire N__9408;
    wire N__9403;
    wire N__9400;
    wire N__9399;
    wire N__9398;
    wire N__9397;
    wire N__9396;
    wire N__9395;
    wire N__9392;
    wire N__9389;
    wire N__9388;
    wire N__9385;
    wire N__9382;
    wire N__9379;
    wire N__9376;
    wire N__9375;
    wire N__9370;
    wire N__9367;
    wire N__9364;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9352;
    wire N__9347;
    wire N__9340;
    wire N__9337;
    wire N__9334;
    wire N__9331;
    wire N__9324;
    wire N__9321;
    wire N__9318;
    wire N__9315;
    wire N__9312;
    wire N__9307;
    wire N__9304;
    wire N__9301;
    wire N__9298;
    wire N__9297;
    wire N__9296;
    wire N__9293;
    wire N__9288;
    wire N__9285;
    wire N__9284;
    wire N__9283;
    wire N__9280;
    wire N__9277;
    wire N__9274;
    wire N__9271;
    wire N__9268;
    wire N__9263;
    wire N__9260;
    wire N__9255;
    wire N__9252;
    wire N__9249;
    wire N__9246;
    wire N__9241;
    wire N__9238;
    wire N__9237;
    wire N__9232;
    wire N__9229;
    wire N__9226;
    wire N__9223;
    wire N__9220;
    wire N__9217;
    wire N__9216;
    wire N__9215;
    wire N__9212;
    wire N__9209;
    wire N__9206;
    wire N__9203;
    wire N__9198;
    wire N__9193;
    wire N__9190;
    wire N__9187;
    wire N__9184;
    wire N__9181;
    wire N__9178;
    wire N__9175;
    wire N__9172;
    wire N__9169;
    wire N__9166;
    wire N__9163;
    wire N__9160;
    wire N__9157;
    wire N__9154;
    wire N__9151;
    wire N__9150;
    wire N__9145;
    wire N__9142;
    wire N__9141;
    wire N__9138;
    wire N__9135;
    wire N__9130;
    wire N__9127;
    wire N__9124;
    wire N__9121;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9109;
    wire N__9106;
    wire N__9103;
    wire N__9100;
    wire N__9097;
    wire N__9096;
    wire N__9093;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9082;
    wire N__9079;
    wire N__9076;
    wire N__9073;
    wire N__9070;
    wire N__9067;
    wire N__9064;
    wire N__9061;
    wire N__9058;
    wire N__9049;
    wire N__9046;
    wire N__9043;
    wire N__9040;
    wire N__9037;
    wire N__9034;
    wire N__9031;
    wire N__9028;
    wire N__9025;
    wire N__9022;
    wire N__9019;
    wire N__9018;
    wire N__9015;
    wire N__9012;
    wire N__9009;
    wire N__9006;
    wire N__9001;
    wire N__8998;
    wire N__8995;
    wire N__8992;
    wire N__8989;
    wire N__8986;
    wire N__8983;
    wire N__8980;
    wire N__8979;
    wire N__8978;
    wire N__8977;
    wire N__8976;
    wire N__8973;
    wire N__8968;
    wire N__8965;
    wire N__8962;
    wire N__8953;
    wire N__8950;
    wire N__8947;
    wire N__8944;
    wire N__8943;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8926;
    wire N__8923;
    wire N__8920;
    wire N__8919;
    wire N__8916;
    wire N__8913;
    wire N__8910;
    wire N__8905;
    wire N__8904;
    wire N__8903;
    wire N__8902;
    wire N__8899;
    wire N__8896;
    wire N__8895;
    wire N__8892;
    wire N__8891;
    wire N__8888;
    wire N__8883;
    wire N__8876;
    wire N__8869;
    wire N__8868;
    wire N__8867;
    wire N__8866;
    wire N__8863;
    wire N__8860;
    wire N__8857;
    wire N__8856;
    wire N__8853;
    wire N__8850;
    wire N__8847;
    wire N__8844;
    wire N__8841;
    wire N__8838;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8826;
    wire N__8823;
    wire N__8820;
    wire N__8817;
    wire N__8814;
    wire N__8811;
    wire N__8806;
    wire N__8799;
    wire N__8796;
    wire N__8793;
    wire N__8790;
    wire N__8787;
    wire N__8782;
    wire N__8779;
    wire N__8778;
    wire N__8777;
    wire N__8774;
    wire N__8771;
    wire N__8770;
    wire N__8769;
    wire N__8768;
    wire N__8765;
    wire N__8762;
    wire N__8759;
    wire N__8752;
    wire N__8743;
    wire N__8742;
    wire N__8739;
    wire N__8736;
    wire N__8733;
    wire N__8730;
    wire N__8727;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8710;
    wire N__8707;
    wire N__8704;
    wire N__8701;
    wire N__8698;
    wire N__8695;
    wire N__8692;
    wire N__8689;
    wire N__8688;
    wire N__8685;
    wire N__8682;
    wire N__8677;
    wire N__8674;
    wire N__8673;
    wire N__8670;
    wire N__8667;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8656;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8638;
    wire N__8635;
    wire N__8632;
    wire N__8629;
    wire N__8626;
    wire N__8623;
    wire N__8622;
    wire N__8621;
    wire N__8620;
    wire N__8619;
    wire N__8616;
    wire N__8609;
    wire N__8604;
    wire N__8599;
    wire N__8596;
    wire N__8595;
    wire N__8592;
    wire N__8591;
    wire N__8590;
    wire N__8587;
    wire N__8586;
    wire N__8579;
    wire N__8574;
    wire N__8569;
    wire N__8568;
    wire N__8567;
    wire N__8566;
    wire N__8565;
    wire N__8560;
    wire N__8553;
    wire N__8548;
    wire N__8545;
    wire N__8544;
    wire N__8543;
    wire N__8542;
    wire N__8539;
    wire N__8536;
    wire N__8533;
    wire N__8532;
    wire N__8529;
    wire N__8524;
    wire N__8521;
    wire N__8518;
    wire N__8515;
    wire N__8508;
    wire N__8503;
    wire N__8500;
    wire N__8497;
    wire N__8496;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8481;
    wire N__8478;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8463;
    wire N__8460;
    wire N__8455;
    wire N__8454;
    wire N__8451;
    wire N__8448;
    wire N__8443;
    wire N__8440;
    wire N__8439;
    wire N__8436;
    wire N__8433;
    wire N__8428;
    wire N__8425;
    wire N__8422;
    wire N__8421;
    wire N__8418;
    wire N__8417;
    wire N__8414;
    wire N__8413;
    wire N__8410;
    wire N__8407;
    wire N__8404;
    wire N__8401;
    wire N__8398;
    wire N__8391;
    wire N__8390;
    wire N__8385;
    wire N__8382;
    wire N__8377;
    wire N__8374;
    wire N__8371;
    wire N__8368;
    wire N__8365;
    wire N__8362;
    wire N__8359;
    wire N__8358;
    wire N__8357;
    wire N__8352;
    wire N__8349;
    wire N__8344;
    wire N__8343;
    wire N__8342;
    wire N__8339;
    wire N__8334;
    wire N__8329;
    wire N__8326;
    wire N__8323;
    wire N__8320;
    wire N__8317;
    wire N__8314;
    wire N__8311;
    wire N__8310;
    wire N__8309;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8299;
    wire N__8294;
    wire N__8287;
    wire N__8284;
    wire N__8283;
    wire N__8278;
    wire N__8275;
    wire N__8274;
    wire N__8273;
    wire N__8270;
    wire N__8269;
    wire N__8264;
    wire N__8259;
    wire N__8254;
    wire N__8251;
    wire N__8248;
    wire N__8245;
    wire N__8244;
    wire N__8243;
    wire N__8242;
    wire N__8239;
    wire N__8236;
    wire N__8231;
    wire N__8224;
    wire N__8223;
    wire N__8222;
    wire N__8221;
    wire N__8218;
    wire N__8211;
    wire N__8206;
    wire N__8205;
    wire N__8202;
    wire N__8199;
    wire N__8196;
    wire N__8191;
    wire N__8190;
    wire N__8189;
    wire N__8188;
    wire N__8187;
    wire N__8184;
    wire N__8181;
    wire N__8178;
    wire N__8173;
    wire N__8164;
    wire N__8161;
    wire N__8160;
    wire N__8155;
    wire N__8152;
    wire N__8149;
    wire N__8148;
    wire N__8147;
    wire N__8144;
    wire N__8139;
    wire N__8138;
    wire N__8137;
    wire N__8134;
    wire N__8131;
    wire N__8128;
    wire N__8125;
    wire N__8120;
    wire N__8115;
    wire N__8110;
    wire N__8107;
    wire N__8104;
    wire N__8101;
    wire N__8098;
    wire N__8097;
    wire N__8094;
    wire N__8091;
    wire N__8088;
    wire N__8085;
    wire N__8080;
    wire N__8077;
    wire N__8076;
    wire N__8073;
    wire N__8070;
    wire N__8067;
    wire N__8062;
    wire N__8061;
    wire N__8058;
    wire N__8055;
    wire N__8052;
    wire N__8049;
    wire N__8048;
    wire N__8047;
    wire N__8046;
    wire N__8043;
    wire N__8040;
    wire N__8033;
    wire N__8030;
    wire N__8025;
    wire N__8020;
    wire N__8017;
    wire N__8014;
    wire N__8013;
    wire N__8012;
    wire N__8011;
    wire N__8008;
    wire N__8003;
    wire N__8000;
    wire N__7993;
    wire N__7990;
    wire N__7989;
    wire N__7986;
    wire N__7983;
    wire N__7980;
    wire N__7977;
    wire N__7972;
    wire N__7971;
    wire N__7970;
    wire N__7969;
    wire N__7964;
    wire N__7959;
    wire N__7954;
    wire N__7953;
    wire N__7952;
    wire N__7949;
    wire N__7946;
    wire N__7943;
    wire N__7940;
    wire N__7937;
    wire N__7930;
    wire N__7927;
    wire N__7924;
    wire N__7921;
    wire N__7918;
    wire N__7917;
    wire N__7914;
    wire N__7911;
    wire N__7910;
    wire N__7909;
    wire N__7908;
    wire N__7907;
    wire N__7906;
    wire N__7905;
    wire N__7904;
    wire N__7891;
    wire N__7890;
    wire N__7889;
    wire N__7888;
    wire N__7881;
    wire N__7878;
    wire N__7877;
    wire N__7876;
    wire N__7875;
    wire N__7874;
    wire N__7873;
    wire N__7866;
    wire N__7865;
    wire N__7862;
    wire N__7859;
    wire N__7854;
    wire N__7847;
    wire N__7844;
    wire N__7841;
    wire N__7832;
    wire N__7825;
    wire N__7822;
    wire N__7819;
    wire N__7816;
    wire N__7813;
    wire N__7810;
    wire N__7809;
    wire N__7806;
    wire N__7805;
    wire N__7802;
    wire N__7799;
    wire N__7798;
    wire N__7797;
    wire N__7794;
    wire N__7791;
    wire N__7788;
    wire N__7783;
    wire N__7780;
    wire N__7777;
    wire N__7774;
    wire N__7771;
    wire N__7768;
    wire N__7765;
    wire N__7762;
    wire N__7759;
    wire N__7754;
    wire N__7747;
    wire N__7746;
    wire N__7743;
    wire N__7740;
    wire N__7735;
    wire N__7734;
    wire N__7733;
    wire N__7732;
    wire N__7729;
    wire N__7724;
    wire N__7723;
    wire N__7720;
    wire N__7717;
    wire N__7714;
    wire N__7711;
    wire N__7710;
    wire N__7707;
    wire N__7704;
    wire N__7701;
    wire N__7698;
    wire N__7695;
    wire N__7692;
    wire N__7689;
    wire N__7686;
    wire N__7681;
    wire N__7678;
    wire N__7675;
    wire N__7670;
    wire N__7667;
    wire N__7662;
    wire N__7657;
    wire N__7654;
    wire N__7653;
    wire N__7650;
    wire N__7647;
    wire N__7642;
    wire N__7639;
    wire N__7636;
    wire N__7635;
    wire N__7632;
    wire N__7631;
    wire N__7626;
    wire N__7625;
    wire N__7624;
    wire N__7621;
    wire N__7620;
    wire N__7617;
    wire N__7614;
    wire N__7613;
    wire N__7612;
    wire N__7609;
    wire N__7608;
    wire N__7605;
    wire N__7602;
    wire N__7597;
    wire N__7594;
    wire N__7591;
    wire N__7588;
    wire N__7585;
    wire N__7570;
    wire N__7567;
    wire N__7564;
    wire N__7561;
    wire N__7560;
    wire N__7557;
    wire N__7554;
    wire N__7549;
    wire N__7548;
    wire N__7545;
    wire N__7542;
    wire N__7537;
    wire N__7534;
    wire N__7531;
    wire N__7530;
    wire N__7529;
    wire N__7526;
    wire N__7521;
    wire N__7516;
    wire N__7513;
    wire N__7512;
    wire N__7509;
    wire N__7506;
    wire N__7503;
    wire N__7500;
    wire N__7495;
    wire N__7494;
    wire N__7493;
    wire N__7490;
    wire N__7485;
    wire N__7482;
    wire N__7477;
    wire N__7474;
    wire N__7471;
    wire N__7468;
    wire N__7467;
    wire N__7464;
    wire N__7461;
    wire N__7456;
    wire N__7455;
    wire N__7452;
    wire N__7451;
    wire N__7450;
    wire N__7449;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7439;
    wire N__7438;
    wire N__7437;
    wire N__7436;
    wire N__7435;
    wire N__7432;
    wire N__7429;
    wire N__7428;
    wire N__7427;
    wire N__7424;
    wire N__7417;
    wire N__7408;
    wire N__7407;
    wire N__7406;
    wire N__7403;
    wire N__7400;
    wire N__7397;
    wire N__7394;
    wire N__7387;
    wire N__7384;
    wire N__7381;
    wire N__7366;
    wire N__7363;
    wire N__7360;
    wire N__7359;
    wire N__7358;
    wire N__7357;
    wire N__7354;
    wire N__7351;
    wire N__7346;
    wire N__7339;
    wire N__7338;
    wire N__7337;
    wire N__7336;
    wire N__7333;
    wire N__7330;
    wire N__7327;
    wire N__7324;
    wire N__7321;
    wire N__7312;
    wire N__7311;
    wire N__7308;
    wire N__7307;
    wire N__7306;
    wire N__7303;
    wire N__7300;
    wire N__7297;
    wire N__7294;
    wire N__7285;
    wire N__7284;
    wire N__7283;
    wire N__7282;
    wire N__7279;
    wire N__7276;
    wire N__7271;
    wire N__7264;
    wire N__7261;
    wire N__7260;
    wire N__7255;
    wire N__7252;
    wire N__7251;
    wire N__7250;
    wire N__7249;
    wire N__7248;
    wire N__7247;
    wire N__7242;
    wire N__7233;
    wire N__7228;
    wire N__7227;
    wire N__7226;
    wire N__7225;
    wire N__7224;
    wire N__7221;
    wire N__7218;
    wire N__7215;
    wire N__7214;
    wire N__7211;
    wire N__7206;
    wire N__7199;
    wire N__7192;
    wire N__7191;
    wire N__7188;
    wire N__7187;
    wire N__7182;
    wire N__7179;
    wire N__7174;
    wire N__7173;
    wire N__7172;
    wire N__7167;
    wire N__7164;
    wire N__7159;
    wire N__7158;
    wire N__7155;
    wire N__7152;
    wire N__7147;
    wire N__7144;
    wire N__7141;
    wire N__7138;
    wire N__7135;
    wire N__7132;
    wire N__7129;
    wire N__7126;
    wire N__7123;
    wire N__7120;
    wire N__7117;
    wire N__7116;
    wire N__7113;
    wire N__7110;
    wire N__7107;
    wire N__7104;
    wire N__7099;
    wire N__7096;
    wire N__7093;
    wire N__7090;
    wire N__7087;
    wire N__7084;
    wire N__7083;
    wire N__7078;
    wire N__7075;
    wire N__7074;
    wire N__7073;
    wire N__7070;
    wire N__7069;
    wire N__7066;
    wire N__7063;
    wire N__7060;
    wire N__7057;
    wire N__7052;
    wire N__7049;
    wire N__7046;
    wire N__7045;
    wire N__7044;
    wire N__7041;
    wire N__7036;
    wire N__7033;
    wire N__7030;
    wire N__7021;
    wire N__7018;
    wire N__7017;
    wire N__7016;
    wire N__7013;
    wire N__7010;
    wire N__7007;
    wire N__7004;
    wire N__7003;
    wire N__6998;
    wire N__6997;
    wire N__6994;
    wire N__6991;
    wire N__6988;
    wire N__6985;
    wire N__6976;
    wire N__6973;
    wire N__6970;
    wire N__6967;
    wire N__6964;
    wire N__6961;
    wire N__6958;
    wire N__6955;
    wire N__6954;
    wire N__6953;
    wire N__6950;
    wire N__6945;
    wire N__6940;
    wire N__6939;
    wire N__6938;
    wire N__6935;
    wire N__6934;
    wire N__6933;
    wire N__6932;
    wire N__6929;
    wire N__6928;
    wire N__6927;
    wire N__6924;
    wire N__6923;
    wire N__6922;
    wire N__6921;
    wire N__6916;
    wire N__6913;
    wire N__6912;
    wire N__6911;
    wire N__6904;
    wire N__6901;
    wire N__6900;
    wire N__6895;
    wire N__6894;
    wire N__6891;
    wire N__6888;
    wire N__6887;
    wire N__6886;
    wire N__6885;
    wire N__6882;
    wire N__6879;
    wire N__6876;
    wire N__6873;
    wire N__6868;
    wire N__6865;
    wire N__6864;
    wire N__6861;
    wire N__6854;
    wire N__6851;
    wire N__6850;
    wire N__6849;
    wire N__6846;
    wire N__6843;
    wire N__6838;
    wire N__6835;
    wire N__6832;
    wire N__6829;
    wire N__6826;
    wire N__6823;
    wire N__6818;
    wire N__6813;
    wire N__6806;
    wire N__6803;
    wire N__6798;
    wire N__6793;
    wire N__6784;
    wire N__6779;
    wire N__6776;
    wire N__6773;
    wire N__6768;
    wire N__6765;
    wire N__6762;
    wire N__6757;
    wire N__6754;
    wire N__6753;
    wire N__6752;
    wire N__6749;
    wire N__6746;
    wire N__6745;
    wire N__6744;
    wire N__6741;
    wire N__6738;
    wire N__6735;
    wire N__6728;
    wire N__6725;
    wire N__6722;
    wire N__6719;
    wire N__6716;
    wire N__6713;
    wire N__6710;
    wire N__6707;
    wire N__6702;
    wire N__6699;
    wire N__6696;
    wire N__6691;
    wire N__6688;
    wire N__6685;
    wire N__6684;
    wire N__6679;
    wire N__6676;
    wire N__6673;
    wire N__6672;
    wire N__6669;
    wire N__6666;
    wire N__6661;
    wire N__6658;
    wire N__6655;
    wire N__6652;
    wire N__6649;
    wire N__6646;
    wire N__6643;
    wire N__6640;
    wire N__6637;
    wire N__6634;
    wire N__6631;
    wire N__6628;
    wire N__6625;
    wire N__6624;
    wire N__6621;
    wire N__6618;
    wire N__6617;
    wire N__6614;
    wire N__6611;
    wire N__6608;
    wire N__6601;
    wire N__6600;
    wire N__6595;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6577;
    wire N__6574;
    wire N__6571;
    wire N__6568;
    wire N__6565;
    wire N__6562;
    wire N__6559;
    wire N__6556;
    wire N__6553;
    wire N__6550;
    wire N__6547;
    wire N__6544;
    wire N__6543;
    wire N__6540;
    wire N__6539;
    wire N__6536;
    wire N__6535;
    wire N__6534;
    wire N__6533;
    wire N__6530;
    wire N__6527;
    wire N__6524;
    wire N__6519;
    wire N__6518;
    wire N__6515;
    wire N__6506;
    wire N__6503;
    wire N__6496;
    wire N__6493;
    wire N__6490;
    wire N__6487;
    wire N__6484;
    wire N__6483;
    wire N__6480;
    wire N__6477;
    wire N__6472;
    wire N__6469;
    wire N__6466;
    wire N__6463;
    wire N__6460;
    wire N__6457;
    wire N__6454;
    wire N__6451;
    wire N__6448;
    wire N__6445;
    wire N__6442;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6430;
    wire N__6429;
    wire N__6426;
    wire N__6423;
    wire N__6418;
    wire N__6415;
    wire N__6412;
    wire N__6409;
    wire N__6406;
    wire N__6403;
    wire N__6400;
    wire N__6397;
    wire N__6394;
    wire N__6391;
    wire N__6388;
    wire N__6385;
    wire N__6382;
    wire N__6381;
    wire N__6380;
    wire N__6375;
    wire N__6372;
    wire N__6367;
    wire N__6364;
    wire N__6361;
    wire N__6358;
    wire N__6355;
    wire N__6352;
    wire N__6349;
    wire N__6348;
    wire N__6345;
    wire N__6342;
    wire N__6337;
    wire N__6334;
    wire N__6331;
    wire N__6328;
    wire N__6325;
    wire N__6322;
    wire N__6319;
    wire N__6316;
    wire N__6313;
    wire N__6310;
    wire N__6307;
    wire N__6306;
    wire N__6303;
    wire N__6300;
    wire N__6295;
    wire N__6292;
    wire N__6289;
    wire N__6286;
    wire N__6283;
    wire N__6280;
    wire N__6279;
    wire N__6278;
    wire N__6275;
    wire N__6272;
    wire N__6269;
    wire N__6268;
    wire N__6267;
    wire N__6264;
    wire N__6261;
    wire N__6258;
    wire N__6255;
    wire N__6252;
    wire N__6249;
    wire N__6246;
    wire N__6243;
    wire N__6240;
    wire N__6237;
    wire N__6226;
    wire N__6225;
    wire N__6224;
    wire N__6223;
    wire N__6222;
    wire N__6221;
    wire N__6220;
    wire N__6219;
    wire N__6218;
    wire N__6217;
    wire N__6216;
    wire N__6215;
    wire N__6214;
    wire N__6213;
    wire N__6212;
    wire N__6211;
    wire N__6210;
    wire N__6205;
    wire N__6202;
    wire N__6199;
    wire N__6196;
    wire N__6187;
    wire N__6182;
    wire N__6177;
    wire N__6174;
    wire N__6169;
    wire N__6166;
    wire N__6161;
    wire N__6156;
    wire N__6143;
    wire N__6142;
    wire N__6139;
    wire N__6136;
    wire N__6133;
    wire N__6130;
    wire N__6121;
    wire N__6118;
    wire N__6117;
    wire N__6116;
    wire N__6113;
    wire N__6112;
    wire N__6111;
    wire N__6110;
    wire N__6107;
    wire N__6106;
    wire N__6105;
    wire N__6100;
    wire N__6095;
    wire N__6092;
    wire N__6091;
    wire N__6088;
    wire N__6085;
    wire N__6084;
    wire N__6081;
    wire N__6080;
    wire N__6073;
    wire N__6070;
    wire N__6067;
    wire N__6064;
    wire N__6061;
    wire N__6058;
    wire N__6055;
    wire N__6052;
    wire N__6051;
    wire N__6050;
    wire N__6049;
    wire N__6046;
    wire N__6045;
    wire N__6036;
    wire N__6033;
    wire N__6030;
    wire N__6023;
    wire N__6020;
    wire N__6017;
    wire N__6014;
    wire N__6011;
    wire N__6002;
    wire N__5997;
    wire N__5994;
    wire N__5991;
    wire N__5988;
    wire N__5985;
    wire N__5980;
    wire N__5979;
    wire N__5978;
    wire N__5977;
    wire N__5972;
    wire N__5969;
    wire N__5968;
    wire N__5965;
    wire N__5964;
    wire N__5963;
    wire N__5962;
    wire N__5961;
    wire N__5960;
    wire N__5957;
    wire N__5954;
    wire N__5951;
    wire N__5950;
    wire N__5947;
    wire N__5940;
    wire N__5939;
    wire N__5936;
    wire N__5935;
    wire N__5932;
    wire N__5931;
    wire N__5928;
    wire N__5925;
    wire N__5922;
    wire N__5919;
    wire N__5914;
    wire N__5911;
    wire N__5902;
    wire N__5887;
    wire N__5886;
    wire N__5883;
    wire N__5878;
    wire N__5875;
    wire N__5872;
    wire N__5869;
    wire N__5866;
    wire N__5865;
    wire N__5862;
    wire N__5859;
    wire N__5856;
    wire N__5853;
    wire N__5848;
    wire N__5845;
    wire N__5842;
    wire N__5839;
    wire N__5836;
    wire N__5833;
    wire N__5830;
    wire N__5827;
    wire N__5824;
    wire N__5821;
    wire N__5818;
    wire N__5815;
    wire N__5812;
    wire N__5809;
    wire N__5806;
    wire N__5803;
    wire N__5800;
    wire N__5797;
    wire N__5794;
    wire N__5791;
    wire N__5788;
    wire N__5785;
    wire N__5782;
    wire N__5779;
    wire N__5776;
    wire N__5773;
    wire N__5770;
    wire N__5767;
    wire N__5764;
    wire N__5761;
    wire N__5758;
    wire N__5755;
    wire N__5754;
    wire N__5751;
    wire N__5748;
    wire N__5747;
    wire N__5744;
    wire N__5741;
    wire N__5738;
    wire N__5737;
    wire N__5736;
    wire N__5731;
    wire N__5730;
    wire N__5727;
    wire N__5724;
    wire N__5721;
    wire N__5718;
    wire N__5715;
    wire N__5708;
    wire N__5705;
    wire N__5702;
    wire N__5699;
    wire N__5694;
    wire N__5691;
    wire N__5688;
    wire N__5683;
    wire N__5682;
    wire N__5679;
    wire N__5676;
    wire N__5675;
    wire N__5674;
    wire N__5671;
    wire N__5670;
    wire N__5669;
    wire N__5666;
    wire N__5661;
    wire N__5658;
    wire N__5655;
    wire N__5652;
    wire N__5649;
    wire N__5640;
    wire N__5637;
    wire N__5632;
    wire N__5629;
    wire N__5628;
    wire N__5625;
    wire N__5620;
    wire N__5617;
    wire N__5614;
    wire N__5613;
    wire N__5610;
    wire N__5607;
    wire N__5602;
    wire N__5599;
    wire N__5596;
    wire N__5593;
    wire N__5590;
    wire N__5587;
    wire N__5584;
    wire N__5581;
    wire N__5578;
    wire N__5575;
    wire N__5572;
    wire N__5569;
    wire N__5566;
    wire N__5563;
    wire N__5560;
    wire N__5557;
    wire N__5554;
    wire N__5551;
    wire N__5548;
    wire N__5547;
    wire N__5542;
    wire N__5539;
    wire N__5536;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5518;
    wire N__5515;
    wire N__5514;
    wire N__5511;
    wire N__5508;
    wire N__5505;
    wire N__5502;
    wire N__5497;
    wire N__5494;
    wire N__5493;
    wire N__5492;
    wire N__5489;
    wire N__5486;
    wire N__5483;
    wire N__5476;
    wire N__5473;
    wire N__5470;
    wire N__5467;
    wire N__5464;
    wire N__5461;
    wire N__5458;
    wire N__5455;
    wire N__5452;
    wire N__5449;
    wire N__5446;
    wire N__5443;
    wire N__5440;
    wire N__5437;
    wire N__5434;
    wire N__5431;
    wire N__5428;
    wire N__5425;
    wire N__5422;
    wire N__5419;
    wire N__5416;
    wire N__5413;
    wire N__5410;
    wire N__5407;
    wire N__5404;
    wire N__5401;
    wire N__5398;
    wire N__5395;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5373;
    wire N__5370;
    wire N__5367;
    wire N__5362;
    wire N__5359;
    wire N__5358;
    wire N__5357;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5332;
    wire N__5329;
    wire N__5326;
    wire N__5323;
    wire N__5320;
    wire N__5317;
    wire N__5314;
    wire N__5311;
    wire N__5308;
    wire N__5305;
    wire N__5304;
    wire N__5301;
    wire N__5298;
    wire N__5293;
    wire N__5290;
    wire N__5287;
    wire N__5284;
    wire N__5281;
    wire N__5278;
    wire N__5277;
    wire N__5274;
    wire N__5271;
    wire N__5268;
    wire N__5265;
    wire N__5260;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5248;
    wire N__5245;
    wire N__5242;
    wire N__5239;
    wire N__5236;
    wire N__5233;
    wire N__5232;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5222;
    wire N__5221;
    wire N__5214;
    wire N__5211;
    wire N__5208;
    wire N__5205;
    wire N__5200;
    wire N__5197;
    wire N__5194;
    wire N__5191;
    wire N__5188;
    wire N__5185;
    wire N__5184;
    wire N__5181;
    wire N__5178;
    wire N__5175;
    wire N__5172;
    wire N__5167;
    wire N__5166;
    wire N__5163;
    wire N__5160;
    wire N__5155;
    wire N__5154;
    wire N__5151;
    wire N__5148;
    wire N__5143;
    wire N__5140;
    wire N__5137;
    wire N__5134;
    wire N__5131;
    wire N__5128;
    wire N__5125;
    wire N__5122;
    wire N__5121;
    wire N__5120;
    wire N__5117;
    wire N__5114;
    wire N__5111;
    wire N__5108;
    wire N__5103;
    wire N__5100;
    wire N__5097;
    wire N__5094;
    wire N__5091;
    wire N__5086;
    wire N__5083;
    wire N__5080;
    wire N__5077;
    wire N__5074;
    wire N__5071;
    wire N__5068;
    wire N__5065;
    wire N__5062;
    wire N__5059;
    wire N__5056;
    wire N__5055;
    wire N__5052;
    wire N__5049;
    wire N__5044;
    wire N__5043;
    wire N__5040;
    wire N__5037;
    wire N__5032;
    wire N__5029;
    wire N__5026;
    wire N__5023;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5013;
    wire N__5012;
    wire N__5009;
    wire N__5006;
    wire N__5003;
    wire N__5000;
    wire N__4995;
    wire N__4992;
    wire N__4989;
    wire N__4986;
    wire N__4983;
    wire N__4978;
    wire N__4975;
    wire N__4972;
    wire N__4969;
    wire N__4966;
    wire N__4963;
    wire N__4960;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4950;
    wire N__4947;
    wire N__4944;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4930;
    wire N__4927;
    wire N__4926;
    wire N__4923;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4905;
    wire N__4902;
    wire N__4899;
    wire N__4894;
    wire N__4891;
    wire N__4888;
    wire N__4885;
    wire N__4884;
    wire N__4879;
    wire N__4876;
    wire N__4873;
    wire N__4870;
    wire N__4867;
    wire N__4866;
    wire N__4863;
    wire N__4860;
    wire N__4857;
    wire N__4854;
    wire N__4851;
    wire N__4846;
    wire N__4843;
    wire N__4840;
    wire N__4837;
    wire N__4834;
    wire N__4833;
    wire N__4830;
    wire N__4827;
    wire N__4824;
    wire N__4821;
    wire N__4818;
    wire N__4815;
    wire N__4812;
    wire N__4809;
    wire N__4806;
    wire N__4803;
    wire N__4798;
    wire N__4795;
    wire N__4792;
    wire N__4789;
    wire N__4786;
    wire N__4783;
    wire N__4780;
    wire N__4777;
    wire N__4774;
    wire N__4771;
    wire N__4768;
    wire N__4765;
    wire N__4762;
    wire N__4761;
    wire N__4760;
    wire N__4759;
    wire N__4758;
    wire N__4757;
    wire N__4756;
    wire N__4755;
    wire N__4754;
    wire N__4753;
    wire N__4752;
    wire N__4751;
    wire N__4750;
    wire N__4723;
    wire CLK80_OUT;
    wire PPIO_c;
    wire GNDG0;
    wire SPIO_c;
    wire VCCG0;
    wire A_c_27;
    wire A_c_28;
    wire A_c_26;
    wire \U409_ADDRESS_DECODE.m12Z0Z_5 ;
    wire \U409_ADDRESS_DECODE.m12Z0Z_0_cascade_ ;
    wire \U409_AUTOCONFIG.un1_A_13Z0Z_1 ;
    wire A_c_25;
    wire A_c_24;
    wire \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_3 ;
    wire \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4_cascade_ ;
    wire U409_ADDRESS_DECODE_un1_BPRO_ENn_i;
    wire A_c_29;
    wire \U409_ADDRESS_DECODE.N_26_cascade_ ;
    wire \U409_ADDRESS_DECODE.m54Z0Z_1 ;
    wire \U409_AUTOCONFIG.un1_A_13Z0Z_3 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a4_0_0Z0Z_0 ;
    wire A_c_30;
    wire A_c_31;
    wire \U409_ADDRESS_DECODE.N_59 ;
    wire \U409_ADDRESS_DECODE.N_59_cascade_ ;
    wire \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7 ;
    wire TT_c_1;
    wire TT_c_0;
    wire TM_c_2;
    wire D_1_i;
    wire CONFIGENn_c;
    wire \INVU409_AUTOCONFIG.CONFIGENnC_net ;
    wire PRO_BASE_2;
    wire PRO_BASE_0;
    wire PRO_BASE_1;
    wire \INVU409_AUTOCONFIG.LIDE_CONFC_net ;
    wire \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1_cascade_ ;
    wire \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa ;
    wire \U409_AUTOCONFIG.LIDE_OUT_7_i_a4_0_0 ;
    wire \U409_AUTOCONFIG.N_216_3_cascade_ ;
    wire \U409_AUTOCONFIG.N_108 ;
    wire \U409_AUTOCONFIG.N_108_cascade_ ;
    wire U409_ADDRESS_DECODE_AUTOVECTOR_8;
    wire U409_ADDRESS_DECODE_AUTOVECTOR_9;
    wire U409_ADDRESS_DECODE_AUTOVECTOR_10;
    wire \U409_AUTOCONFIG.N_99 ;
    wire \U409_AUTOCONFIG.N_100 ;
    wire \U409_AUTOCONFIG.LIDE_OUT_RNI9FMPZ0Z_2_cascade_ ;
    wire D_OUT_2;
    wire D_OUT_1;
    wire \INVU409_AUTOCONFIG.LIDE_OUT_0C_net ;
    wire \U409_AUTOCONFIG.N_111 ;
    wire \U409_AUTOCONFIG.N_105_cascade_ ;
    wire \U409_AUTOCONFIG.PR_OUTZ0Z_1 ;
    wire \U409_AUTOCONFIG.N_91 ;
    wire \U409_AUTOCONFIG.N_91_cascade_ ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2 ;
    wire \INVU409_AUTOCONFIG.PR_OUT_1C_net ;
    wire \U409_AUTOCONFIG.N_216_3 ;
    wire \U409_AUTOCONFIG.LIDE_OUT_7_i_0_1_cascade_ ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ;
    wire \U409_AUTOCONFIG.LIDE_OUT_RNI7DMPZ0Z_1 ;
    wire \U409_AUTOCONFIG.N_116 ;
    wire \U409_AUTOCONFIG.N_89 ;
    wire \U409_AUTOCONFIG.PR_OUT_cnst_i_i_0_2_cascade_ ;
    wire \U409_AUTOCONFIG.PR_OUTZ0Z_2 ;
    wire \INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net ;
    wire PORTSIZE_0_i;
    wire A_c_3;
    wire A_c_6;
    wire \U409_AUTOCONFIG.N_109_cascade_ ;
    wire \U409_AUTOCONFIG.N_117 ;
    wire \U409_AUTOCONFIG.N_113 ;
    wire AUTOBOOT_c;
    wire \U409_AUTOCONFIG.N_101 ;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0_cascade_ ;
    wire \U409_AUTOCONFIG.N_119 ;
    wire \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net ;
    wire \U409_AUTOCONFIG.PR_OUTZ0Z_3 ;
    wire \U409_AUTOCONFIG.D_OUT_sm0_0_cascade_ ;
    wire D_OUT_3;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ;
    wire \U409_AUTOCONFIG.LIDE_OUT_RNIBHMPZ0Z_3 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_0 ;
    wire \U409_AUTOCONFIG.PR_OUTZ0Z_0 ;
    wire \U409_AUTOCONFIG.LIDE_OUT_RNI5BMPZ0Z_0_cascade_ ;
    wire \U409_AUTOCONFIG.D_OUT_sm0_0 ;
    wire D_OUT_0;
    wire \U409_AUTOCONFIG.N_90 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ;
    wire \U409_AUTOCONFIG.N_98 ;
    wire CPUCONFn_c;
    wire \U409_AUTOCONFIG.STATE4_cascade_ ;
    wire \U409_AUTOCONFIG.N_104 ;
    wire \U409_AUTOCONFIG.N_103_cascade_ ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ;
    wire \INVU409_AUTOCONFIG.LIDE_OUT_2C_net ;
    wire \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i ;
    wire A_c_4;
    wire A_c_2;
    wire \U409_AUTOCONFIG.N_109 ;
    wire \U409_AUTOCONFIG.N_115 ;
    wire \U409_AUTOCONFIG.AC_STARTZ0 ;
    wire \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_a3_0 ;
    wire \U409_CIA.CLK_CIA_r_1_0_cascade_ ;
    wire bfn_8_12_0_;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_1 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_5 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_6 ;
    wire \U409_CIA.CLK_CIA6_3 ;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0 ;
    wire U409_ADDRESS_DECODE_un1_RTC_ENn_i;
    wire BRIDGE_BASE_2;
    wire \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1 ;
    wire \INVU409_AUTOCONFIG.LIDE_BASE_1C_net ;
    wire \INVU409_AUTOCONFIG.BRIDGE_BASE_0C_net ;
    wire BRIDGE_BASE_0;
    wire \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_4 ;
    wire \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_3 ;
    wire \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_1_cascade_ ;
    wire \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_2 ;
    wire U409_ADDRESS_DECODE_un1_BREG_ENn_i;
    wire \U409_AUTOCONFIG.LIDE_CONFZ0 ;
    wire \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_0 ;
    wire BRIDGE_BASE_4;
    wire BRIDGE_BASE_7;
    wire A_c_7;
    wire A_c_5;
    wire \U409_AUTOCONFIG.un1_STATE_6Z0Z_1 ;
    wire \U409_AUTOCONFIG.un1_STATE_6_0 ;
    wire A_c_1;
    wire \U409_AUTOCONFIG.un1_STATE_6_0_cascade_ ;
    wire D_in_6;
    wire \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1Z0Z_0_cascade_ ;
    wire BRIDGE_BASE_6;
    wire \INVU409_AUTOCONFIG.BRIDGE_BASE_4C_net ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ;
    wire CIA_SPACE;
    wire \U409_CIA.VMA_RNOZ0Z_0_cascade_ ;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENn_2_cascade_ ;
    wire U409_ADDRESS_DECODE_un1_REGSPACEn_i;
    wire \U409_CIA.un1_CIA_CLK_COUNT_3_2 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_2 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_5 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_3 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_4 ;
    wire \U409_CIA.CIA_CLK_COUNT11_3_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNT11 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_0 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_1 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_7 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_6 ;
    wire \U409_CIA.CLK_CIA6_4 ;
    wire \U409_ADDRESS_DECODE.N_77_mux_cascade_ ;
    wire N_22_0_i;
    wire U409_ADDRESS_DECODE_un1_RTC_ENn;
    wire \U409_ADDRESS_DECODE.PORTSIZE_2 ;
    wire A_c_18;
    wire LIDE_BASE_1;
    wire A_c_17;
    wire LIDE_BASE_2;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_0_cascade_ ;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_ ;
    wire CONFIGURED;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3 ;
    wire LIDE_BASE_6;
    wire LIDE_BASE_5;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2 ;
    wire \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1Z0Z_0 ;
    wire BRIDGE_BASE_5;
    wire \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2Z0Z_0 ;
    wire \U409_AUTOCONFIG.un1_AZ0Z_13 ;
    wire \U409_AUTOCONFIG.BRIDGE_CONFZ0 ;
    wire D_in_5;
    wire BRIDGE_BASE_1;
    wire LIDE_BASE_7;
    wire D_in_7;
    wire \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FUZ0Z1 ;
    wire BRIDGE_BASE_3;
    wire \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2Z0Z_1 ;
    wire D_in_4;
    wire un1_AUTOCONFIG_SPACE;
    wire \INVU409_AUTOCONFIG.BRIDGE_BASE_5C_net ;
    wire N_71_mux_cascade_;
    wire N_23_cascade_;
    wire \U409_ADDRESS_DECODE.m33Z0Z_3 ;
    wire \U409_ADDRESS_DECODE.m27Z0Z_3_cascade_ ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ;
    wire U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_4;
    wire U409_ADDRESS_DECODE_m33_1;
    wire U409_ADDRESS_DECODE_m33_1_cascade_;
    wire U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_5;
    wire U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_1;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c2 ;
    wire U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_2;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c2_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ;
    wire N_23;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ;
    wire U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_3;
    wire U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_0;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net ;
    wire \U409_ADDRESS_DECODE.CIA_SPACE_4 ;
    wire \U409_ADDRESS_DECODE.CIA_SPACE_5 ;
    wire LIDE_BASE_4;
    wire LIDE_BASE_3;
    wire \U409_ADDRESS_DECODE.ATA_SPACE_1Z0Z_0 ;
    wire AUTOCONFIG_SPACE;
    wire BUFENn_c;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0 ;
    wire \U409_ADDRESS_DECODE.ATA_ENZ0 ;
    wire U409_ADDRESS_DECODE_un1_ATA_ENn_i;
    wire U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_7;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_EN_nerC_net ;
    wire \U409_AUTOCONFIG.STATE4 ;
    wire \INVU409_AUTOCONFIG.STATE_1C_net ;
    wire U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_6;
    wire N_71_mux;
    wire N_70_mux;
    wire \U409_TRANSFER_ACK.N_20_0 ;
    wire \U409_AUTOCONFIG.STATE_d_2 ;
    wire \U409_AUTOCONFIG.STATEZ0Z_1 ;
    wire RnW_c;
    wire \U409_AUTOCONFIG.STATEZ0Z_0 ;
    wire \INVU409_AUTOCONFIG.AC_TACKC_net ;
    wire U409_ADDRESS_DECODE_un1_REGSPACEn;
    wire TACKn_in;
    wire U409_ADDRESS_DECODE_un1_RAMSPACEn;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ;
    wire GB_BUFFER_CLK40_IN_c_g_THRU_CO;
    wire A_c_16;
    wire A_c_15;
    wire A_c_13;
    wire U409_ADDRESS_DECODE_un1_CIACS1n_i;
    wire CIA_ENABLE;
    wire CIA_ENABLE_cascade_;
    wire A_c_12;
    wire U409_ADDRESS_DECODE_un1_CIACS0n_i;
    wire \U409_ADDRESS_DECODE.N_75 ;
    wire N_77_mux_i;
    wire \U409_ADDRESS_DECODE.N_60_1 ;
    wire U409_ADDRESS_DECODE_un1_RAMSPACEn_i;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ;
    wire AC_TACK;
    wire \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_ ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ;
    wire \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ;
    wire TACK_OUTn;
    wire \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER6 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net ;
    wire \U409_ADDRESS_DECODE.Z2_SPACE ;
    wire ROMEN_cascade_;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0_cascade_ ;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENn_2 ;
    wire \U409_ADDRESS_DECODE.N_61 ;
    wire \U409_TRANSFER_ACK.N_42_i_cascade_ ;
    wire A_c_23;
    wire A_c_20;
    wire \U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_1 ;
    wire A_c_19;
    wire A_c_22;
    wire OVL_c;
    wire A_c_21;
    wire \U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_2 ;
    wire ROMEN;
    wire TACK_EN;
    wire TCIn_1_i;
    wire RESETn_c_i;
    wire \U409_TRANSFER_ACK.un1_AUTOVECTOR_0 ;
    wire TSn_c;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1_cascade_ ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER22_NE_1_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_NE_1_0_cascade_ ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0_0 ;
    wire ROMENn_c;
    wire \INVU409_TRANSFER_ACK.ROMENnC_net ;
    wire \U409_TRANSFER_ACK.N_42_i ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER21_0 ;
    wire PCIAT_c_1;
    wire TM_c_0;
    wire \U409_ADDRESS_DECODE.N_58_mux ;
    wire TM_c_1;
    wire PCIAT_c_0;
    wire bfn_14_6_0_;
    wire \U409_TICK.un3_COUNTER60_1_cry_1 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_2 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_3 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_4 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_6 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_8 ;
    wire bfn_14_7_0_;
    wire \U409_TICK.un3_COUNTER60_1_cry_9 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_10 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_13 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_15 ;
    wire \U409_TRANSFER_ACK.CIA_TACK_ENZ0 ;
    wire \U409_CIA.VMAZ0 ;
    wire \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.N_33 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER21_NE_0_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER22_NE_0_0 ;
    wire ROM_DELAY_c_0;
    wire ROM_DELAY_c_1;
    wire \U409_TRANSFER_ACK.N_31_i ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_9 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_8 ;
    wire \U409_TICK.COUNTER60Z0Z_5 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_4 ;
    wire \U409_TICK.COUNTER60Z0Z_4 ;
    wire \U409_TICK.COUNTER60Z0Z_9 ;
    wire \U409_TICK.COUNTER60Z0Z_8 ;
    wire \U409_TICK.TICK603_9_cascade_ ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_6 ;
    wire \U409_TICK.COUNTER60Z0Z_6 ;
    wire \U409_TICK.COUNTER60Z0Z_13 ;
    wire \U409_TICK.COUNTER60Z0Z_10 ;
    wire \U409_TICK.COUNTER60Z0Z_7 ;
    wire \U409_TICK.TICK603_10_cascade_ ;
    wire \U409_TICK.COUNTER60Z0Z_0 ;
    wire \U409_TICK.COUNTER60Z0Z_12 ;
    wire \U409_TICK.COUNTER60Z0Z_2 ;
    wire \U409_TICK.COUNTER60Z0Z_1 ;
    wire \U409_TICK.COUNTER60Z0Z_16 ;
    wire \U409_TICK.TICK603_8 ;
    wire \U409_TICK.COUNTER60Z0Z_11 ;
    wire \U409_TICK.TICK603_11_cascade_ ;
    wire \U409_TICK.COUNTER60Z0Z_3 ;
    wire \U409_TICK.TICK603_14_cascade_ ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_14 ;
    wire \U409_TICK.COUNTER60Z0Z_14 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER60Z0Z_15 ;
    wire \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_ ;
    wire CLK40_IN_c_g;
    wire \U409_TRANSFER_ACK.N_17_mux ;
    wire \U409_TRANSFER_ACK.N_3_0_cascade_ ;
    wire \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ;
    wire \U409_TRANSFER_ACK.N_3_0 ;
    wire RESETn_c;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ;
    wire \U409_TRANSFER_ACK.N_55_cascade_ ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_0C_net ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_1 ;
    wire CLK_CIA_c;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_0 ;
    wire \INVU409_TRANSFER_ACK.LASTCLK_1C_net ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0 ;
    wire N_52_1;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ;
    wire RESETn_c_i_g;
    wire \U409_TICK.TICK503_10_cascade_ ;
    wire \U409_TICK.TICK603_10 ;
    wire \U409_TICK.TICK603_9 ;
    wire \U409_TICK.TICK603_14 ;
    wire TICK60_c;
    wire CONSTANT_ONE_NET;
    wire \U409_TICK.TICK503_8 ;
    wire \U409_TICK.TICK503_11_cascade_ ;
    wire \U409_TICK.TICK503_14_cascade_ ;
    wire TICK50_c;
    wire \U409_TICK.TICK503_9_cascade_ ;
    wire \U409_TICK.COUNTER50Z0Z_1 ;
    wire \U409_TICK.COUNTER50Z0Z_0 ;
    wire bfn_17_5_0_;
    wire \U409_TICK.COUNTER50Z0Z_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_1 ;
    wire \U409_TICK.COUNTER50Z0Z_3 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_2 ;
    wire \U409_TICK.COUNTER50Z0Z_4 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_3 ;
    wire \U409_TICK.COUNTER50Z0Z_5 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_4 ;
    wire \U409_TICK.COUNTER50Z0Z_6 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_6 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_5 ;
    wire \U409_TICK.COUNTER50Z0Z_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_6 ;
    wire \U409_TICK.COUNTER50Z0Z_8 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_8 ;
    wire \U409_TICK.COUNTER50Z0Z_9 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_9 ;
    wire bfn_17_6_0_;
    wire \U409_TICK.COUNTER50Z0Z_10 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_9 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_10 ;
    wire \U409_TICK.COUNTER50Z0Z_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_11 ;
    wire \U409_TICK.COUNTER50Z0Z_13 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_13 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_12 ;
    wire \U409_TICK.COUNTER50Z0Z_14 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_13 ;
    wire \U409_TICK.COUNTER50Z0Z_15 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_15 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_15 ;
    wire \U409_TICK.COUNTER50Z0Z_16 ;
    wire \U409_TICK.TICK503_14 ;
    wire \U409_TICK.TICK503_9 ;
    wire \U409_TICK.TICK503_10 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_11 ;
    wire \U409_TICK.COUNTER50Z0Z_11 ;
    wire CLK6_c_g;
    wire PCS0_c;
    wire SCS1_c;
    wire \U409_ADDRESS_DECODE.CSZ0Z0 ;
    wire PCS1_c;
    wire \U409_ADDRESS_DECODE.CSZ0Z1 ;
    wire A_c_14;
    wire SCS0_c;
    wire XCLK_ENn_c;
    wire XCLK_c;
    wire CLK28_IN_c_g;
    wire AGNUS_CLK_c;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="SIMPLE";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0001111;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE pll (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__8638),
            .RESETB(N__11981),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(CLK80_OUT));
    PRE_IO_GBUF CLK40_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__13651),
            .GLOBALBUFFEROUTPUT(CLK40_IN_c_g));
    IO_PAD CLK40_IN_ibuf_gb_io_iopad (
            .OE(N__13653),
            .DIN(N__13652),
            .DOUT(N__13651),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_gb_io_preio (
            .PADOEN(N__13653),
            .PADOUT(N__13652),
            .PADIN(N__13651),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK28_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__13641),
            .GLOBALBUFFEROUTPUT(CLK28_IN_c_g));
    IO_PAD CLK28_IN_ibuf_gb_io_iopad (
            .OE(N__13643),
            .DIN(N__13642),
            .DOUT(N__13641),
            .PACKAGEPIN(CLK28_IN));
    defparam CLK28_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK28_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK28_IN_ibuf_gb_io_preio (
            .PADOEN(N__13643),
            .PADOUT(N__13642),
            .PADIN(N__13641),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK6_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__13631),
            .GLOBALBUFFEROUTPUT(CLK6_c_g));
    IO_PAD CLK6_ibuf_gb_io_iopad (
            .OE(N__13633),
            .DIN(N__13632),
            .DOUT(N__13631),
            .PACKAGEPIN(CLK6));
    defparam CLK6_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK6_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK6_ibuf_gb_io_preio (
            .PADOEN(N__13633),
            .PADOUT(N__13632),
            .PADIN(N__13631),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__13622),
            .DIN(N__13621),
            .DOUT(N__13620),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__13622),
            .PADOUT(N__13621),
            .PADIN(N__13620),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_0_iopad (
            .OE(N__13613),
            .DIN(N__13612),
            .DOUT(N__13611),
            .PACKAGEPIN(TT[0]));
    defparam TT_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_0_preio (
            .PADOEN(N__13613),
            .PADOUT(N__13612),
            .PADIN(N__13611),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ROM_DELAY_ibuf_1_iopad.PULLUP=1'b1;
    IO_PAD ROM_DELAY_ibuf_1_iopad (
            .OE(N__13604),
            .DIN(N__13603),
            .DOUT(N__13602),
            .PACKAGEPIN(ROM_DELAY[1]));
    defparam ROM_DELAY_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam ROM_DELAY_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ROM_DELAY_ibuf_1_preio (
            .PADOEN(N__13604),
            .PADOUT(N__13603),
            .PADIN(N__13602),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ROM_DELAY_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_7_iopad (
            .OE(N__13595),
            .DIN(N__13594),
            .DOUT(N__13593),
            .PACKAGEPIN(D[7]));
    defparam D_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_7_preio (
            .PADOEN(N__13595),
            .PADOUT(N__13594),
            .PADIN(N__13593),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5236),
            .DIN0(D_in_7),
            .DOUT0(N__5836),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__13586),
            .DIN(N__13585),
            .DOUT(N__13584),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__13586),
            .PADOUT(N__13585),
            .PADIN(N__13584),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CPUCONFn_ibuf_iopad (
            .OE(N__13577),
            .DIN(N__13576),
            .DOUT(N__13575),
            .PACKAGEPIN(CPUCONFn));
    defparam CPUCONFn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CPUCONFn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CPUCONFn_ibuf_preio (
            .PADOEN(N__13577),
            .PADOUT(N__13576),
            .PADIN(N__13575),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CPUCONFn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RTC_ENn_obuf_iopad (
            .OE(N__13568),
            .DIN(N__13567),
            .DOUT(N__13566),
            .PACKAGEPIN(RTC_ENn));
    defparam RTC_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RTC_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RTC_ENn_obuf_preio (
            .PADOEN(N__13568),
            .PADOUT(N__13567),
            .PADIN(N__13566),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6454),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_24_iopad (
            .OE(N__13559),
            .DIN(N__13558),
            .DOUT(N__13557),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__13559),
            .PADOUT(N__13558),
            .PADIN(N__13557),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SPIO_J_ibuf_iopad.PULLUP=1'b1;
    IO_PAD SPIO_J_ibuf_iopad (
            .OE(N__13550),
            .DIN(N__13549),
            .DOUT(N__13548),
            .PACKAGEPIN(SPIO_J));
    defparam SPIO_J_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam SPIO_J_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO SPIO_J_ibuf_preio (
            .PADOEN(N__13550),
            .PADOUT(N__13549),
            .PADIN(N__13548),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SPIO_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_4_iopad (
            .OE(N__13541),
            .DIN(N__13540),
            .DOUT(N__13539),
            .PACKAGEPIN(D[4]));
    defparam D_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_4_preio (
            .PADOEN(N__13541),
            .PADOUT(N__13540),
            .PADIN(N__13539),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5221),
            .DIN0(D_in_4),
            .DOUT0(N__6367),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PPIO_obuf_iopad (
            .OE(N__13532),
            .DIN(N__13531),
            .DOUT(N__13530),
            .PACKAGEPIN(PPIO));
    defparam PPIO_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PPIO_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PPIO_obuf_preio (
            .PADOEN(N__13532),
            .PADOUT(N__13531),
            .PADIN(N__13530),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4798),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__13523),
            .DIN(N__13522),
            .DOUT(N__13521),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__13523),
            .PADOUT(N__13522),
            .PADIN(N__13521),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TM_ibuf_1_iopad (
            .OE(N__13514),
            .DIN(N__13513),
            .DOUT(N__13512),
            .PACKAGEPIN(TM[1]));
    defparam TM_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TM_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TM_ibuf_1_preio (
            .PADOEN(N__13514),
            .PADOUT(N__13513),
            .PADIN(N__13512),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TM_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_21_iopad (
            .OE(N__13505),
            .DIN(N__13504),
            .DOUT(N__13503),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__13505),
            .PADOUT(N__13504),
            .PADIN(N__13503),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam PPIO_J_ibuf_iopad.PULLUP=1'b1;
    IO_PAD PPIO_J_ibuf_iopad (
            .OE(N__13496),
            .DIN(N__13495),
            .DOUT(N__13494),
            .PACKAGEPIN(PPIO_J));
    defparam PPIO_J_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam PPIO_J_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO PPIO_J_ibuf_preio (
            .PADOEN(N__13496),
            .PADOUT(N__13495),
            .PADIN(N__13494),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(PPIO_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_obuf_iopad (
            .OE(N__13487),
            .DIN(N__13486),
            .DOUT(N__13485),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMSPACEn_obuf_preio (
            .PADOEN(N__13487),
            .PADOUT(N__13486),
            .PADIN(N__13485),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9001),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__13478),
            .DIN(N__13477),
            .DOUT(N__13476),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__13478),
            .PADOUT(N__13477),
            .PADIN(N__13476),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ROMENn_obuf_iopad (
            .OE(N__13469),
            .DIN(N__13468),
            .DOUT(N__13467),
            .PACKAGEPIN(ROMENn));
    defparam ROMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ROMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ROMENn_obuf_preio (
            .PADOEN(N__13469),
            .PADOUT(N__13468),
            .PADIN(N__13467),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10291),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuft_iopad (
            .OE(N__13460),
            .DIN(N__13459),
            .DOUT(N__13458),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TBIn_obuft_preio (
            .PADOEN(N__13460),
            .PADOUT(N__13459),
            .PADIN(N__13458),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9607),
            .DIN0(),
            .DOUT0(N__9498),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam AUTOBOOT_ibuf_iopad.PULLUP=1'b1;
    IO_PAD AUTOBOOT_ibuf_iopad (
            .OE(N__13451),
            .DIN(N__13450),
            .DOUT(N__13449),
            .PACKAGEPIN(AUTOBOOT));
    defparam AUTOBOOT_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AUTOBOOT_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AUTOBOOT_ibuf_preio (
            .PADOEN(N__13451),
            .PADOUT(N__13450),
            .PADIN(N__13449),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AUTOBOOT_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD F_READn_obuf_iopad (
            .OE(N__13442),
            .DIN(N__13441),
            .DOUT(N__13440),
            .PACKAGEPIN(F_READn));
    defparam F_READn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam F_READn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO F_READn_obuf_preio (
            .PADOEN(N__13442),
            .PADOUT(N__13441),
            .PADIN(N__13440),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12001),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__13433),
            .DIN(N__13432),
            .DOUT(N__13431),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__13433),
            .PADOUT(N__13432),
            .PADIN(N__13431),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORTSIZE_obuf_iopad (
            .OE(N__13424),
            .DIN(N__13423),
            .DOUT(N__13422),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PORTSIZE_obuf_preio (
            .PADOEN(N__13424),
            .PADOUT(N__13423),
            .PADIN(N__13422),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5776),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD F_ENn_obuf_iopad (
            .OE(N__13415),
            .DIN(N__13414),
            .DOUT(N__13413),
            .PACKAGEPIN(F_ENn));
    defparam F_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam F_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO F_ENn_obuf_preio (
            .PADOEN(N__13415),
            .PADOUT(N__13414),
            .PADIN(N__13413),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12000),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__13406),
            .DIN(N__13405),
            .DOUT(N__13404),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__13406),
            .PADOUT(N__13405),
            .PADIN(N__13404),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TM_ibuf_2_iopad (
            .OE(N__13397),
            .DIN(N__13396),
            .DOUT(N__13395),
            .PACKAGEPIN(TM[2]));
    defparam TM_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam TM_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO TM_ibuf_2_preio (
            .PADOEN(N__13397),
            .PADOUT(N__13396),
            .PADIN(N__13395),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TM_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_22_iopad (
            .OE(N__13388),
            .DIN(N__13387),
            .DOUT(N__13386),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__13388),
            .PADOUT(N__13387),
            .PADIN(N__13386),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__13379),
            .DIN(N__13378),
            .DOUT(N__13377),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__13379),
            .PADOUT(N__13378),
            .PADIN(N__13377),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__13370),
            .DIN(N__13369),
            .DOUT(N__13368),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__13370),
            .PADOUT(N__13369),
            .PADIN(N__13368),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__13361),
            .DIN(N__13360),
            .DOUT(N__13359),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__13361),
            .PADOUT(N__13360),
            .PADIN(N__13359),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ROM_DELAY_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD ROM_DELAY_ibuf_0_iopad (
            .OE(N__13352),
            .DIN(N__13351),
            .DOUT(N__13350),
            .PACKAGEPIN(ROM_DELAY[0]));
    defparam ROM_DELAY_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam ROM_DELAY_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO ROM_DELAY_ibuf_0_preio (
            .PADOEN(N__13352),
            .PADOUT(N__13351),
            .PADIN(N__13350),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ROM_DELAY_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SCS1_obuf_iopad (
            .OE(N__13343),
            .DIN(N__13342),
            .DOUT(N__13341),
            .PACKAGEPIN(SCS1));
    defparam SCS1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SCS1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SCS1_obuf_preio (
            .PADOEN(N__13343),
            .PADOUT(N__13342),
            .PADIN(N__13341),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12553),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_CLK_obuf_iopad (
            .OE(N__13334),
            .DIN(N__13333),
            .DOUT(N__13332),
            .PACKAGEPIN(AGNUS_CLK));
    defparam AGNUS_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO AGNUS_CLK_obuf_preio (
            .PADOEN(N__13334),
            .PADOUT(N__13333),
            .PADIN(N__13332),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12823),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_25_iopad (
            .OE(N__13325),
            .DIN(N__13324),
            .DOUT(N__13323),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__13325),
            .PADOUT(N__13324),
            .PADIN(N__13323),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS0n_obuf_iopad (
            .OE(N__13316),
            .DIN(N__13315),
            .DOUT(N__13314),
            .PACKAGEPIN(CIACS0n));
    defparam CIACS0n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS0n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS0n_obuf_preio (
            .PADOEN(N__13316),
            .PADOUT(N__13315),
            .PADIN(N__13314),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9124),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK50_obuf_iopad (
            .OE(N__13307),
            .DIN(N__13306),
            .DOUT(N__13305),
            .PACKAGEPIN(TICK50));
    defparam TICK50_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK50_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK50_obuf_preio (
            .PADOEN(N__13307),
            .PADOUT(N__13306),
            .PADIN(N__13305),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12277),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_28_iopad (
            .OE(N__13298),
            .DIN(N__13297),
            .DOUT(N__13296),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__13298),
            .PADOUT(N__13297),
            .PADIN(N__13296),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BREG_ENn_obuf_iopad (
            .OE(N__13289),
            .DIN(N__13288),
            .DOUT(N__13287),
            .PACKAGEPIN(BREG_ENn));
    defparam BREG_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BREG_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BREG_ENn_obuf_preio (
            .PADOEN(N__13289),
            .PADOUT(N__13288),
            .PADIN(N__13287),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6565),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_5_iopad (
            .OE(N__13280),
            .DIN(N__13279),
            .DOUT(N__13278),
            .PACKAGEPIN(D[5]));
    defparam D_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_5_preio (
            .PADOEN(N__13280),
            .PADOUT(N__13279),
            .PADIN(N__13278),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5231),
            .DIN0(D_in_5),
            .DOUT0(N__5404),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD F_BANK_obuf_0_iopad (
            .OE(N__13271),
            .DIN(N__13270),
            .DOUT(N__13269),
            .PACKAGEPIN(F_BANK[0]));
    defparam F_BANK_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam F_BANK_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO F_BANK_obuf_0_preio (
            .PADOEN(N__13271),
            .PADOUT(N__13270),
            .PADIN(N__13269),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7144),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD XCLK_ENn_ibuf_iopad (
            .OE(N__13262),
            .DIN(N__13261),
            .DOUT(N__13260),
            .PACKAGEPIN(XCLK_ENn));
    defparam XCLK_ENn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam XCLK_ENn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO XCLK_ENn_ibuf_preio (
            .PADOEN(N__13262),
            .PADOUT(N__13261),
            .PADIN(N__13260),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(XCLK_ENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__13253),
            .DIN(N__13252),
            .DOUT(N__13251),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__13253),
            .PADOUT(N__13252),
            .PADIN(N__13251),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK60_obuf_iopad (
            .OE(N__13244),
            .DIN(N__13243),
            .DOUT(N__13242),
            .PACKAGEPIN(TICK60));
    defparam TICK60_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK60_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK60_obuf_preio (
            .PADOEN(N__13244),
            .PADOUT(N__13243),
            .PADIN(N__13242),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12025),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_26_iopad (
            .OE(N__13235),
            .DIN(N__13234),
            .DOUT(N__13233),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__13235),
            .PADOUT(N__13234),
            .PADIN(N__13233),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_23_iopad (
            .OE(N__13226),
            .DIN(N__13225),
            .DOUT(N__13224),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__13226),
            .PADOUT(N__13225),
            .PADIN(N__13224),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__13217),
            .DIN(N__13216),
            .DOUT(N__13215),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__13217),
            .PADOUT(N__13216),
            .PADIN(N__13215),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ATA_ENn_obuf_iopad (
            .OE(N__13208),
            .DIN(N__13207),
            .DOUT(N__13206),
            .PACKAGEPIN(ATA_ENn));
    defparam ATA_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ATA_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ATA_ENn_obuf_preio (
            .PADOEN(N__13208),
            .PADOUT(N__13207),
            .PADIN(N__13206),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8329),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_31_iopad (
            .OE(N__13199),
            .DIN(N__13198),
            .DOUT(N__13197),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__13199),
            .PADOUT(N__13198),
            .PADIN(N__13197),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS1n_obuf_iopad (
            .OE(N__13190),
            .DIN(N__13189),
            .DOUT(N__13188),
            .PACKAGEPIN(CIACS1n));
    defparam CIACS1n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS1n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS1n_obuf_preio (
            .PADOEN(N__13190),
            .PADOUT(N__13189),
            .PADIN(N__13188),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9181),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_obuf_iopad (
            .OE(N__13181),
            .DIN(N__13180),
            .DOUT(N__13179),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGSPACEn_obuf_preio (
            .PADOEN(N__13181),
            .PADOUT(N__13180),
            .PADIN(N__13179),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6652),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PCS0_obuf_iopad (
            .OE(N__13172),
            .DIN(N__13171),
            .DOUT(N__13170),
            .PACKAGEPIN(PCS0));
    defparam PCS0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PCS0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PCS0_obuf_preio (
            .PADOEN(N__13172),
            .PADOUT(N__13171),
            .PADIN(N__13170),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12571),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PCIAT_obuf_0_iopad (
            .OE(N__13163),
            .DIN(N__13162),
            .DOUT(N__13161),
            .PACKAGEPIN(PCIAT[0]));
    defparam PCIAT_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam PCIAT_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO PCIAT_obuf_0_preio (
            .PADOEN(N__13163),
            .PADOUT(N__13162),
            .PADIN(N__13161),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10465),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__13154),
            .DIN(N__13153),
            .DOUT(N__13152),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__13154),
            .PADOUT(N__13153),
            .PADIN(N__13152),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_CIA_obuf_iopad (
            .OE(N__13145),
            .DIN(N__13144),
            .DOUT(N__13143),
            .PACKAGEPIN(CLK_CIA));
    defparam CLK_CIA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_CIA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_CIA_obuf_preio (
            .PADOEN(N__13145),
            .PADOUT(N__13144),
            .PADIN(N__13143),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11593),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__13136),
            .DIN(N__13135),
            .DOUT(N__13134),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__13136),
            .PADOUT(N__13135),
            .PADIN(N__13134),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PCS1_obuf_iopad (
            .OE(N__13127),
            .DIN(N__13126),
            .DOUT(N__13125),
            .PACKAGEPIN(PCS1));
    defparam PCS1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PCS1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PCS1_obuf_preio (
            .PADOEN(N__13127),
            .PADOUT(N__13126),
            .PADIN(N__13125),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12505),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__13118),
            .DIN(N__13117),
            .DOUT(N__13116),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__13118),
            .PADOUT(N__13117),
            .PADIN(N__13116),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9603),
            .DIN0(TACKn_in),
            .DOUT0(N__9491),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_1_iopad (
            .OE(N__13109),
            .DIN(N__13108),
            .DOUT(N__13107),
            .PACKAGEPIN(TT[1]));
    defparam TT_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_1_preio (
            .PADOEN(N__13109),
            .PADOUT(N__13108),
            .PADIN(N__13107),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__13100),
            .DIN(N__13099),
            .DOUT(N__13098),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__13100),
            .PADOUT(N__13099),
            .PADIN(N__13098),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8377),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_29_iopad (
            .OE(N__13091),
            .DIN(N__13090),
            .DOUT(N__13089),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__13091),
            .PADOUT(N__13090),
            .PADIN(N__13089),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_6_iopad (
            .OE(N__13082),
            .DIN(N__13081),
            .DOUT(N__13080),
            .PACKAGEPIN(D[6]));
    defparam D_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_6_preio (
            .PADOEN(N__13082),
            .PADOUT(N__13081),
            .PADIN(N__13080),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5232),
            .DIN0(D_in_6),
            .DOUT0(N__5422),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD F_BANK_obuf_1_iopad (
            .OE(N__13073),
            .DIN(N__13072),
            .DOUT(N__13071),
            .PACKAGEPIN(F_BANK[1]));
    defparam F_BANK_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam F_BANK_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO F_BANK_obuf_1_preio (
            .PADOEN(N__13073),
            .PADOUT(N__13072),
            .PADIN(N__13071),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9049),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD F_WRITEn_obuf_iopad (
            .OE(N__13064),
            .DIN(N__13063),
            .DOUT(N__13062),
            .PACKAGEPIN(F_WRITEn));
    defparam F_WRITEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam F_WRITEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO F_WRITEn_obuf_preio (
            .PADOEN(N__13064),
            .PADOUT(N__13063),
            .PADIN(N__13062),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11977),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__13055),
            .DIN(N__13054),
            .DOUT(N__13053),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__13055),
            .PADOUT(N__13054),
            .PADIN(N__13053),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_27_iopad (
            .OE(N__13046),
            .DIN(N__13045),
            .DOUT(N__13044),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__13046),
            .PADOUT(N__13045),
            .PADIN(N__13044),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SCS0_obuf_iopad (
            .OE(N__13037),
            .DIN(N__13036),
            .DOUT(N__13035),
            .PACKAGEPIN(SCS0));
    defparam SCS0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SCS0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SCS0_obuf_preio (
            .PADOEN(N__13037),
            .PADOUT(N__13036),
            .PADIN(N__13035),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12433),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BPRO_ENn_obuf_iopad (
            .OE(N__13028),
            .DIN(N__13027),
            .DOUT(N__13026),
            .PACKAGEPIN(BPRO_ENn));
    defparam BPRO_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BPRO_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BPRO_ENn_obuf_preio (
            .PADOEN(N__13028),
            .PADOUT(N__13027),
            .PADIN(N__13026),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5143),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TM_ibuf_0_iopad (
            .OE(N__13019),
            .DIN(N__13018),
            .DOUT(N__13017),
            .PACKAGEPIN(TM[0]));
    defparam TM_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TM_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TM_ibuf_0_preio (
            .PADOEN(N__13019),
            .PADOUT(N__13018),
            .PADIN(N__13017),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TM_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD XCLK_ibuf_iopad (
            .OE(N__13010),
            .DIN(N__13009),
            .DOUT(N__13008),
            .PACKAGEPIN(XCLK));
    defparam XCLK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam XCLK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO XCLK_ibuf_preio (
            .PADOEN(N__13010),
            .PADOUT(N__13009),
            .PADIN(N__13008),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(XCLK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__13001),
            .DIN(N__13000),
            .DOUT(N__12999),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__13001),
            .PADOUT(N__13000),
            .PADIN(N__12999),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD F_WPn_obuf_iopad (
            .OE(N__12992),
            .DIN(N__12991),
            .DOUT(N__12990),
            .PACKAGEPIN(F_WPn));
    defparam F_WPn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam F_WPn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO F_WPn_obuf_preio (
            .PADOEN(N__12992),
            .PADOUT(N__12991),
            .PADIN(N__12990),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__12983),
            .DIN(N__12982),
            .DOUT(N__12981),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__12983),
            .PADOUT(N__12982),
            .PADIN(N__12981),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__12974),
            .DIN(N__12973),
            .DOUT(N__12972),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__12974),
            .PADOUT(N__12973),
            .PADIN(N__12972),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_30_iopad (
            .OE(N__12965),
            .DIN(N__12964),
            .DOUT(N__12963),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__12965),
            .PADOUT(N__12964),
            .PADIN(N__12963),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD OVL_ibuf_iopad (
            .OE(N__12956),
            .DIN(N__12955),
            .DOUT(N__12954),
            .PACKAGEPIN(OVL));
    defparam OVL_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam OVL_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO OVL_ibuf_preio (
            .PADOEN(N__12956),
            .PADOUT(N__12955),
            .PADIN(N__12954),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(OVL_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuft_iopad (
            .OE(N__12947),
            .DIN(N__12946),
            .DOUT(N__12945),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TCIn_obuft_preio (
            .PADOEN(N__12947),
            .PADOUT(N__12946),
            .PADIN(N__12945),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9559),
            .DIN0(),
            .DOUT0(N__9499),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PCIAT_obuf_1_iopad (
            .OE(N__12938),
            .DIN(N__12937),
            .DOUT(N__12936),
            .PACKAGEPIN(PCIAT[1]));
    defparam PCIAT_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam PCIAT_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO PCIAT_obuf_1_preio (
            .PADOEN(N__12938),
            .PADOUT(N__12937),
            .PADIN(N__12936),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10555),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__12929),
            .DIN(N__12928),
            .DOUT(N__12927),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__12929),
            .PADOUT(N__12928),
            .PADIN(N__12927),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__12920),
            .DIN(N__12919),
            .DOUT(N__12918),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__12920),
            .PADOUT(N__12919),
            .PADIN(N__12918),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CONFIGENn_obuf_iopad (
            .OE(N__12911),
            .DIN(N__12910),
            .DOUT(N__12909),
            .PACKAGEPIN(CONFIGENn));
    defparam CONFIGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CONFIGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CONFIGENn_obuf_preio (
            .PADOEN(N__12911),
            .PADOUT(N__12910),
            .PADIN(N__12909),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5194),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SPIO_obuf_iopad (
            .OE(N__12902),
            .DIN(N__12901),
            .DOUT(N__12900),
            .PACKAGEPIN(SPIO));
    defparam SPIO_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SPIO_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SPIO_obuf_preio (
            .PADOEN(N__12902),
            .PADOUT(N__12901),
            .PADIN(N__12900),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4777),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD F_RSTn_obuf_iopad (
            .OE(N__12893),
            .DIN(N__12892),
            .DOUT(N__12891),
            .PACKAGEPIN(F_RSTn));
    defparam F_RSTn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam F_RSTn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO F_RSTn_obuf_preio (
            .PADOEN(N__12893),
            .PADOUT(N__12892),
            .PADIN(N__12891),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11993),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__3133 (
            .O(N__12874),
            .I(N__12871));
    LocalMux I__3132 (
            .O(N__12871),
            .I(N__12868));
    Span12Mux_v I__3131 (
            .O(N__12868),
            .I(N__12865));
    Odrv12 I__3130 (
            .O(N__12865),
            .I(XCLK_ENn_c));
    InMux I__3129 (
            .O(N__12862),
            .I(N__12859));
    LocalMux I__3128 (
            .O(N__12859),
            .I(N__12856));
    Span4Mux_v I__3127 (
            .O(N__12856),
            .I(N__12853));
    Odrv4 I__3126 (
            .O(N__12853),
            .I(XCLK_c));
    InMux I__3125 (
            .O(N__12850),
            .I(N__12847));
    LocalMux I__3124 (
            .O(N__12847),
            .I(N__12840));
    ClkMux I__3123 (
            .O(N__12846),
            .I(N__12829));
    ClkMux I__3122 (
            .O(N__12845),
            .I(N__12829));
    ClkMux I__3121 (
            .O(N__12844),
            .I(N__12829));
    ClkMux I__3120 (
            .O(N__12843),
            .I(N__12829));
    Glb2LocalMux I__3119 (
            .O(N__12840),
            .I(N__12829));
    GlobalMux I__3118 (
            .O(N__12829),
            .I(N__12826));
    gio2CtrlBuf I__3117 (
            .O(N__12826),
            .I(CLK28_IN_c_g));
    IoInMux I__3116 (
            .O(N__12823),
            .I(N__12820));
    LocalMux I__3115 (
            .O(N__12820),
            .I(N__12817));
    Span4Mux_s3_h I__3114 (
            .O(N__12817),
            .I(N__12814));
    Odrv4 I__3113 (
            .O(N__12814),
            .I(AGNUS_CLK_c));
    InMux I__3112 (
            .O(N__12811),
            .I(N__12807));
    InMux I__3111 (
            .O(N__12810),
            .I(N__12804));
    LocalMux I__3110 (
            .O(N__12807),
            .I(N__12801));
    LocalMux I__3109 (
            .O(N__12804),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    Odrv4 I__3108 (
            .O(N__12801),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    InMux I__3107 (
            .O(N__12796),
            .I(N__12793));
    LocalMux I__3106 (
            .O(N__12793),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ));
    InMux I__3105 (
            .O(N__12790),
            .I(\U409_TICK.un2_COUNTER50_1_cry_13 ));
    InMux I__3104 (
            .O(N__12787),
            .I(N__12783));
    InMux I__3103 (
            .O(N__12786),
            .I(N__12780));
    LocalMux I__3102 (
            .O(N__12783),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    LocalMux I__3101 (
            .O(N__12780),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    CascadeMux I__3100 (
            .O(N__12775),
            .I(N__12772));
    InMux I__3099 (
            .O(N__12772),
            .I(N__12769));
    LocalMux I__3098 (
            .O(N__12769),
            .I(N__12766));
    Odrv4 I__3097 (
            .O(N__12766),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ));
    InMux I__3096 (
            .O(N__12763),
            .I(\U409_TICK.un2_COUNTER50_1_cry_14 ));
    InMux I__3095 (
            .O(N__12760),
            .I(\U409_TICK.un2_COUNTER50_1_cry_15 ));
    InMux I__3094 (
            .O(N__12757),
            .I(N__12753));
    InMux I__3093 (
            .O(N__12756),
            .I(N__12750));
    LocalMux I__3092 (
            .O(N__12753),
            .I(N__12747));
    LocalMux I__3091 (
            .O(N__12750),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    Odrv4 I__3090 (
            .O(N__12747),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    CascadeMux I__3089 (
            .O(N__12742),
            .I(N__12739));
    InMux I__3088 (
            .O(N__12739),
            .I(N__12725));
    InMux I__3087 (
            .O(N__12738),
            .I(N__12725));
    InMux I__3086 (
            .O(N__12737),
            .I(N__12725));
    InMux I__3085 (
            .O(N__12736),
            .I(N__12716));
    InMux I__3084 (
            .O(N__12735),
            .I(N__12716));
    InMux I__3083 (
            .O(N__12734),
            .I(N__12716));
    InMux I__3082 (
            .O(N__12733),
            .I(N__12716));
    InMux I__3081 (
            .O(N__12732),
            .I(N__12713));
    LocalMux I__3080 (
            .O(N__12725),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__3079 (
            .O(N__12716),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__3078 (
            .O(N__12713),
            .I(\U409_TICK.TICK503_14 ));
    CascadeMux I__3077 (
            .O(N__12706),
            .I(N__12698));
    InMux I__3076 (
            .O(N__12705),
            .I(N__12687));
    InMux I__3075 (
            .O(N__12704),
            .I(N__12687));
    InMux I__3074 (
            .O(N__12703),
            .I(N__12687));
    InMux I__3073 (
            .O(N__12702),
            .I(N__12687));
    InMux I__3072 (
            .O(N__12701),
            .I(N__12684));
    InMux I__3071 (
            .O(N__12698),
            .I(N__12677));
    InMux I__3070 (
            .O(N__12697),
            .I(N__12677));
    InMux I__3069 (
            .O(N__12696),
            .I(N__12677));
    LocalMux I__3068 (
            .O(N__12687),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__3067 (
            .O(N__12684),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__3066 (
            .O(N__12677),
            .I(\U409_TICK.TICK503_9 ));
    CascadeMux I__3065 (
            .O(N__12670),
            .I(N__12665));
    CascadeMux I__3064 (
            .O(N__12669),
            .I(N__12657));
    CascadeMux I__3063 (
            .O(N__12668),
            .I(N__12654));
    InMux I__3062 (
            .O(N__12665),
            .I(N__12651));
    InMux I__3061 (
            .O(N__12664),
            .I(N__12642));
    InMux I__3060 (
            .O(N__12663),
            .I(N__12642));
    InMux I__3059 (
            .O(N__12662),
            .I(N__12642));
    InMux I__3058 (
            .O(N__12661),
            .I(N__12642));
    InMux I__3057 (
            .O(N__12660),
            .I(N__12635));
    InMux I__3056 (
            .O(N__12657),
            .I(N__12635));
    InMux I__3055 (
            .O(N__12654),
            .I(N__12635));
    LocalMux I__3054 (
            .O(N__12651),
            .I(N__12632));
    LocalMux I__3053 (
            .O(N__12642),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__3052 (
            .O(N__12635),
            .I(\U409_TICK.TICK503_10 ));
    Odrv12 I__3051 (
            .O(N__12632),
            .I(\U409_TICK.TICK503_10 ));
    InMux I__3050 (
            .O(N__12625),
            .I(N__12622));
    LocalMux I__3049 (
            .O(N__12622),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ));
    InMux I__3048 (
            .O(N__12619),
            .I(N__12615));
    InMux I__3047 (
            .O(N__12618),
            .I(N__12612));
    LocalMux I__3046 (
            .O(N__12615),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    LocalMux I__3045 (
            .O(N__12612),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    ClkMux I__3044 (
            .O(N__12607),
            .I(N__12577));
    ClkMux I__3043 (
            .O(N__12606),
            .I(N__12577));
    ClkMux I__3042 (
            .O(N__12605),
            .I(N__12577));
    ClkMux I__3041 (
            .O(N__12604),
            .I(N__12577));
    ClkMux I__3040 (
            .O(N__12603),
            .I(N__12577));
    ClkMux I__3039 (
            .O(N__12602),
            .I(N__12577));
    ClkMux I__3038 (
            .O(N__12601),
            .I(N__12577));
    ClkMux I__3037 (
            .O(N__12600),
            .I(N__12577));
    ClkMux I__3036 (
            .O(N__12599),
            .I(N__12577));
    ClkMux I__3035 (
            .O(N__12598),
            .I(N__12577));
    GlobalMux I__3034 (
            .O(N__12577),
            .I(N__12574));
    gio2CtrlBuf I__3033 (
            .O(N__12574),
            .I(CLK6_c_g));
    IoInMux I__3032 (
            .O(N__12571),
            .I(N__12568));
    LocalMux I__3031 (
            .O(N__12568),
            .I(N__12565));
    IoSpan4Mux I__3030 (
            .O(N__12565),
            .I(N__12562));
    Sp12to4 I__3029 (
            .O(N__12562),
            .I(N__12559));
    Span12Mux_s9_h I__3028 (
            .O(N__12559),
            .I(N__12556));
    Odrv12 I__3027 (
            .O(N__12556),
            .I(PCS0_c));
    IoInMux I__3026 (
            .O(N__12553),
            .I(N__12550));
    LocalMux I__3025 (
            .O(N__12550),
            .I(N__12547));
    IoSpan4Mux I__3024 (
            .O(N__12547),
            .I(N__12544));
    IoSpan4Mux I__3023 (
            .O(N__12544),
            .I(N__12541));
    Span4Mux_s2_h I__3022 (
            .O(N__12541),
            .I(N__12538));
    Span4Mux_h I__3021 (
            .O(N__12538),
            .I(N__12535));
    Odrv4 I__3020 (
            .O(N__12535),
            .I(SCS1_c));
    InMux I__3019 (
            .O(N__12532),
            .I(N__12529));
    LocalMux I__3018 (
            .O(N__12529),
            .I(N__12525));
    InMux I__3017 (
            .O(N__12528),
            .I(N__12522));
    Span4Mux_v I__3016 (
            .O(N__12525),
            .I(N__12519));
    LocalMux I__3015 (
            .O(N__12522),
            .I(N__12516));
    Span4Mux_h I__3014 (
            .O(N__12519),
            .I(N__12513));
    Span12Mux_s8_v I__3013 (
            .O(N__12516),
            .I(N__12510));
    Odrv4 I__3012 (
            .O(N__12513),
            .I(\U409_ADDRESS_DECODE.CSZ0Z0 ));
    Odrv12 I__3011 (
            .O(N__12510),
            .I(\U409_ADDRESS_DECODE.CSZ0Z0 ));
    IoInMux I__3010 (
            .O(N__12505),
            .I(N__12502));
    LocalMux I__3009 (
            .O(N__12502),
            .I(N__12499));
    Span4Mux_s2_h I__3008 (
            .O(N__12499),
            .I(N__12496));
    Sp12to4 I__3007 (
            .O(N__12496),
            .I(N__12493));
    Span12Mux_s7_v I__3006 (
            .O(N__12493),
            .I(N__12490));
    Odrv12 I__3005 (
            .O(N__12490),
            .I(PCS1_c));
    InMux I__3004 (
            .O(N__12487),
            .I(N__12483));
    InMux I__3003 (
            .O(N__12486),
            .I(N__12480));
    LocalMux I__3002 (
            .O(N__12483),
            .I(N__12475));
    LocalMux I__3001 (
            .O(N__12480),
            .I(N__12475));
    Odrv12 I__3000 (
            .O(N__12475),
            .I(\U409_ADDRESS_DECODE.CSZ0Z1 ));
    InMux I__2999 (
            .O(N__12472),
            .I(N__12466));
    InMux I__2998 (
            .O(N__12471),
            .I(N__12463));
    InMux I__2997 (
            .O(N__12470),
            .I(N__12460));
    InMux I__2996 (
            .O(N__12469),
            .I(N__12457));
    LocalMux I__2995 (
            .O(N__12466),
            .I(N__12452));
    LocalMux I__2994 (
            .O(N__12463),
            .I(N__12452));
    LocalMux I__2993 (
            .O(N__12460),
            .I(N__12447));
    LocalMux I__2992 (
            .O(N__12457),
            .I(N__12447));
    Span4Mux_v I__2991 (
            .O(N__12452),
            .I(N__12444));
    Span12Mux_v I__2990 (
            .O(N__12447),
            .I(N__12439));
    Sp12to4 I__2989 (
            .O(N__12444),
            .I(N__12439));
    Span12Mux_h I__2988 (
            .O(N__12439),
            .I(N__12436));
    Odrv12 I__2987 (
            .O(N__12436),
            .I(A_c_14));
    IoInMux I__2986 (
            .O(N__12433),
            .I(N__12430));
    LocalMux I__2985 (
            .O(N__12430),
            .I(N__12427));
    Span4Mux_s3_h I__2984 (
            .O(N__12427),
            .I(N__12424));
    Span4Mux_v I__2983 (
            .O(N__12424),
            .I(N__12421));
    Span4Mux_h I__2982 (
            .O(N__12421),
            .I(N__12418));
    Odrv4 I__2981 (
            .O(N__12418),
            .I(SCS0_c));
    CascadeMux I__2980 (
            .O(N__12415),
            .I(N__12411));
    CascadeMux I__2979 (
            .O(N__12414),
            .I(N__12408));
    InMux I__2978 (
            .O(N__12411),
            .I(N__12405));
    InMux I__2977 (
            .O(N__12408),
            .I(N__12402));
    LocalMux I__2976 (
            .O(N__12405),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    LocalMux I__2975 (
            .O(N__12402),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    InMux I__2974 (
            .O(N__12397),
            .I(N__12394));
    LocalMux I__2973 (
            .O(N__12394),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ));
    InMux I__2972 (
            .O(N__12391),
            .I(\U409_TICK.un2_COUNTER50_1_cry_5 ));
    InMux I__2971 (
            .O(N__12388),
            .I(N__12384));
    InMux I__2970 (
            .O(N__12387),
            .I(N__12381));
    LocalMux I__2969 (
            .O(N__12384),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    LocalMux I__2968 (
            .O(N__12381),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    InMux I__2967 (
            .O(N__12376),
            .I(\U409_TICK.un2_COUNTER50_1_cry_6 ));
    InMux I__2966 (
            .O(N__12373),
            .I(N__12369));
    InMux I__2965 (
            .O(N__12372),
            .I(N__12366));
    LocalMux I__2964 (
            .O(N__12369),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    LocalMux I__2963 (
            .O(N__12366),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    InMux I__2962 (
            .O(N__12361),
            .I(\U409_TICK.un2_COUNTER50_1_cry_7 ));
    InMux I__2961 (
            .O(N__12358),
            .I(N__12354));
    InMux I__2960 (
            .O(N__12357),
            .I(N__12351));
    LocalMux I__2959 (
            .O(N__12354),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    LocalMux I__2958 (
            .O(N__12351),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    InMux I__2957 (
            .O(N__12346),
            .I(N__12343));
    LocalMux I__2956 (
            .O(N__12343),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ));
    InMux I__2955 (
            .O(N__12340),
            .I(bfn_17_6_0_));
    InMux I__2954 (
            .O(N__12337),
            .I(N__12334));
    LocalMux I__2953 (
            .O(N__12334),
            .I(N__12330));
    InMux I__2952 (
            .O(N__12333),
            .I(N__12327));
    Odrv4 I__2951 (
            .O(N__12330),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    LocalMux I__2950 (
            .O(N__12327),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    InMux I__2949 (
            .O(N__12322),
            .I(\U409_TICK.un2_COUNTER50_1_cry_9 ));
    InMux I__2948 (
            .O(N__12319),
            .I(\U409_TICK.un2_COUNTER50_1_cry_10 ));
    InMux I__2947 (
            .O(N__12316),
            .I(N__12313));
    LocalMux I__2946 (
            .O(N__12313),
            .I(N__12309));
    InMux I__2945 (
            .O(N__12312),
            .I(N__12306));
    Odrv4 I__2944 (
            .O(N__12309),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    LocalMux I__2943 (
            .O(N__12306),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    InMux I__2942 (
            .O(N__12301),
            .I(\U409_TICK.un2_COUNTER50_1_cry_11 ));
    InMux I__2941 (
            .O(N__12298),
            .I(N__12294));
    InMux I__2940 (
            .O(N__12297),
            .I(N__12291));
    LocalMux I__2939 (
            .O(N__12294),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    LocalMux I__2938 (
            .O(N__12291),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    InMux I__2937 (
            .O(N__12286),
            .I(N__12283));
    LocalMux I__2936 (
            .O(N__12283),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ));
    InMux I__2935 (
            .O(N__12280),
            .I(\U409_TICK.un2_COUNTER50_1_cry_12 ));
    IoInMux I__2934 (
            .O(N__12277),
            .I(N__12274));
    LocalMux I__2933 (
            .O(N__12274),
            .I(N__12271));
    Span4Mux_s1_v I__2932 (
            .O(N__12271),
            .I(N__12268));
    Span4Mux_v I__2931 (
            .O(N__12268),
            .I(N__12265));
    Span4Mux_v I__2930 (
            .O(N__12265),
            .I(N__12262));
    Span4Mux_h I__2929 (
            .O(N__12262),
            .I(N__12258));
    InMux I__2928 (
            .O(N__12261),
            .I(N__12255));
    Odrv4 I__2927 (
            .O(N__12258),
            .I(TICK50_c));
    LocalMux I__2926 (
            .O(N__12255),
            .I(TICK50_c));
    CascadeMux I__2925 (
            .O(N__12250),
            .I(\U409_TICK.TICK503_9_cascade_ ));
    InMux I__2924 (
            .O(N__12247),
            .I(N__12243));
    InMux I__2923 (
            .O(N__12246),
            .I(N__12239));
    LocalMux I__2922 (
            .O(N__12243),
            .I(N__12236));
    InMux I__2921 (
            .O(N__12242),
            .I(N__12233));
    LocalMux I__2920 (
            .O(N__12239),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    Odrv4 I__2919 (
            .O(N__12236),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__2918 (
            .O(N__12233),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    InMux I__2917 (
            .O(N__12226),
            .I(N__12222));
    CascadeMux I__2916 (
            .O(N__12225),
            .I(N__12217));
    LocalMux I__2915 (
            .O(N__12222),
            .I(N__12214));
    InMux I__2914 (
            .O(N__12221),
            .I(N__12209));
    InMux I__2913 (
            .O(N__12220),
            .I(N__12209));
    InMux I__2912 (
            .O(N__12217),
            .I(N__12206));
    Odrv4 I__2911 (
            .O(N__12214),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__2910 (
            .O(N__12209),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__2909 (
            .O(N__12206),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    CascadeMux I__2908 (
            .O(N__12199),
            .I(N__12196));
    InMux I__2907 (
            .O(N__12196),
            .I(N__12192));
    InMux I__2906 (
            .O(N__12195),
            .I(N__12189));
    LocalMux I__2905 (
            .O(N__12192),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    LocalMux I__2904 (
            .O(N__12189),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    InMux I__2903 (
            .O(N__12184),
            .I(\U409_TICK.un2_COUNTER50_1_cry_1 ));
    InMux I__2902 (
            .O(N__12181),
            .I(N__12177));
    InMux I__2901 (
            .O(N__12180),
            .I(N__12174));
    LocalMux I__2900 (
            .O(N__12177),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    LocalMux I__2899 (
            .O(N__12174),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    InMux I__2898 (
            .O(N__12169),
            .I(\U409_TICK.un2_COUNTER50_1_cry_2 ));
    CascadeMux I__2897 (
            .O(N__12166),
            .I(N__12163));
    InMux I__2896 (
            .O(N__12163),
            .I(N__12159));
    InMux I__2895 (
            .O(N__12162),
            .I(N__12156));
    LocalMux I__2894 (
            .O(N__12159),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    LocalMux I__2893 (
            .O(N__12156),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    InMux I__2892 (
            .O(N__12151),
            .I(\U409_TICK.un2_COUNTER50_1_cry_3 ));
    InMux I__2891 (
            .O(N__12148),
            .I(N__12144));
    InMux I__2890 (
            .O(N__12147),
            .I(N__12141));
    LocalMux I__2889 (
            .O(N__12144),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    LocalMux I__2888 (
            .O(N__12141),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    InMux I__2887 (
            .O(N__12136),
            .I(N__12133));
    LocalMux I__2886 (
            .O(N__12133),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ));
    InMux I__2885 (
            .O(N__12130),
            .I(\U409_TICK.un2_COUNTER50_1_cry_4 ));
    CascadeMux I__2884 (
            .O(N__12127),
            .I(\U409_TICK.TICK503_10_cascade_ ));
    CascadeMux I__2883 (
            .O(N__12124),
            .I(N__12117));
    InMux I__2882 (
            .O(N__12123),
            .I(N__12112));
    InMux I__2881 (
            .O(N__12122),
            .I(N__12103));
    InMux I__2880 (
            .O(N__12121),
            .I(N__12103));
    InMux I__2879 (
            .O(N__12120),
            .I(N__12103));
    InMux I__2878 (
            .O(N__12117),
            .I(N__12103));
    InMux I__2877 (
            .O(N__12116),
            .I(N__12098));
    InMux I__2876 (
            .O(N__12115),
            .I(N__12098));
    LocalMux I__2875 (
            .O(N__12112),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__2874 (
            .O(N__12103),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__2873 (
            .O(N__12098),
            .I(\U409_TICK.TICK603_10 ));
    CascadeMux I__2872 (
            .O(N__12091),
            .I(N__12087));
    CascadeMux I__2871 (
            .O(N__12090),
            .I(N__12083));
    InMux I__2870 (
            .O(N__12087),
            .I(N__12076));
    InMux I__2869 (
            .O(N__12086),
            .I(N__12069));
    InMux I__2868 (
            .O(N__12083),
            .I(N__12069));
    InMux I__2867 (
            .O(N__12082),
            .I(N__12069));
    InMux I__2866 (
            .O(N__12081),
            .I(N__12062));
    InMux I__2865 (
            .O(N__12080),
            .I(N__12062));
    InMux I__2864 (
            .O(N__12079),
            .I(N__12062));
    LocalMux I__2863 (
            .O(N__12076),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__2862 (
            .O(N__12069),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__2861 (
            .O(N__12062),
            .I(\U409_TICK.TICK603_9 ));
    InMux I__2860 (
            .O(N__12055),
            .I(N__12046));
    InMux I__2859 (
            .O(N__12054),
            .I(N__12041));
    InMux I__2858 (
            .O(N__12053),
            .I(N__12041));
    InMux I__2857 (
            .O(N__12052),
            .I(N__12032));
    InMux I__2856 (
            .O(N__12051),
            .I(N__12032));
    InMux I__2855 (
            .O(N__12050),
            .I(N__12032));
    InMux I__2854 (
            .O(N__12049),
            .I(N__12032));
    LocalMux I__2853 (
            .O(N__12046),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__2852 (
            .O(N__12041),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__2851 (
            .O(N__12032),
            .I(\U409_TICK.TICK603_14 ));
    IoInMux I__2850 (
            .O(N__12025),
            .I(N__12022));
    LocalMux I__2849 (
            .O(N__12022),
            .I(N__12019));
    Span4Mux_s3_v I__2848 (
            .O(N__12019),
            .I(N__12016));
    Sp12to4 I__2847 (
            .O(N__12016),
            .I(N__12013));
    Span12Mux_h I__2846 (
            .O(N__12013),
            .I(N__12009));
    InMux I__2845 (
            .O(N__12012),
            .I(N__12006));
    Odrv12 I__2844 (
            .O(N__12009),
            .I(TICK60_c));
    LocalMux I__2843 (
            .O(N__12006),
            .I(TICK60_c));
    IoInMux I__2842 (
            .O(N__12001),
            .I(N__11997));
    IoInMux I__2841 (
            .O(N__12000),
            .I(N__11994));
    LocalMux I__2840 (
            .O(N__11997),
            .I(N__11988));
    LocalMux I__2839 (
            .O(N__11994),
            .I(N__11988));
    IoInMux I__2838 (
            .O(N__11993),
            .I(N__11985));
    IoSpan4Mux I__2837 (
            .O(N__11988),
            .I(N__11982));
    LocalMux I__2836 (
            .O(N__11985),
            .I(N__11978));
    Span4Mux_s0_h I__2835 (
            .O(N__11982),
            .I(N__11974));
    IoInMux I__2834 (
            .O(N__11981),
            .I(N__11971));
    Span4Mux_s0_v I__2833 (
            .O(N__11978),
            .I(N__11968));
    IoInMux I__2832 (
            .O(N__11977),
            .I(N__11965));
    Sp12to4 I__2831 (
            .O(N__11974),
            .I(N__11962));
    LocalMux I__2830 (
            .O(N__11971),
            .I(N__11959));
    Span4Mux_v I__2829 (
            .O(N__11968),
            .I(N__11956));
    LocalMux I__2828 (
            .O(N__11965),
            .I(N__11953));
    Span12Mux_v I__2827 (
            .O(N__11962),
            .I(N__11948));
    Span12Mux_s8_v I__2826 (
            .O(N__11959),
            .I(N__11948));
    Span4Mux_v I__2825 (
            .O(N__11956),
            .I(N__11945));
    Span12Mux_s8_v I__2824 (
            .O(N__11953),
            .I(N__11942));
    Odrv12 I__2823 (
            .O(N__11948),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2822 (
            .O(N__11945),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__2821 (
            .O(N__11942),
            .I(CONSTANT_ONE_NET));
    InMux I__2820 (
            .O(N__11935),
            .I(N__11932));
    LocalMux I__2819 (
            .O(N__11932),
            .I(\U409_TICK.TICK503_8 ));
    CascadeMux I__2818 (
            .O(N__11929),
            .I(\U409_TICK.TICK503_11_cascade_ ));
    CascadeMux I__2817 (
            .O(N__11926),
            .I(\U409_TICK.TICK503_14_cascade_ ));
    InMux I__2816 (
            .O(N__11923),
            .I(N__11914));
    InMux I__2815 (
            .O(N__11922),
            .I(N__11914));
    InMux I__2814 (
            .O(N__11921),
            .I(N__11914));
    LocalMux I__2813 (
            .O(N__11914),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    InMux I__2812 (
            .O(N__11911),
            .I(N__11905));
    InMux I__2811 (
            .O(N__11910),
            .I(N__11898));
    InMux I__2810 (
            .O(N__11909),
            .I(N__11898));
    InMux I__2809 (
            .O(N__11908),
            .I(N__11898));
    LocalMux I__2808 (
            .O(N__11905),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__2807 (
            .O(N__11898),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    InMux I__2806 (
            .O(N__11893),
            .I(N__11890));
    LocalMux I__2805 (
            .O(N__11890),
            .I(\U409_TRANSFER_ACK.N_3_0 ));
    InMux I__2804 (
            .O(N__11887),
            .I(N__11884));
    LocalMux I__2803 (
            .O(N__11884),
            .I(N__11880));
    InMux I__2802 (
            .O(N__11883),
            .I(N__11877));
    Span4Mux_v I__2801 (
            .O(N__11880),
            .I(N__11870));
    LocalMux I__2800 (
            .O(N__11877),
            .I(N__11870));
    InMux I__2799 (
            .O(N__11876),
            .I(N__11867));
    InMux I__2798 (
            .O(N__11875),
            .I(N__11864));
    Span4Mux_v I__2797 (
            .O(N__11870),
            .I(N__11859));
    LocalMux I__2796 (
            .O(N__11867),
            .I(N__11859));
    LocalMux I__2795 (
            .O(N__11864),
            .I(N__11856));
    Span4Mux_v I__2794 (
            .O(N__11859),
            .I(N__11843));
    Span4Mux_v I__2793 (
            .O(N__11856),
            .I(N__11839));
    InMux I__2792 (
            .O(N__11855),
            .I(N__11829));
    InMux I__2791 (
            .O(N__11854),
            .I(N__11829));
    InMux I__2790 (
            .O(N__11853),
            .I(N__11829));
    InMux I__2789 (
            .O(N__11852),
            .I(N__11826));
    InMux I__2788 (
            .O(N__11851),
            .I(N__11821));
    InMux I__2787 (
            .O(N__11850),
            .I(N__11821));
    InMux I__2786 (
            .O(N__11849),
            .I(N__11816));
    InMux I__2785 (
            .O(N__11848),
            .I(N__11816));
    InMux I__2784 (
            .O(N__11847),
            .I(N__11810));
    InMux I__2783 (
            .O(N__11846),
            .I(N__11810));
    Span4Mux_h I__2782 (
            .O(N__11843),
            .I(N__11806));
    InMux I__2781 (
            .O(N__11842),
            .I(N__11803));
    Span4Mux_h I__2780 (
            .O(N__11839),
            .I(N__11800));
    InMux I__2779 (
            .O(N__11838),
            .I(N__11797));
    InMux I__2778 (
            .O(N__11837),
            .I(N__11792));
    CascadeMux I__2777 (
            .O(N__11836),
            .I(N__11789));
    LocalMux I__2776 (
            .O(N__11829),
            .I(N__11779));
    LocalMux I__2775 (
            .O(N__11826),
            .I(N__11779));
    LocalMux I__2774 (
            .O(N__11821),
            .I(N__11779));
    LocalMux I__2773 (
            .O(N__11816),
            .I(N__11779));
    InMux I__2772 (
            .O(N__11815),
            .I(N__11776));
    LocalMux I__2771 (
            .O(N__11810),
            .I(N__11772));
    InMux I__2770 (
            .O(N__11809),
            .I(N__11769));
    Span4Mux_h I__2769 (
            .O(N__11806),
            .I(N__11764));
    LocalMux I__2768 (
            .O(N__11803),
            .I(N__11764));
    Span4Mux_h I__2767 (
            .O(N__11800),
            .I(N__11759));
    LocalMux I__2766 (
            .O(N__11797),
            .I(N__11759));
    InMux I__2765 (
            .O(N__11796),
            .I(N__11756));
    InMux I__2764 (
            .O(N__11795),
            .I(N__11753));
    LocalMux I__2763 (
            .O(N__11792),
            .I(N__11750));
    InMux I__2762 (
            .O(N__11789),
            .I(N__11745));
    InMux I__2761 (
            .O(N__11788),
            .I(N__11745));
    Span4Mux_v I__2760 (
            .O(N__11779),
            .I(N__11740));
    LocalMux I__2759 (
            .O(N__11776),
            .I(N__11740));
    CascadeMux I__2758 (
            .O(N__11775),
            .I(N__11735));
    Span4Mux_v I__2757 (
            .O(N__11772),
            .I(N__11732));
    LocalMux I__2756 (
            .O(N__11769),
            .I(N__11728));
    Span4Mux_v I__2755 (
            .O(N__11764),
            .I(N__11725));
    Span4Mux_v I__2754 (
            .O(N__11759),
            .I(N__11722));
    LocalMux I__2753 (
            .O(N__11756),
            .I(N__11719));
    LocalMux I__2752 (
            .O(N__11753),
            .I(N__11716));
    Span4Mux_h I__2751 (
            .O(N__11750),
            .I(N__11711));
    LocalMux I__2750 (
            .O(N__11745),
            .I(N__11711));
    Span4Mux_h I__2749 (
            .O(N__11740),
            .I(N__11708));
    InMux I__2748 (
            .O(N__11739),
            .I(N__11701));
    InMux I__2747 (
            .O(N__11738),
            .I(N__11701));
    InMux I__2746 (
            .O(N__11735),
            .I(N__11701));
    Span4Mux_h I__2745 (
            .O(N__11732),
            .I(N__11698));
    InMux I__2744 (
            .O(N__11731),
            .I(N__11695));
    Span12Mux_h I__2743 (
            .O(N__11728),
            .I(N__11692));
    Sp12to4 I__2742 (
            .O(N__11725),
            .I(N__11687));
    Sp12to4 I__2741 (
            .O(N__11722),
            .I(N__11687));
    Span12Mux_v I__2740 (
            .O(N__11719),
            .I(N__11672));
    Sp12to4 I__2739 (
            .O(N__11716),
            .I(N__11672));
    Sp12to4 I__2738 (
            .O(N__11711),
            .I(N__11672));
    Sp12to4 I__2737 (
            .O(N__11708),
            .I(N__11672));
    LocalMux I__2736 (
            .O(N__11701),
            .I(N__11672));
    Sp12to4 I__2735 (
            .O(N__11698),
            .I(N__11672));
    LocalMux I__2734 (
            .O(N__11695),
            .I(N__11672));
    Span12Mux_v I__2733 (
            .O(N__11692),
            .I(N__11669));
    Span12Mux_h I__2732 (
            .O(N__11687),
            .I(N__11666));
    Span12Mux_v I__2731 (
            .O(N__11672),
            .I(N__11663));
    Span12Mux_h I__2730 (
            .O(N__11669),
            .I(N__11660));
    Span12Mux_v I__2729 (
            .O(N__11666),
            .I(N__11655));
    Span12Mux_h I__2728 (
            .O(N__11663),
            .I(N__11655));
    Odrv12 I__2727 (
            .O(N__11660),
            .I(RESETn_c));
    Odrv12 I__2726 (
            .O(N__11655),
            .I(RESETn_c));
    CascadeMux I__2725 (
            .O(N__11650),
            .I(N__11645));
    InMux I__2724 (
            .O(N__11649),
            .I(N__11640));
    InMux I__2723 (
            .O(N__11648),
            .I(N__11640));
    InMux I__2722 (
            .O(N__11645),
            .I(N__11637));
    LocalMux I__2721 (
            .O(N__11640),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__2720 (
            .O(N__11637),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    CascadeMux I__2719 (
            .O(N__11632),
            .I(\U409_TRANSFER_ACK.N_55_cascade_ ));
    CascadeMux I__2718 (
            .O(N__11629),
            .I(N__11622));
    CascadeMux I__2717 (
            .O(N__11628),
            .I(N__11619));
    InMux I__2716 (
            .O(N__11627),
            .I(N__11616));
    InMux I__2715 (
            .O(N__11626),
            .I(N__11607));
    InMux I__2714 (
            .O(N__11625),
            .I(N__11607));
    InMux I__2713 (
            .O(N__11622),
            .I(N__11607));
    InMux I__2712 (
            .O(N__11619),
            .I(N__11607));
    LocalMux I__2711 (
            .O(N__11616),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__2710 (
            .O(N__11607),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    InMux I__2709 (
            .O(N__11602),
            .I(N__11596));
    InMux I__2708 (
            .O(N__11601),
            .I(N__11596));
    LocalMux I__2707 (
            .O(N__11596),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    IoInMux I__2706 (
            .O(N__11593),
            .I(N__11590));
    LocalMux I__2705 (
            .O(N__11590),
            .I(N__11587));
    Span4Mux_s3_v I__2704 (
            .O(N__11587),
            .I(N__11583));
    InMux I__2703 (
            .O(N__11586),
            .I(N__11580));
    Span4Mux_h I__2702 (
            .O(N__11583),
            .I(N__11577));
    LocalMux I__2701 (
            .O(N__11580),
            .I(N__11574));
    Span4Mux_h I__2700 (
            .O(N__11577),
            .I(N__11570));
    Span4Mux_v I__2699 (
            .O(N__11574),
            .I(N__11567));
    CascadeMux I__2698 (
            .O(N__11573),
            .I(N__11563));
    Sp12to4 I__2697 (
            .O(N__11570),
            .I(N__11560));
    Span4Mux_h I__2696 (
            .O(N__11567),
            .I(N__11557));
    InMux I__2695 (
            .O(N__11566),
            .I(N__11554));
    InMux I__2694 (
            .O(N__11563),
            .I(N__11551));
    Odrv12 I__2693 (
            .O(N__11560),
            .I(CLK_CIA_c));
    Odrv4 I__2692 (
            .O(N__11557),
            .I(CLK_CIA_c));
    LocalMux I__2691 (
            .O(N__11554),
            .I(CLK_CIA_c));
    LocalMux I__2690 (
            .O(N__11551),
            .I(CLK_CIA_c));
    InMux I__2689 (
            .O(N__11542),
            .I(N__11537));
    InMux I__2688 (
            .O(N__11541),
            .I(N__11532));
    InMux I__2687 (
            .O(N__11540),
            .I(N__11532));
    LocalMux I__2686 (
            .O(N__11537),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__2685 (
            .O(N__11532),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    InMux I__2684 (
            .O(N__11527),
            .I(N__11524));
    LocalMux I__2683 (
            .O(N__11524),
            .I(N__11521));
    Odrv4 I__2682 (
            .O(N__11521),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0 ));
    InMux I__2681 (
            .O(N__11518),
            .I(N__11515));
    LocalMux I__2680 (
            .O(N__11515),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0 ));
    CascadeMux I__2679 (
            .O(N__11512),
            .I(N__11509));
    InMux I__2678 (
            .O(N__11509),
            .I(N__11506));
    LocalMux I__2677 (
            .O(N__11506),
            .I(N__11502));
    InMux I__2676 (
            .O(N__11505),
            .I(N__11499));
    Span4Mux_v I__2675 (
            .O(N__11502),
            .I(N__11494));
    LocalMux I__2674 (
            .O(N__11499),
            .I(N__11491));
    InMux I__2673 (
            .O(N__11498),
            .I(N__11488));
    CascadeMux I__2672 (
            .O(N__11497),
            .I(N__11485));
    Span4Mux_h I__2671 (
            .O(N__11494),
            .I(N__11482));
    Span4Mux_v I__2670 (
            .O(N__11491),
            .I(N__11479));
    LocalMux I__2669 (
            .O(N__11488),
            .I(N__11476));
    InMux I__2668 (
            .O(N__11485),
            .I(N__11473));
    Odrv4 I__2667 (
            .O(N__11482),
            .I(N_52_1));
    Odrv4 I__2666 (
            .O(N__11479),
            .I(N_52_1));
    Odrv4 I__2665 (
            .O(N__11476),
            .I(N_52_1));
    LocalMux I__2664 (
            .O(N__11473),
            .I(N_52_1));
    InMux I__2663 (
            .O(N__11464),
            .I(N__11460));
    InMux I__2662 (
            .O(N__11463),
            .I(N__11455));
    LocalMux I__2661 (
            .O(N__11460),
            .I(N__11452));
    InMux I__2660 (
            .O(N__11459),
            .I(N__11447));
    InMux I__2659 (
            .O(N__11458),
            .I(N__11447));
    LocalMux I__2658 (
            .O(N__11455),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ));
    Odrv4 I__2657 (
            .O(N__11452),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ));
    LocalMux I__2656 (
            .O(N__11447),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ));
    InMux I__2655 (
            .O(N__11440),
            .I(N__11437));
    LocalMux I__2654 (
            .O(N__11437),
            .I(N__11431));
    InMux I__2653 (
            .O(N__11436),
            .I(N__11426));
    InMux I__2652 (
            .O(N__11435),
            .I(N__11421));
    InMux I__2651 (
            .O(N__11434),
            .I(N__11421));
    Span4Mux_h I__2650 (
            .O(N__11431),
            .I(N__11417));
    InMux I__2649 (
            .O(N__11430),
            .I(N__11412));
    InMux I__2648 (
            .O(N__11429),
            .I(N__11412));
    LocalMux I__2647 (
            .O(N__11426),
            .I(N__11407));
    LocalMux I__2646 (
            .O(N__11421),
            .I(N__11407));
    InMux I__2645 (
            .O(N__11420),
            .I(N__11404));
    Odrv4 I__2644 (
            .O(N__11417),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__2643 (
            .O(N__11412),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    Odrv4 I__2642 (
            .O(N__11407),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__2641 (
            .O(N__11404),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    SRMux I__2640 (
            .O(N__11395),
            .I(N__11353));
    SRMux I__2639 (
            .O(N__11394),
            .I(N__11353));
    SRMux I__2638 (
            .O(N__11393),
            .I(N__11353));
    SRMux I__2637 (
            .O(N__11392),
            .I(N__11353));
    SRMux I__2636 (
            .O(N__11391),
            .I(N__11353));
    SRMux I__2635 (
            .O(N__11390),
            .I(N__11353));
    SRMux I__2634 (
            .O(N__11389),
            .I(N__11353));
    SRMux I__2633 (
            .O(N__11388),
            .I(N__11353));
    SRMux I__2632 (
            .O(N__11387),
            .I(N__11353));
    SRMux I__2631 (
            .O(N__11386),
            .I(N__11353));
    SRMux I__2630 (
            .O(N__11385),
            .I(N__11353));
    SRMux I__2629 (
            .O(N__11384),
            .I(N__11353));
    SRMux I__2628 (
            .O(N__11383),
            .I(N__11353));
    SRMux I__2627 (
            .O(N__11382),
            .I(N__11353));
    GlobalMux I__2626 (
            .O(N__11353),
            .I(N__11350));
    gio2CtrlBuf I__2625 (
            .O(N__11350),
            .I(RESETn_c_i_g));
    InMux I__2624 (
            .O(N__11347),
            .I(N__11343));
    InMux I__2623 (
            .O(N__11346),
            .I(N__11340));
    LocalMux I__2622 (
            .O(N__11343),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    LocalMux I__2621 (
            .O(N__11340),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    InMux I__2620 (
            .O(N__11335),
            .I(N__11331));
    InMux I__2619 (
            .O(N__11334),
            .I(N__11328));
    LocalMux I__2618 (
            .O(N__11331),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    LocalMux I__2617 (
            .O(N__11328),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    CascadeMux I__2616 (
            .O(N__11323),
            .I(N__11320));
    InMux I__2615 (
            .O(N__11320),
            .I(N__11316));
    InMux I__2614 (
            .O(N__11319),
            .I(N__11312));
    LocalMux I__2613 (
            .O(N__11316),
            .I(N__11309));
    InMux I__2612 (
            .O(N__11315),
            .I(N__11306));
    LocalMux I__2611 (
            .O(N__11312),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    Odrv12 I__2610 (
            .O(N__11309),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__2609 (
            .O(N__11306),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    InMux I__2608 (
            .O(N__11299),
            .I(N__11295));
    InMux I__2607 (
            .O(N__11298),
            .I(N__11292));
    LocalMux I__2606 (
            .O(N__11295),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    LocalMux I__2605 (
            .O(N__11292),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    InMux I__2604 (
            .O(N__11287),
            .I(N__11284));
    LocalMux I__2603 (
            .O(N__11284),
            .I(\U409_TICK.TICK603_8 ));
    InMux I__2602 (
            .O(N__11281),
            .I(N__11277));
    InMux I__2601 (
            .O(N__11280),
            .I(N__11274));
    LocalMux I__2600 (
            .O(N__11277),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    LocalMux I__2599 (
            .O(N__11274),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    CascadeMux I__2598 (
            .O(N__11269),
            .I(\U409_TICK.TICK603_11_cascade_ ));
    InMux I__2597 (
            .O(N__11266),
            .I(N__11262));
    InMux I__2596 (
            .O(N__11265),
            .I(N__11259));
    LocalMux I__2595 (
            .O(N__11262),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    LocalMux I__2594 (
            .O(N__11259),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    CascadeMux I__2593 (
            .O(N__11254),
            .I(\U409_TICK.TICK603_14_cascade_ ));
    InMux I__2592 (
            .O(N__11251),
            .I(N__11248));
    LocalMux I__2591 (
            .O(N__11248),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ));
    InMux I__2590 (
            .O(N__11245),
            .I(N__11241));
    InMux I__2589 (
            .O(N__11244),
            .I(N__11238));
    LocalMux I__2588 (
            .O(N__11241),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    LocalMux I__2587 (
            .O(N__11238),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    CascadeMux I__2586 (
            .O(N__11233),
            .I(N__11230));
    InMux I__2585 (
            .O(N__11230),
            .I(N__11227));
    LocalMux I__2584 (
            .O(N__11227),
            .I(N__11224));
    Odrv4 I__2583 (
            .O(N__11224),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ));
    InMux I__2582 (
            .O(N__11221),
            .I(N__11217));
    InMux I__2581 (
            .O(N__11220),
            .I(N__11214));
    LocalMux I__2580 (
            .O(N__11217),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    LocalMux I__2579 (
            .O(N__11214),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    CascadeMux I__2578 (
            .O(N__11209),
            .I(\U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_ ));
    InMux I__2577 (
            .O(N__11206),
            .I(N__11199));
    InMux I__2576 (
            .O(N__11205),
            .I(N__11196));
    InMux I__2575 (
            .O(N__11204),
            .I(N__11191));
    InMux I__2574 (
            .O(N__11203),
            .I(N__11191));
    InMux I__2573 (
            .O(N__11202),
            .I(N__11188));
    LocalMux I__2572 (
            .O(N__11199),
            .I(N__11184));
    LocalMux I__2571 (
            .O(N__11196),
            .I(N__11176));
    LocalMux I__2570 (
            .O(N__11191),
            .I(N__11166));
    LocalMux I__2569 (
            .O(N__11188),
            .I(N__11162));
    ClkMux I__2568 (
            .O(N__11187),
            .I(N__11122));
    Glb2LocalMux I__2567 (
            .O(N__11184),
            .I(N__11122));
    ClkMux I__2566 (
            .O(N__11183),
            .I(N__11122));
    ClkMux I__2565 (
            .O(N__11182),
            .I(N__11122));
    ClkMux I__2564 (
            .O(N__11181),
            .I(N__11122));
    ClkMux I__2563 (
            .O(N__11180),
            .I(N__11122));
    ClkMux I__2562 (
            .O(N__11179),
            .I(N__11122));
    Glb2LocalMux I__2561 (
            .O(N__11176),
            .I(N__11122));
    ClkMux I__2560 (
            .O(N__11175),
            .I(N__11122));
    ClkMux I__2559 (
            .O(N__11174),
            .I(N__11122));
    ClkMux I__2558 (
            .O(N__11173),
            .I(N__11122));
    ClkMux I__2557 (
            .O(N__11172),
            .I(N__11122));
    ClkMux I__2556 (
            .O(N__11171),
            .I(N__11122));
    ClkMux I__2555 (
            .O(N__11170),
            .I(N__11122));
    ClkMux I__2554 (
            .O(N__11169),
            .I(N__11122));
    Glb2LocalMux I__2553 (
            .O(N__11166),
            .I(N__11122));
    ClkMux I__2552 (
            .O(N__11165),
            .I(N__11122));
    Glb2LocalMux I__2551 (
            .O(N__11162),
            .I(N__11122));
    ClkMux I__2550 (
            .O(N__11161),
            .I(N__11122));
    GlobalMux I__2549 (
            .O(N__11122),
            .I(N__11119));
    gio2CtrlBuf I__2548 (
            .O(N__11119),
            .I(CLK40_IN_c_g));
    InMux I__2547 (
            .O(N__11116),
            .I(N__11112));
    InMux I__2546 (
            .O(N__11115),
            .I(N__11109));
    LocalMux I__2545 (
            .O(N__11112),
            .I(\U409_TRANSFER_ACK.N_17_mux ));
    LocalMux I__2544 (
            .O(N__11109),
            .I(\U409_TRANSFER_ACK.N_17_mux ));
    CascadeMux I__2543 (
            .O(N__11104),
            .I(\U409_TRANSFER_ACK.N_3_0_cascade_ ));
    InMux I__2542 (
            .O(N__11101),
            .I(N__11098));
    LocalMux I__2541 (
            .O(N__11098),
            .I(\U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0 ));
    CascadeMux I__2540 (
            .O(N__11095),
            .I(N__11092));
    InMux I__2539 (
            .O(N__11092),
            .I(N__11089));
    LocalMux I__2538 (
            .O(N__11089),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ));
    InMux I__2537 (
            .O(N__11086),
            .I(N__11082));
    InMux I__2536 (
            .O(N__11085),
            .I(N__11079));
    LocalMux I__2535 (
            .O(N__11082),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    LocalMux I__2534 (
            .O(N__11079),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    InMux I__2533 (
            .O(N__11074),
            .I(N__11071));
    LocalMux I__2532 (
            .O(N__11071),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ));
    InMux I__2531 (
            .O(N__11068),
            .I(N__11064));
    InMux I__2530 (
            .O(N__11067),
            .I(N__11061));
    LocalMux I__2529 (
            .O(N__11064),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    LocalMux I__2528 (
            .O(N__11061),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    InMux I__2527 (
            .O(N__11056),
            .I(N__11052));
    InMux I__2526 (
            .O(N__11055),
            .I(N__11049));
    LocalMux I__2525 (
            .O(N__11052),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    LocalMux I__2524 (
            .O(N__11049),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    CascadeMux I__2523 (
            .O(N__11044),
            .I(N__11040));
    InMux I__2522 (
            .O(N__11043),
            .I(N__11037));
    InMux I__2521 (
            .O(N__11040),
            .I(N__11034));
    LocalMux I__2520 (
            .O(N__11037),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    LocalMux I__2519 (
            .O(N__11034),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    CascadeMux I__2518 (
            .O(N__11029),
            .I(\U409_TICK.TICK603_9_cascade_ ));
    InMux I__2517 (
            .O(N__11026),
            .I(N__11023));
    LocalMux I__2516 (
            .O(N__11023),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ));
    CascadeMux I__2515 (
            .O(N__11020),
            .I(N__11017));
    InMux I__2514 (
            .O(N__11017),
            .I(N__11013));
    InMux I__2513 (
            .O(N__11016),
            .I(N__11010));
    LocalMux I__2512 (
            .O(N__11013),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    LocalMux I__2511 (
            .O(N__11010),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    InMux I__2510 (
            .O(N__11005),
            .I(N__11001));
    InMux I__2509 (
            .O(N__11004),
            .I(N__10998));
    LocalMux I__2508 (
            .O(N__11001),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    LocalMux I__2507 (
            .O(N__10998),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    InMux I__2506 (
            .O(N__10993),
            .I(N__10989));
    InMux I__2505 (
            .O(N__10992),
            .I(N__10986));
    LocalMux I__2504 (
            .O(N__10989),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    LocalMux I__2503 (
            .O(N__10986),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    CascadeMux I__2502 (
            .O(N__10981),
            .I(N__10978));
    InMux I__2501 (
            .O(N__10978),
            .I(N__10974));
    InMux I__2500 (
            .O(N__10977),
            .I(N__10971));
    LocalMux I__2499 (
            .O(N__10974),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    LocalMux I__2498 (
            .O(N__10971),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    CascadeMux I__2497 (
            .O(N__10966),
            .I(\U409_TICK.TICK603_10_cascade_ ));
    CascadeMux I__2496 (
            .O(N__10963),
            .I(N__10957));
    InMux I__2495 (
            .O(N__10962),
            .I(N__10954));
    InMux I__2494 (
            .O(N__10961),
            .I(N__10949));
    InMux I__2493 (
            .O(N__10960),
            .I(N__10949));
    InMux I__2492 (
            .O(N__10957),
            .I(N__10946));
    LocalMux I__2491 (
            .O(N__10954),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__2490 (
            .O(N__10949),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__2489 (
            .O(N__10946),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    InMux I__2488 (
            .O(N__10939),
            .I(N__10935));
    InMux I__2487 (
            .O(N__10938),
            .I(N__10932));
    LocalMux I__2486 (
            .O(N__10935),
            .I(N__10929));
    LocalMux I__2485 (
            .O(N__10932),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    Odrv4 I__2484 (
            .O(N__10929),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    InMux I__2483 (
            .O(N__10924),
            .I(N__10920));
    InMux I__2482 (
            .O(N__10923),
            .I(N__10917));
    LocalMux I__2481 (
            .O(N__10920),
            .I(N__10914));
    LocalMux I__2480 (
            .O(N__10917),
            .I(N__10911));
    Span4Mux_v I__2479 (
            .O(N__10914),
            .I(N__10908));
    Span4Mux_v I__2478 (
            .O(N__10911),
            .I(N__10905));
    Span4Mux_v I__2477 (
            .O(N__10908),
            .I(N__10901));
    Sp12to4 I__2476 (
            .O(N__10905),
            .I(N__10898));
    InMux I__2475 (
            .O(N__10904),
            .I(N__10895));
    Odrv4 I__2474 (
            .O(N__10901),
            .I(\U409_CIA.VMAZ0 ));
    Odrv12 I__2473 (
            .O(N__10898),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__2472 (
            .O(N__10895),
            .I(\U409_CIA.VMAZ0 ));
    InMux I__2471 (
            .O(N__10888),
            .I(N__10884));
    CascadeMux I__2470 (
            .O(N__10887),
            .I(N__10881));
    LocalMux I__2469 (
            .O(N__10884),
            .I(N__10878));
    InMux I__2468 (
            .O(N__10881),
            .I(N__10875));
    Span4Mux_h I__2467 (
            .O(N__10878),
            .I(N__10870));
    LocalMux I__2466 (
            .O(N__10875),
            .I(N__10870));
    Odrv4 I__2465 (
            .O(N__10870),
            .I(\U409_TRANSFER_ACK.N_33 ));
    InMux I__2464 (
            .O(N__10867),
            .I(N__10864));
    LocalMux I__2463 (
            .O(N__10864),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER21_NE_0_0 ));
    InMux I__2462 (
            .O(N__10861),
            .I(N__10855));
    CascadeMux I__2461 (
            .O(N__10860),
            .I(N__10852));
    InMux I__2460 (
            .O(N__10859),
            .I(N__10845));
    InMux I__2459 (
            .O(N__10858),
            .I(N__10842));
    LocalMux I__2458 (
            .O(N__10855),
            .I(N__10839));
    InMux I__2457 (
            .O(N__10852),
            .I(N__10834));
    InMux I__2456 (
            .O(N__10851),
            .I(N__10834));
    InMux I__2455 (
            .O(N__10850),
            .I(N__10829));
    InMux I__2454 (
            .O(N__10849),
            .I(N__10829));
    InMux I__2453 (
            .O(N__10848),
            .I(N__10826));
    LocalMux I__2452 (
            .O(N__10845),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__2451 (
            .O(N__10842),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    Odrv4 I__2450 (
            .O(N__10839),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__2449 (
            .O(N__10834),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__2448 (
            .O(N__10829),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__2447 (
            .O(N__10826),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    InMux I__2446 (
            .O(N__10813),
            .I(N__10809));
    InMux I__2445 (
            .O(N__10812),
            .I(N__10802));
    LocalMux I__2444 (
            .O(N__10809),
            .I(N__10799));
    CascadeMux I__2443 (
            .O(N__10808),
            .I(N__10796));
    InMux I__2442 (
            .O(N__10807),
            .I(N__10792));
    InMux I__2441 (
            .O(N__10806),
            .I(N__10789));
    InMux I__2440 (
            .O(N__10805),
            .I(N__10786));
    LocalMux I__2439 (
            .O(N__10802),
            .I(N__10783));
    Span4Mux_h I__2438 (
            .O(N__10799),
            .I(N__10780));
    InMux I__2437 (
            .O(N__10796),
            .I(N__10777));
    InMux I__2436 (
            .O(N__10795),
            .I(N__10774));
    LocalMux I__2435 (
            .O(N__10792),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__2434 (
            .O(N__10789),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__2433 (
            .O(N__10786),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    Odrv4 I__2432 (
            .O(N__10783),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    Odrv4 I__2431 (
            .O(N__10780),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__2430 (
            .O(N__10777),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__2429 (
            .O(N__10774),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    InMux I__2428 (
            .O(N__10759),
            .I(N__10751));
    InMux I__2427 (
            .O(N__10758),
            .I(N__10748));
    InMux I__2426 (
            .O(N__10757),
            .I(N__10745));
    InMux I__2425 (
            .O(N__10756),
            .I(N__10742));
    InMux I__2424 (
            .O(N__10755),
            .I(N__10737));
    InMux I__2423 (
            .O(N__10754),
            .I(N__10737));
    LocalMux I__2422 (
            .O(N__10751),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__2421 (
            .O(N__10748),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__2420 (
            .O(N__10745),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__2419 (
            .O(N__10742),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__2418 (
            .O(N__10737),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    CascadeMux I__2417 (
            .O(N__10726),
            .I(N__10723));
    InMux I__2416 (
            .O(N__10723),
            .I(N__10720));
    LocalMux I__2415 (
            .O(N__10720),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER22_NE_0_0 ));
    CascadeMux I__2414 (
            .O(N__10717),
            .I(N__10712));
    CascadeMux I__2413 (
            .O(N__10716),
            .I(N__10709));
    InMux I__2412 (
            .O(N__10715),
            .I(N__10704));
    InMux I__2411 (
            .O(N__10712),
            .I(N__10701));
    InMux I__2410 (
            .O(N__10709),
            .I(N__10698));
    InMux I__2409 (
            .O(N__10708),
            .I(N__10695));
    InMux I__2408 (
            .O(N__10707),
            .I(N__10692));
    LocalMux I__2407 (
            .O(N__10704),
            .I(N__10687));
    LocalMux I__2406 (
            .O(N__10701),
            .I(N__10687));
    LocalMux I__2405 (
            .O(N__10698),
            .I(N__10682));
    LocalMux I__2404 (
            .O(N__10695),
            .I(N__10682));
    LocalMux I__2403 (
            .O(N__10692),
            .I(N__10679));
    Span4Mux_v I__2402 (
            .O(N__10687),
            .I(N__10676));
    Span4Mux_v I__2401 (
            .O(N__10682),
            .I(N__10673));
    Span12Mux_v I__2400 (
            .O(N__10679),
            .I(N__10668));
    Sp12to4 I__2399 (
            .O(N__10676),
            .I(N__10668));
    Sp12to4 I__2398 (
            .O(N__10673),
            .I(N__10665));
    Span12Mux_h I__2397 (
            .O(N__10668),
            .I(N__10662));
    Span12Mux_h I__2396 (
            .O(N__10665),
            .I(N__10659));
    Span12Mux_v I__2395 (
            .O(N__10662),
            .I(N__10656));
    Span12Mux_v I__2394 (
            .O(N__10659),
            .I(N__10653));
    Odrv12 I__2393 (
            .O(N__10656),
            .I(ROM_DELAY_c_0));
    Odrv12 I__2392 (
            .O(N__10653),
            .I(ROM_DELAY_c_0));
    InMux I__2391 (
            .O(N__10648),
            .I(N__10641));
    InMux I__2390 (
            .O(N__10647),
            .I(N__10641));
    InMux I__2389 (
            .O(N__10646),
            .I(N__10638));
    LocalMux I__2388 (
            .O(N__10641),
            .I(N__10632));
    LocalMux I__2387 (
            .O(N__10638),
            .I(N__10632));
    InMux I__2386 (
            .O(N__10637),
            .I(N__10629));
    Span4Mux_h I__2385 (
            .O(N__10632),
            .I(N__10623));
    LocalMux I__2384 (
            .O(N__10629),
            .I(N__10623));
    InMux I__2383 (
            .O(N__10628),
            .I(N__10620));
    Span4Mux_h I__2382 (
            .O(N__10623),
            .I(N__10615));
    LocalMux I__2381 (
            .O(N__10620),
            .I(N__10615));
    Sp12to4 I__2380 (
            .O(N__10615),
            .I(N__10612));
    Span12Mux_v I__2379 (
            .O(N__10612),
            .I(N__10609));
    Span12Mux_h I__2378 (
            .O(N__10609),
            .I(N__10606));
    Odrv12 I__2377 (
            .O(N__10606),
            .I(ROM_DELAY_c_1));
    CascadeMux I__2376 (
            .O(N__10603),
            .I(N__10599));
    InMux I__2375 (
            .O(N__10602),
            .I(N__10596));
    InMux I__2374 (
            .O(N__10599),
            .I(N__10593));
    LocalMux I__2373 (
            .O(N__10596),
            .I(\U409_TRANSFER_ACK.N_31_i ));
    LocalMux I__2372 (
            .O(N__10593),
            .I(\U409_TRANSFER_ACK.N_31_i ));
    InMux I__2371 (
            .O(N__10588),
            .I(N__10585));
    LocalMux I__2370 (
            .O(N__10585),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ));
    InMux I__2369 (
            .O(N__10582),
            .I(\U409_TICK.un3_COUNTER60_1_cry_7 ));
    InMux I__2368 (
            .O(N__10579),
            .I(bfn_14_7_0_));
    InMux I__2367 (
            .O(N__10576),
            .I(\U409_TICK.un3_COUNTER60_1_cry_9 ));
    InMux I__2366 (
            .O(N__10573),
            .I(\U409_TICK.un3_COUNTER60_1_cry_10 ));
    InMux I__2365 (
            .O(N__10570),
            .I(\U409_TICK.un3_COUNTER60_1_cry_11 ));
    InMux I__2364 (
            .O(N__10567),
            .I(\U409_TICK.un3_COUNTER60_1_cry_12 ));
    InMux I__2363 (
            .O(N__10564),
            .I(\U409_TICK.un3_COUNTER60_1_cry_13 ));
    InMux I__2362 (
            .O(N__10561),
            .I(\U409_TICK.un3_COUNTER60_1_cry_14 ));
    InMux I__2361 (
            .O(N__10558),
            .I(\U409_TICK.un3_COUNTER60_1_cry_15 ));
    IoInMux I__2360 (
            .O(N__10555),
            .I(N__10552));
    LocalMux I__2359 (
            .O(N__10552),
            .I(N__10549));
    IoSpan4Mux I__2358 (
            .O(N__10549),
            .I(N__10546));
    Sp12to4 I__2357 (
            .O(N__10546),
            .I(N__10543));
    Span12Mux_s7_v I__2356 (
            .O(N__10543),
            .I(N__10540));
    Span12Mux_v I__2355 (
            .O(N__10540),
            .I(N__10537));
    Odrv12 I__2354 (
            .O(N__10537),
            .I(PCIAT_c_1));
    InMux I__2353 (
            .O(N__10534),
            .I(N__10530));
    InMux I__2352 (
            .O(N__10533),
            .I(N__10527));
    LocalMux I__2351 (
            .O(N__10530),
            .I(N__10522));
    LocalMux I__2350 (
            .O(N__10527),
            .I(N__10522));
    Span4Mux_v I__2349 (
            .O(N__10522),
            .I(N__10519));
    Sp12to4 I__2348 (
            .O(N__10519),
            .I(N__10516));
    Span12Mux_h I__2347 (
            .O(N__10516),
            .I(N__10513));
    Odrv12 I__2346 (
            .O(N__10513),
            .I(TM_c_0));
    InMux I__2345 (
            .O(N__10510),
            .I(N__10506));
    InMux I__2344 (
            .O(N__10509),
            .I(N__10503));
    LocalMux I__2343 (
            .O(N__10506),
            .I(N__10498));
    LocalMux I__2342 (
            .O(N__10503),
            .I(N__10498));
    Span4Mux_v I__2341 (
            .O(N__10498),
            .I(N__10495));
    Sp12to4 I__2340 (
            .O(N__10495),
            .I(N__10492));
    Odrv12 I__2339 (
            .O(N__10492),
            .I(\U409_ADDRESS_DECODE.N_58_mux ));
    InMux I__2338 (
            .O(N__10489),
            .I(N__10486));
    LocalMux I__2337 (
            .O(N__10486),
            .I(N__10483));
    Span4Mux_v I__2336 (
            .O(N__10483),
            .I(N__10479));
    InMux I__2335 (
            .O(N__10482),
            .I(N__10476));
    Sp12to4 I__2334 (
            .O(N__10479),
            .I(N__10471));
    LocalMux I__2333 (
            .O(N__10476),
            .I(N__10471));
    Span12Mux_h I__2332 (
            .O(N__10471),
            .I(N__10468));
    Odrv12 I__2331 (
            .O(N__10468),
            .I(TM_c_1));
    IoInMux I__2330 (
            .O(N__10465),
            .I(N__10462));
    LocalMux I__2329 (
            .O(N__10462),
            .I(N__10459));
    Span4Mux_s3_h I__2328 (
            .O(N__10459),
            .I(N__10456));
    Sp12to4 I__2327 (
            .O(N__10456),
            .I(N__10453));
    Span12Mux_s11_v I__2326 (
            .O(N__10453),
            .I(N__10450));
    Span12Mux_h I__2325 (
            .O(N__10450),
            .I(N__10447));
    Odrv12 I__2324 (
            .O(N__10447),
            .I(PCIAT_c_0));
    InMux I__2323 (
            .O(N__10444),
            .I(\U409_TICK.un3_COUNTER60_1_cry_1 ));
    InMux I__2322 (
            .O(N__10441),
            .I(\U409_TICK.un3_COUNTER60_1_cry_2 ));
    InMux I__2321 (
            .O(N__10438),
            .I(\U409_TICK.un3_COUNTER60_1_cry_3 ));
    InMux I__2320 (
            .O(N__10435),
            .I(\U409_TICK.un3_COUNTER60_1_cry_4 ));
    InMux I__2319 (
            .O(N__10432),
            .I(\U409_TICK.un3_COUNTER60_1_cry_5 ));
    InMux I__2318 (
            .O(N__10429),
            .I(\U409_TICK.un3_COUNTER60_1_cry_6 ));
    InMux I__2317 (
            .O(N__10426),
            .I(N__10420));
    InMux I__2316 (
            .O(N__10425),
            .I(N__10420));
    LocalMux I__2315 (
            .O(N__10420),
            .I(N__10417));
    Span4Mux_v I__2314 (
            .O(N__10417),
            .I(N__10414));
    Span4Mux_h I__2313 (
            .O(N__10414),
            .I(N__10411));
    Odrv4 I__2312 (
            .O(N__10411),
            .I(\U409_TRANSFER_ACK.un1_AUTOVECTOR_0 ));
    CascadeMux I__2311 (
            .O(N__10408),
            .I(N__10404));
    CascadeMux I__2310 (
            .O(N__10407),
            .I(N__10401));
    InMux I__2309 (
            .O(N__10404),
            .I(N__10396));
    InMux I__2308 (
            .O(N__10401),
            .I(N__10396));
    LocalMux I__2307 (
            .O(N__10396),
            .I(N__10391));
    InMux I__2306 (
            .O(N__10395),
            .I(N__10388));
    InMux I__2305 (
            .O(N__10394),
            .I(N__10385));
    Span4Mux_v I__2304 (
            .O(N__10391),
            .I(N__10382));
    LocalMux I__2303 (
            .O(N__10388),
            .I(N__10379));
    LocalMux I__2302 (
            .O(N__10385),
            .I(N__10376));
    Span4Mux_v I__2301 (
            .O(N__10382),
            .I(N__10373));
    Span4Mux_v I__2300 (
            .O(N__10379),
            .I(N__10370));
    Span4Mux_v I__2299 (
            .O(N__10376),
            .I(N__10367));
    Sp12to4 I__2298 (
            .O(N__10373),
            .I(N__10362));
    Sp12to4 I__2297 (
            .O(N__10370),
            .I(N__10362));
    Span4Mux_h I__2296 (
            .O(N__10367),
            .I(N__10359));
    Span12Mux_h I__2295 (
            .O(N__10362),
            .I(N__10354));
    Sp12to4 I__2294 (
            .O(N__10359),
            .I(N__10354));
    Span12Mux_v I__2293 (
            .O(N__10354),
            .I(N__10351));
    Odrv12 I__2292 (
            .O(N__10351),
            .I(TSn_c));
    InMux I__2291 (
            .O(N__10348),
            .I(N__10344));
    InMux I__2290 (
            .O(N__10347),
            .I(N__10341));
    LocalMux I__2289 (
            .O(N__10344),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    LocalMux I__2288 (
            .O(N__10341),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    CascadeMux I__2287 (
            .O(N__10336),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1_cascade_ ));
    InMux I__2286 (
            .O(N__10333),
            .I(N__10329));
    InMux I__2285 (
            .O(N__10332),
            .I(N__10326));
    LocalMux I__2284 (
            .O(N__10329),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    LocalMux I__2283 (
            .O(N__10326),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    InMux I__2282 (
            .O(N__10321),
            .I(N__10318));
    LocalMux I__2281 (
            .O(N__10318),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER22_NE_1_0 ));
    InMux I__2280 (
            .O(N__10315),
            .I(N__10311));
    InMux I__2279 (
            .O(N__10314),
            .I(N__10308));
    LocalMux I__2278 (
            .O(N__10311),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    LocalMux I__2277 (
            .O(N__10308),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    CascadeMux I__2276 (
            .O(N__10303),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_NE_1_0_cascade_ ));
    CascadeMux I__2275 (
            .O(N__10300),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0_cascade_ ));
    InMux I__2274 (
            .O(N__10297),
            .I(N__10294));
    LocalMux I__2273 (
            .O(N__10294),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0_0 ));
    IoInMux I__2272 (
            .O(N__10291),
            .I(N__10288));
    LocalMux I__2271 (
            .O(N__10288),
            .I(N__10285));
    IoSpan4Mux I__2270 (
            .O(N__10285),
            .I(N__10282));
    Span4Mux_s2_v I__2269 (
            .O(N__10282),
            .I(N__10279));
    Span4Mux_v I__2268 (
            .O(N__10279),
            .I(N__10276));
    Sp12to4 I__2267 (
            .O(N__10276),
            .I(N__10272));
    InMux I__2266 (
            .O(N__10275),
            .I(N__10269));
    Odrv12 I__2265 (
            .O(N__10272),
            .I(ROMENn_c));
    LocalMux I__2264 (
            .O(N__10269),
            .I(ROMENn_c));
    InMux I__2263 (
            .O(N__10264),
            .I(N__10261));
    LocalMux I__2262 (
            .O(N__10261),
            .I(\U409_TRANSFER_ACK.N_42_i ));
    InMux I__2261 (
            .O(N__10258),
            .I(N__10255));
    LocalMux I__2260 (
            .O(N__10255),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER21_0 ));
    InMux I__2259 (
            .O(N__10252),
            .I(N__10249));
    LocalMux I__2258 (
            .O(N__10249),
            .I(N__10246));
    Span4Mux_h I__2257 (
            .O(N__10246),
            .I(N__10242));
    InMux I__2256 (
            .O(N__10245),
            .I(N__10239));
    Odrv4 I__2255 (
            .O(N__10242),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENn_2 ));
    LocalMux I__2254 (
            .O(N__10239),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENn_2 ));
    CascadeMux I__2253 (
            .O(N__10234),
            .I(N__10231));
    InMux I__2252 (
            .O(N__10231),
            .I(N__10228));
    LocalMux I__2251 (
            .O(N__10228),
            .I(N__10225));
    Odrv4 I__2250 (
            .O(N__10225),
            .I(\U409_ADDRESS_DECODE.N_61 ));
    CascadeMux I__2249 (
            .O(N__10222),
            .I(\U409_TRANSFER_ACK.N_42_i_cascade_ ));
    CascadeMux I__2248 (
            .O(N__10219),
            .I(N__10215));
    CascadeMux I__2247 (
            .O(N__10218),
            .I(N__10210));
    InMux I__2246 (
            .O(N__10215),
            .I(N__10206));
    InMux I__2245 (
            .O(N__10214),
            .I(N__10203));
    InMux I__2244 (
            .O(N__10213),
            .I(N__10198));
    InMux I__2243 (
            .O(N__10210),
            .I(N__10198));
    InMux I__2242 (
            .O(N__10209),
            .I(N__10195));
    LocalMux I__2241 (
            .O(N__10206),
            .I(N__10191));
    LocalMux I__2240 (
            .O(N__10203),
            .I(N__10187));
    LocalMux I__2239 (
            .O(N__10198),
            .I(N__10184));
    LocalMux I__2238 (
            .O(N__10195),
            .I(N__10181));
    InMux I__2237 (
            .O(N__10194),
            .I(N__10178));
    Span4Mux_v I__2236 (
            .O(N__10191),
            .I(N__10175));
    InMux I__2235 (
            .O(N__10190),
            .I(N__10171));
    Span4Mux_v I__2234 (
            .O(N__10187),
            .I(N__10168));
    Span4Mux_h I__2233 (
            .O(N__10184),
            .I(N__10163));
    Span4Mux_v I__2232 (
            .O(N__10181),
            .I(N__10163));
    LocalMux I__2231 (
            .O(N__10178),
            .I(N__10160));
    Span4Mux_h I__2230 (
            .O(N__10175),
            .I(N__10157));
    InMux I__2229 (
            .O(N__10174),
            .I(N__10154));
    LocalMux I__2228 (
            .O(N__10171),
            .I(N__10151));
    Span4Mux_v I__2227 (
            .O(N__10168),
            .I(N__10148));
    Span4Mux_h I__2226 (
            .O(N__10163),
            .I(N__10143));
    Span4Mux_v I__2225 (
            .O(N__10160),
            .I(N__10143));
    Span4Mux_h I__2224 (
            .O(N__10157),
            .I(N__10138));
    LocalMux I__2223 (
            .O(N__10154),
            .I(N__10138));
    Span12Mux_v I__2222 (
            .O(N__10151),
            .I(N__10135));
    Sp12to4 I__2221 (
            .O(N__10148),
            .I(N__10132));
    Span4Mux_v I__2220 (
            .O(N__10143),
            .I(N__10129));
    Sp12to4 I__2219 (
            .O(N__10138),
            .I(N__10126));
    Span12Mux_h I__2218 (
            .O(N__10135),
            .I(N__10123));
    Span12Mux_h I__2217 (
            .O(N__10132),
            .I(N__10116));
    Sp12to4 I__2216 (
            .O(N__10129),
            .I(N__10116));
    Span12Mux_v I__2215 (
            .O(N__10126),
            .I(N__10116));
    Odrv12 I__2214 (
            .O(N__10123),
            .I(A_c_23));
    Odrv12 I__2213 (
            .O(N__10116),
            .I(A_c_23));
    InMux I__2212 (
            .O(N__10111),
            .I(N__10104));
    InMux I__2211 (
            .O(N__10110),
            .I(N__10101));
    InMux I__2210 (
            .O(N__10109),
            .I(N__10097));
    InMux I__2209 (
            .O(N__10108),
            .I(N__10094));
    InMux I__2208 (
            .O(N__10107),
            .I(N__10091));
    LocalMux I__2207 (
            .O(N__10104),
            .I(N__10085));
    LocalMux I__2206 (
            .O(N__10101),
            .I(N__10085));
    InMux I__2205 (
            .O(N__10100),
            .I(N__10082));
    LocalMux I__2204 (
            .O(N__10097),
            .I(N__10079));
    LocalMux I__2203 (
            .O(N__10094),
            .I(N__10074));
    LocalMux I__2202 (
            .O(N__10091),
            .I(N__10074));
    InMux I__2201 (
            .O(N__10090),
            .I(N__10071));
    Span4Mux_v I__2200 (
            .O(N__10085),
            .I(N__10068));
    LocalMux I__2199 (
            .O(N__10082),
            .I(N__10065));
    Span4Mux_v I__2198 (
            .O(N__10079),
            .I(N__10062));
    Span4Mux_v I__2197 (
            .O(N__10074),
            .I(N__10057));
    LocalMux I__2196 (
            .O(N__10071),
            .I(N__10057));
    Span4Mux_v I__2195 (
            .O(N__10068),
            .I(N__10054));
    Span4Mux_v I__2194 (
            .O(N__10065),
            .I(N__10051));
    Span4Mux_h I__2193 (
            .O(N__10062),
            .I(N__10046));
    Span4Mux_v I__2192 (
            .O(N__10057),
            .I(N__10046));
    Span4Mux_h I__2191 (
            .O(N__10054),
            .I(N__10042));
    Span4Mux_v I__2190 (
            .O(N__10051),
            .I(N__10037));
    Span4Mux_h I__2189 (
            .O(N__10046),
            .I(N__10037));
    InMux I__2188 (
            .O(N__10045),
            .I(N__10034));
    Sp12to4 I__2187 (
            .O(N__10042),
            .I(N__10027));
    Sp12to4 I__2186 (
            .O(N__10037),
            .I(N__10027));
    LocalMux I__2185 (
            .O(N__10034),
            .I(N__10027));
    Odrv12 I__2184 (
            .O(N__10027),
            .I(A_c_20));
    InMux I__2183 (
            .O(N__10024),
            .I(N__10021));
    LocalMux I__2182 (
            .O(N__10021),
            .I(\U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_1 ));
    CascadeMux I__2181 (
            .O(N__10018),
            .I(N__10013));
    InMux I__2180 (
            .O(N__10017),
            .I(N__10006));
    InMux I__2179 (
            .O(N__10016),
            .I(N__10002));
    InMux I__2178 (
            .O(N__10013),
            .I(N__9999));
    InMux I__2177 (
            .O(N__10012),
            .I(N__9996));
    InMux I__2176 (
            .O(N__10011),
            .I(N__9993));
    CascadeMux I__2175 (
            .O(N__10010),
            .I(N__9990));
    CascadeMux I__2174 (
            .O(N__10009),
            .I(N__9987));
    LocalMux I__2173 (
            .O(N__10006),
            .I(N__9984));
    CascadeMux I__2172 (
            .O(N__10005),
            .I(N__9981));
    LocalMux I__2171 (
            .O(N__10002),
            .I(N__9978));
    LocalMux I__2170 (
            .O(N__9999),
            .I(N__9975));
    LocalMux I__2169 (
            .O(N__9996),
            .I(N__9969));
    LocalMux I__2168 (
            .O(N__9993),
            .I(N__9969));
    InMux I__2167 (
            .O(N__9990),
            .I(N__9966));
    InMux I__2166 (
            .O(N__9987),
            .I(N__9963));
    Span4Mux_v I__2165 (
            .O(N__9984),
            .I(N__9960));
    InMux I__2164 (
            .O(N__9981),
            .I(N__9957));
    Span4Mux_v I__2163 (
            .O(N__9978),
            .I(N__9954));
    Span4Mux_v I__2162 (
            .O(N__9975),
            .I(N__9951));
    InMux I__2161 (
            .O(N__9974),
            .I(N__9948));
    Span12Mux_v I__2160 (
            .O(N__9969),
            .I(N__9943));
    LocalMux I__2159 (
            .O(N__9966),
            .I(N__9943));
    LocalMux I__2158 (
            .O(N__9963),
            .I(N__9930));
    Sp12to4 I__2157 (
            .O(N__9960),
            .I(N__9930));
    LocalMux I__2156 (
            .O(N__9957),
            .I(N__9930));
    Sp12to4 I__2155 (
            .O(N__9954),
            .I(N__9930));
    Sp12to4 I__2154 (
            .O(N__9951),
            .I(N__9930));
    LocalMux I__2153 (
            .O(N__9948),
            .I(N__9930));
    Span12Mux_v I__2152 (
            .O(N__9943),
            .I(N__9927));
    Span12Mux_h I__2151 (
            .O(N__9930),
            .I(N__9924));
    Span12Mux_h I__2150 (
            .O(N__9927),
            .I(N__9919));
    Span12Mux_v I__2149 (
            .O(N__9924),
            .I(N__9919));
    Odrv12 I__2148 (
            .O(N__9919),
            .I(A_c_19));
    InMux I__2147 (
            .O(N__9916),
            .I(N__9909));
    InMux I__2146 (
            .O(N__9915),
            .I(N__9906));
    InMux I__2145 (
            .O(N__9914),
            .I(N__9903));
    InMux I__2144 (
            .O(N__9913),
            .I(N__9900));
    InMux I__2143 (
            .O(N__9912),
            .I(N__9896));
    LocalMux I__2142 (
            .O(N__9909),
            .I(N__9892));
    LocalMux I__2141 (
            .O(N__9906),
            .I(N__9889));
    LocalMux I__2140 (
            .O(N__9903),
            .I(N__9886));
    LocalMux I__2139 (
            .O(N__9900),
            .I(N__9883));
    InMux I__2138 (
            .O(N__9899),
            .I(N__9880));
    LocalMux I__2137 (
            .O(N__9896),
            .I(N__9877));
    InMux I__2136 (
            .O(N__9895),
            .I(N__9874));
    Span4Mux_v I__2135 (
            .O(N__9892),
            .I(N__9871));
    Span4Mux_v I__2134 (
            .O(N__9889),
            .I(N__9868));
    Span4Mux_v I__2133 (
            .O(N__9886),
            .I(N__9864));
    Span4Mux_v I__2132 (
            .O(N__9883),
            .I(N__9861));
    LocalMux I__2131 (
            .O(N__9880),
            .I(N__9854));
    Span4Mux_h I__2130 (
            .O(N__9877),
            .I(N__9854));
    LocalMux I__2129 (
            .O(N__9874),
            .I(N__9854));
    Span4Mux_v I__2128 (
            .O(N__9871),
            .I(N__9851));
    Span4Mux_v I__2127 (
            .O(N__9868),
            .I(N__9848));
    InMux I__2126 (
            .O(N__9867),
            .I(N__9845));
    Sp12to4 I__2125 (
            .O(N__9864),
            .I(N__9840));
    Sp12to4 I__2124 (
            .O(N__9861),
            .I(N__9840));
    Sp12to4 I__2123 (
            .O(N__9854),
            .I(N__9837));
    Span4Mux_v I__2122 (
            .O(N__9851),
            .I(N__9834));
    Span4Mux_v I__2121 (
            .O(N__9848),
            .I(N__9831));
    LocalMux I__2120 (
            .O(N__9845),
            .I(N__9828));
    Span12Mux_h I__2119 (
            .O(N__9840),
            .I(N__9825));
    Span12Mux_v I__2118 (
            .O(N__9837),
            .I(N__9822));
    Sp12to4 I__2117 (
            .O(N__9834),
            .I(N__9819));
    Span4Mux_v I__2116 (
            .O(N__9831),
            .I(N__9816));
    Sp12to4 I__2115 (
            .O(N__9828),
            .I(N__9813));
    Span12Mux_v I__2114 (
            .O(N__9825),
            .I(N__9808));
    Span12Mux_h I__2113 (
            .O(N__9822),
            .I(N__9808));
    Span12Mux_h I__2112 (
            .O(N__9819),
            .I(N__9801));
    Sp12to4 I__2111 (
            .O(N__9816),
            .I(N__9801));
    Span12Mux_v I__2110 (
            .O(N__9813),
            .I(N__9801));
    Odrv12 I__2109 (
            .O(N__9808),
            .I(A_c_22));
    Odrv12 I__2108 (
            .O(N__9801),
            .I(A_c_22));
    InMux I__2107 (
            .O(N__9796),
            .I(N__9792));
    CascadeMux I__2106 (
            .O(N__9795),
            .I(N__9789));
    LocalMux I__2105 (
            .O(N__9792),
            .I(N__9786));
    InMux I__2104 (
            .O(N__9789),
            .I(N__9782));
    Span4Mux_v I__2103 (
            .O(N__9786),
            .I(N__9779));
    InMux I__2102 (
            .O(N__9785),
            .I(N__9776));
    LocalMux I__2101 (
            .O(N__9782),
            .I(N__9769));
    Sp12to4 I__2100 (
            .O(N__9779),
            .I(N__9769));
    LocalMux I__2099 (
            .O(N__9776),
            .I(N__9769));
    Span12Mux_v I__2098 (
            .O(N__9769),
            .I(N__9766));
    Span12Mux_h I__2097 (
            .O(N__9766),
            .I(N__9763));
    Odrv12 I__2096 (
            .O(N__9763),
            .I(OVL_c));
    CascadeMux I__2095 (
            .O(N__9760),
            .I(N__9755));
    InMux I__2094 (
            .O(N__9759),
            .I(N__9751));
    InMux I__2093 (
            .O(N__9758),
            .I(N__9748));
    InMux I__2092 (
            .O(N__9755),
            .I(N__9745));
    CascadeMux I__2091 (
            .O(N__9754),
            .I(N__9741));
    LocalMux I__2090 (
            .O(N__9751),
            .I(N__9733));
    LocalMux I__2089 (
            .O(N__9748),
            .I(N__9733));
    LocalMux I__2088 (
            .O(N__9745),
            .I(N__9733));
    InMux I__2087 (
            .O(N__9744),
            .I(N__9730));
    InMux I__2086 (
            .O(N__9741),
            .I(N__9725));
    InMux I__2085 (
            .O(N__9740),
            .I(N__9720));
    Span4Mux_h I__2084 (
            .O(N__9733),
            .I(N__9715));
    LocalMux I__2083 (
            .O(N__9730),
            .I(N__9715));
    InMux I__2082 (
            .O(N__9729),
            .I(N__9712));
    InMux I__2081 (
            .O(N__9728),
            .I(N__9709));
    LocalMux I__2080 (
            .O(N__9725),
            .I(N__9705));
    InMux I__2079 (
            .O(N__9724),
            .I(N__9702));
    InMux I__2078 (
            .O(N__9723),
            .I(N__9699));
    LocalMux I__2077 (
            .O(N__9720),
            .I(N__9695));
    Span4Mux_h I__2076 (
            .O(N__9715),
            .I(N__9690));
    LocalMux I__2075 (
            .O(N__9712),
            .I(N__9690));
    LocalMux I__2074 (
            .O(N__9709),
            .I(N__9687));
    InMux I__2073 (
            .O(N__9708),
            .I(N__9684));
    Span4Mux_v I__2072 (
            .O(N__9705),
            .I(N__9676));
    LocalMux I__2071 (
            .O(N__9702),
            .I(N__9676));
    LocalMux I__2070 (
            .O(N__9699),
            .I(N__9676));
    InMux I__2069 (
            .O(N__9698),
            .I(N__9673));
    Span4Mux_h I__2068 (
            .O(N__9695),
            .I(N__9668));
    Span4Mux_v I__2067 (
            .O(N__9690),
            .I(N__9668));
    Span4Mux_v I__2066 (
            .O(N__9687),
            .I(N__9665));
    LocalMux I__2065 (
            .O(N__9684),
            .I(N__9662));
    InMux I__2064 (
            .O(N__9683),
            .I(N__9659));
    Span4Mux_v I__2063 (
            .O(N__9676),
            .I(N__9656));
    LocalMux I__2062 (
            .O(N__9673),
            .I(N__9653));
    Span4Mux_v I__2061 (
            .O(N__9668),
            .I(N__9646));
    Span4Mux_h I__2060 (
            .O(N__9665),
            .I(N__9646));
    Span4Mux_v I__2059 (
            .O(N__9662),
            .I(N__9646));
    LocalMux I__2058 (
            .O(N__9659),
            .I(N__9643));
    Span4Mux_h I__2057 (
            .O(N__9656),
            .I(N__9640));
    Sp12to4 I__2056 (
            .O(N__9653),
            .I(N__9637));
    Span4Mux_h I__2055 (
            .O(N__9646),
            .I(N__9632));
    Span4Mux_v I__2054 (
            .O(N__9643),
            .I(N__9632));
    Sp12to4 I__2053 (
            .O(N__9640),
            .I(N__9625));
    Span12Mux_v I__2052 (
            .O(N__9637),
            .I(N__9625));
    Sp12to4 I__2051 (
            .O(N__9632),
            .I(N__9625));
    Odrv12 I__2050 (
            .O(N__9625),
            .I(A_c_21));
    InMux I__2049 (
            .O(N__9622),
            .I(N__9619));
    LocalMux I__2048 (
            .O(N__9619),
            .I(\U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_2 ));
    InMux I__2047 (
            .O(N__9616),
            .I(N__9613));
    LocalMux I__2046 (
            .O(N__9613),
            .I(N__9610));
    Odrv12 I__2045 (
            .O(N__9610),
            .I(ROMEN));
    IoInMux I__2044 (
            .O(N__9607),
            .I(N__9604));
    LocalMux I__2043 (
            .O(N__9604),
            .I(N__9600));
    IoInMux I__2042 (
            .O(N__9603),
            .I(N__9597));
    Span12Mux_s5_v I__2041 (
            .O(N__9600),
            .I(N__9594));
    LocalMux I__2040 (
            .O(N__9597),
            .I(N__9591));
    Span12Mux_v I__2039 (
            .O(N__9594),
            .I(N__9586));
    Span12Mux_s10_v I__2038 (
            .O(N__9591),
            .I(N__9583));
    InMux I__2037 (
            .O(N__9590),
            .I(N__9580));
    CascadeMux I__2036 (
            .O(N__9589),
            .I(N__9577));
    Span12Mux_h I__2035 (
            .O(N__9586),
            .I(N__9574));
    Span12Mux_h I__2034 (
            .O(N__9583),
            .I(N__9569));
    LocalMux I__2033 (
            .O(N__9580),
            .I(N__9569));
    InMux I__2032 (
            .O(N__9577),
            .I(N__9566));
    Odrv12 I__2031 (
            .O(N__9574),
            .I(TACK_EN));
    Odrv12 I__2030 (
            .O(N__9569),
            .I(TACK_EN));
    LocalMux I__2029 (
            .O(N__9566),
            .I(TACK_EN));
    IoInMux I__2028 (
            .O(N__9559),
            .I(N__9556));
    LocalMux I__2027 (
            .O(N__9556),
            .I(N__9553));
    Span4Mux_s1_v I__2026 (
            .O(N__9553),
            .I(N__9550));
    Sp12to4 I__2025 (
            .O(N__9550),
            .I(N__9547));
    Span12Mux_s9_h I__2024 (
            .O(N__9547),
            .I(N__9544));
    Span12Mux_v I__2023 (
            .O(N__9544),
            .I(N__9541));
    Odrv12 I__2022 (
            .O(N__9541),
            .I(TCIn_1_i));
    IoInMux I__2021 (
            .O(N__9538),
            .I(N__9535));
    LocalMux I__2020 (
            .O(N__9535),
            .I(N__9532));
    Odrv12 I__2019 (
            .O(N__9532),
            .I(RESETn_c_i));
    InMux I__2018 (
            .O(N__9529),
            .I(N__9526));
    LocalMux I__2017 (
            .O(N__9526),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    InMux I__2016 (
            .O(N__9523),
            .I(N__9519));
    InMux I__2015 (
            .O(N__9522),
            .I(N__9516));
    LocalMux I__2014 (
            .O(N__9519),
            .I(N__9513));
    LocalMux I__2013 (
            .O(N__9516),
            .I(AC_TACK));
    Odrv4 I__2012 (
            .O(N__9513),
            .I(AC_TACK));
    CascadeMux I__2011 (
            .O(N__9508),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_ ));
    CascadeMux I__2010 (
            .O(N__9505),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ));
    CascadeMux I__2009 (
            .O(N__9502),
            .I(\U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ));
    IoInMux I__2008 (
            .O(N__9499),
            .I(N__9495));
    IoInMux I__2007 (
            .O(N__9498),
            .I(N__9492));
    LocalMux I__2006 (
            .O(N__9495),
            .I(N__9486));
    LocalMux I__2005 (
            .O(N__9492),
            .I(N__9486));
    IoInMux I__2004 (
            .O(N__9491),
            .I(N__9483));
    Span12Mux_s6_v I__2003 (
            .O(N__9486),
            .I(N__9480));
    LocalMux I__2002 (
            .O(N__9483),
            .I(N__9477));
    Span12Mux_v I__2001 (
            .O(N__9480),
            .I(N__9474));
    Span12Mux_s11_v I__2000 (
            .O(N__9477),
            .I(N__9471));
    Span12Mux_h I__1999 (
            .O(N__9474),
            .I(N__9466));
    Span12Mux_h I__1998 (
            .O(N__9471),
            .I(N__9463));
    InMux I__1997 (
            .O(N__9470),
            .I(N__9458));
    InMux I__1996 (
            .O(N__9469),
            .I(N__9458));
    Odrv12 I__1995 (
            .O(N__9466),
            .I(TACK_OUTn));
    Odrv12 I__1994 (
            .O(N__9463),
            .I(TACK_OUTn));
    LocalMux I__1993 (
            .O(N__9458),
            .I(TACK_OUTn));
    InMux I__1992 (
            .O(N__9451),
            .I(N__9445));
    InMux I__1991 (
            .O(N__9450),
            .I(N__9438));
    InMux I__1990 (
            .O(N__9449),
            .I(N__9438));
    InMux I__1989 (
            .O(N__9448),
            .I(N__9438));
    LocalMux I__1988 (
            .O(N__9445),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    LocalMux I__1987 (
            .O(N__9438),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    InMux I__1986 (
            .O(N__9433),
            .I(N__9427));
    InMux I__1985 (
            .O(N__9432),
            .I(N__9420));
    InMux I__1984 (
            .O(N__9431),
            .I(N__9420));
    InMux I__1983 (
            .O(N__9430),
            .I(N__9420));
    LocalMux I__1982 (
            .O(N__9427),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    LocalMux I__1981 (
            .O(N__9420),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    InMux I__1980 (
            .O(N__9415),
            .I(N__9411));
    InMux I__1979 (
            .O(N__9414),
            .I(N__9408));
    LocalMux I__1978 (
            .O(N__9411),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    LocalMux I__1977 (
            .O(N__9408),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    InMux I__1976 (
            .O(N__9403),
            .I(N__9400));
    LocalMux I__1975 (
            .O(N__9400),
            .I(N__9392));
    InMux I__1974 (
            .O(N__9399),
            .I(N__9389));
    InMux I__1973 (
            .O(N__9398),
            .I(N__9385));
    InMux I__1972 (
            .O(N__9397),
            .I(N__9382));
    InMux I__1971 (
            .O(N__9396),
            .I(N__9379));
    InMux I__1970 (
            .O(N__9395),
            .I(N__9376));
    Span4Mux_v I__1969 (
            .O(N__9392),
            .I(N__9370));
    LocalMux I__1968 (
            .O(N__9389),
            .I(N__9370));
    InMux I__1967 (
            .O(N__9388),
            .I(N__9367));
    LocalMux I__1966 (
            .O(N__9385),
            .I(N__9364));
    LocalMux I__1965 (
            .O(N__9382),
            .I(N__9359));
    LocalMux I__1964 (
            .O(N__9379),
            .I(N__9359));
    LocalMux I__1963 (
            .O(N__9376),
            .I(N__9356));
    InMux I__1962 (
            .O(N__9375),
            .I(N__9353));
    Span4Mux_h I__1961 (
            .O(N__9370),
            .I(N__9347));
    LocalMux I__1960 (
            .O(N__9367),
            .I(N__9347));
    Span4Mux_v I__1959 (
            .O(N__9364),
            .I(N__9340));
    Span4Mux_h I__1958 (
            .O(N__9359),
            .I(N__9340));
    Span4Mux_v I__1957 (
            .O(N__9356),
            .I(N__9340));
    LocalMux I__1956 (
            .O(N__9353),
            .I(N__9337));
    InMux I__1955 (
            .O(N__9352),
            .I(N__9334));
    Span4Mux_v I__1954 (
            .O(N__9347),
            .I(N__9331));
    Span4Mux_h I__1953 (
            .O(N__9340),
            .I(N__9324));
    Span4Mux_v I__1952 (
            .O(N__9337),
            .I(N__9324));
    LocalMux I__1951 (
            .O(N__9334),
            .I(N__9324));
    Sp12to4 I__1950 (
            .O(N__9331),
            .I(N__9321));
    Span4Mux_h I__1949 (
            .O(N__9324),
            .I(N__9318));
    Span12Mux_h I__1948 (
            .O(N__9321),
            .I(N__9315));
    Span4Mux_v I__1947 (
            .O(N__9318),
            .I(N__9312));
    Odrv12 I__1946 (
            .O(N__9315),
            .I(\U409_ADDRESS_DECODE.Z2_SPACE ));
    Odrv4 I__1945 (
            .O(N__9312),
            .I(\U409_ADDRESS_DECODE.Z2_SPACE ));
    CascadeMux I__1944 (
            .O(N__9307),
            .I(ROMEN_cascade_));
    CascadeMux I__1943 (
            .O(N__9304),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0_cascade_ ));
    CascadeMux I__1942 (
            .O(N__9301),
            .I(N__9298));
    InMux I__1941 (
            .O(N__9298),
            .I(N__9293));
    InMux I__1940 (
            .O(N__9297),
            .I(N__9288));
    InMux I__1939 (
            .O(N__9296),
            .I(N__9288));
    LocalMux I__1938 (
            .O(N__9293),
            .I(N__9285));
    LocalMux I__1937 (
            .O(N__9288),
            .I(N__9280));
    Span4Mux_v I__1936 (
            .O(N__9285),
            .I(N__9277));
    InMux I__1935 (
            .O(N__9284),
            .I(N__9274));
    CascadeMux I__1934 (
            .O(N__9283),
            .I(N__9271));
    Span4Mux_h I__1933 (
            .O(N__9280),
            .I(N__9268));
    Span4Mux_h I__1932 (
            .O(N__9277),
            .I(N__9263));
    LocalMux I__1931 (
            .O(N__9274),
            .I(N__9263));
    InMux I__1930 (
            .O(N__9271),
            .I(N__9260));
    Span4Mux_h I__1929 (
            .O(N__9268),
            .I(N__9255));
    Span4Mux_v I__1928 (
            .O(N__9263),
            .I(N__9255));
    LocalMux I__1927 (
            .O(N__9260),
            .I(N__9252));
    Span4Mux_v I__1926 (
            .O(N__9255),
            .I(N__9249));
    Sp12to4 I__1925 (
            .O(N__9252),
            .I(N__9246));
    Sp12to4 I__1924 (
            .O(N__9249),
            .I(N__9241));
    Span12Mux_v I__1923 (
            .O(N__9246),
            .I(N__9241));
    Odrv12 I__1922 (
            .O(N__9241),
            .I(A_c_16));
    InMux I__1921 (
            .O(N__9238),
            .I(N__9232));
    InMux I__1920 (
            .O(N__9237),
            .I(N__9232));
    LocalMux I__1919 (
            .O(N__9232),
            .I(N__9229));
    Span4Mux_v I__1918 (
            .O(N__9229),
            .I(N__9226));
    Sp12to4 I__1917 (
            .O(N__9226),
            .I(N__9223));
    Span12Mux_h I__1916 (
            .O(N__9223),
            .I(N__9220));
    Odrv12 I__1915 (
            .O(N__9220),
            .I(A_c_15));
    InMux I__1914 (
            .O(N__9217),
            .I(N__9212));
    CascadeMux I__1913 (
            .O(N__9216),
            .I(N__9209));
    CascadeMux I__1912 (
            .O(N__9215),
            .I(N__9206));
    LocalMux I__1911 (
            .O(N__9212),
            .I(N__9203));
    InMux I__1910 (
            .O(N__9209),
            .I(N__9198));
    InMux I__1909 (
            .O(N__9206),
            .I(N__9198));
    Span4Mux_v I__1908 (
            .O(N__9203),
            .I(N__9193));
    LocalMux I__1907 (
            .O(N__9198),
            .I(N__9193));
    Span4Mux_v I__1906 (
            .O(N__9193),
            .I(N__9190));
    Sp12to4 I__1905 (
            .O(N__9190),
            .I(N__9187));
    Span12Mux_h I__1904 (
            .O(N__9187),
            .I(N__9184));
    Odrv12 I__1903 (
            .O(N__9184),
            .I(A_c_13));
    IoInMux I__1902 (
            .O(N__9181),
            .I(N__9178));
    LocalMux I__1901 (
            .O(N__9178),
            .I(N__9175));
    IoSpan4Mux I__1900 (
            .O(N__9175),
            .I(N__9172));
    Span4Mux_s2_h I__1899 (
            .O(N__9172),
            .I(N__9169));
    Sp12to4 I__1898 (
            .O(N__9169),
            .I(N__9166));
    Span12Mux_h I__1897 (
            .O(N__9166),
            .I(N__9163));
    Odrv12 I__1896 (
            .O(N__9163),
            .I(U409_ADDRESS_DECODE_un1_CIACS1n_i));
    InMux I__1895 (
            .O(N__9160),
            .I(N__9157));
    LocalMux I__1894 (
            .O(N__9157),
            .I(CIA_ENABLE));
    CascadeMux I__1893 (
            .O(N__9154),
            .I(CIA_ENABLE_cascade_));
    InMux I__1892 (
            .O(N__9151),
            .I(N__9145));
    InMux I__1891 (
            .O(N__9150),
            .I(N__9145));
    LocalMux I__1890 (
            .O(N__9145),
            .I(N__9142));
    Span4Mux_v I__1889 (
            .O(N__9142),
            .I(N__9138));
    InMux I__1888 (
            .O(N__9141),
            .I(N__9135));
    Sp12to4 I__1887 (
            .O(N__9138),
            .I(N__9130));
    LocalMux I__1886 (
            .O(N__9135),
            .I(N__9130));
    Span12Mux_h I__1885 (
            .O(N__9130),
            .I(N__9127));
    Odrv12 I__1884 (
            .O(N__9127),
            .I(A_c_12));
    IoInMux I__1883 (
            .O(N__9124),
            .I(N__9121));
    LocalMux I__1882 (
            .O(N__9121),
            .I(N__9118));
    IoSpan4Mux I__1881 (
            .O(N__9118),
            .I(N__9115));
    IoSpan4Mux I__1880 (
            .O(N__9115),
            .I(N__9112));
    Span4Mux_s3_h I__1879 (
            .O(N__9112),
            .I(N__9109));
    Span4Mux_h I__1878 (
            .O(N__9109),
            .I(N__9106));
    Sp12to4 I__1877 (
            .O(N__9106),
            .I(N__9103));
    Odrv12 I__1876 (
            .O(N__9103),
            .I(U409_ADDRESS_DECODE_un1_CIACS0n_i));
    CascadeMux I__1875 (
            .O(N__9100),
            .I(N__9097));
    InMux I__1874 (
            .O(N__9097),
            .I(N__9093));
    InMux I__1873 (
            .O(N__9096),
            .I(N__9089));
    LocalMux I__1872 (
            .O(N__9093),
            .I(N__9086));
    InMux I__1871 (
            .O(N__9092),
            .I(N__9083));
    LocalMux I__1870 (
            .O(N__9089),
            .I(N__9079));
    Span4Mux_v I__1869 (
            .O(N__9086),
            .I(N__9076));
    LocalMux I__1868 (
            .O(N__9083),
            .I(N__9073));
    InMux I__1867 (
            .O(N__9082),
            .I(N__9070));
    Span12Mux_v I__1866 (
            .O(N__9079),
            .I(N__9067));
    Span4Mux_h I__1865 (
            .O(N__9076),
            .I(N__9064));
    Span4Mux_v I__1864 (
            .O(N__9073),
            .I(N__9061));
    LocalMux I__1863 (
            .O(N__9070),
            .I(N__9058));
    Odrv12 I__1862 (
            .O(N__9067),
            .I(\U409_ADDRESS_DECODE.N_75 ));
    Odrv4 I__1861 (
            .O(N__9064),
            .I(\U409_ADDRESS_DECODE.N_75 ));
    Odrv4 I__1860 (
            .O(N__9061),
            .I(\U409_ADDRESS_DECODE.N_75 ));
    Odrv4 I__1859 (
            .O(N__9058),
            .I(\U409_ADDRESS_DECODE.N_75 ));
    IoInMux I__1858 (
            .O(N__9049),
            .I(N__9046));
    LocalMux I__1857 (
            .O(N__9046),
            .I(N__9043));
    Span4Mux_s3_h I__1856 (
            .O(N__9043),
            .I(N__9040));
    Span4Mux_v I__1855 (
            .O(N__9040),
            .I(N__9037));
    Span4Mux_h I__1854 (
            .O(N__9037),
            .I(N__9034));
    Span4Mux_h I__1853 (
            .O(N__9034),
            .I(N__9031));
    Span4Mux_h I__1852 (
            .O(N__9031),
            .I(N__9028));
    Odrv4 I__1851 (
            .O(N__9028),
            .I(N_77_mux_i));
    CascadeMux I__1850 (
            .O(N__9025),
            .I(N__9022));
    InMux I__1849 (
            .O(N__9022),
            .I(N__9019));
    LocalMux I__1848 (
            .O(N__9019),
            .I(N__9015));
    InMux I__1847 (
            .O(N__9018),
            .I(N__9012));
    Span4Mux_v I__1846 (
            .O(N__9015),
            .I(N__9009));
    LocalMux I__1845 (
            .O(N__9012),
            .I(N__9006));
    Odrv4 I__1844 (
            .O(N__9009),
            .I(\U409_ADDRESS_DECODE.N_60_1 ));
    Odrv4 I__1843 (
            .O(N__9006),
            .I(\U409_ADDRESS_DECODE.N_60_1 ));
    IoInMux I__1842 (
            .O(N__9001),
            .I(N__8998));
    LocalMux I__1841 (
            .O(N__8998),
            .I(N__8995));
    Span12Mux_s11_v I__1840 (
            .O(N__8995),
            .I(N__8992));
    Odrv12 I__1839 (
            .O(N__8992),
            .I(U409_ADDRESS_DECODE_un1_RAMSPACEn_i));
    InMux I__1838 (
            .O(N__8989),
            .I(N__8986));
    LocalMux I__1837 (
            .O(N__8986),
            .I(N__8983));
    Odrv4 I__1836 (
            .O(N__8983),
            .I(\U409_AUTOCONFIG.STATE4 ));
    InMux I__1835 (
            .O(N__8980),
            .I(N__8973));
    InMux I__1834 (
            .O(N__8979),
            .I(N__8968));
    InMux I__1833 (
            .O(N__8978),
            .I(N__8968));
    InMux I__1832 (
            .O(N__8977),
            .I(N__8965));
    InMux I__1831 (
            .O(N__8976),
            .I(N__8962));
    LocalMux I__1830 (
            .O(N__8973),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_6));
    LocalMux I__1829 (
            .O(N__8968),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_6));
    LocalMux I__1828 (
            .O(N__8965),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_6));
    LocalMux I__1827 (
            .O(N__8962),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_6));
    CascadeMux I__1826 (
            .O(N__8953),
            .I(N__8950));
    InMux I__1825 (
            .O(N__8950),
            .I(N__8947));
    LocalMux I__1824 (
            .O(N__8947),
            .I(N_71_mux));
    InMux I__1823 (
            .O(N__8944),
            .I(N__8939));
    InMux I__1822 (
            .O(N__8943),
            .I(N__8936));
    InMux I__1821 (
            .O(N__8942),
            .I(N__8933));
    LocalMux I__1820 (
            .O(N__8939),
            .I(N_70_mux));
    LocalMux I__1819 (
            .O(N__8936),
            .I(N_70_mux));
    LocalMux I__1818 (
            .O(N__8933),
            .I(N_70_mux));
    CEMux I__1817 (
            .O(N__8926),
            .I(N__8923));
    LocalMux I__1816 (
            .O(N__8923),
            .I(\U409_TRANSFER_ACK.N_20_0 ));
    InMux I__1815 (
            .O(N__8920),
            .I(N__8916));
    InMux I__1814 (
            .O(N__8919),
            .I(N__8913));
    LocalMux I__1813 (
            .O(N__8916),
            .I(N__8910));
    LocalMux I__1812 (
            .O(N__8913),
            .I(\U409_AUTOCONFIG.STATE_d_2 ));
    Odrv4 I__1811 (
            .O(N__8910),
            .I(\U409_AUTOCONFIG.STATE_d_2 ));
    InMux I__1810 (
            .O(N__8905),
            .I(N__8899));
    InMux I__1809 (
            .O(N__8904),
            .I(N__8896));
    CascadeMux I__1808 (
            .O(N__8903),
            .I(N__8892));
    InMux I__1807 (
            .O(N__8902),
            .I(N__8888));
    LocalMux I__1806 (
            .O(N__8899),
            .I(N__8883));
    LocalMux I__1805 (
            .O(N__8896),
            .I(N__8883));
    InMux I__1804 (
            .O(N__8895),
            .I(N__8876));
    InMux I__1803 (
            .O(N__8892),
            .I(N__8876));
    InMux I__1802 (
            .O(N__8891),
            .I(N__8876));
    LocalMux I__1801 (
            .O(N__8888),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    Odrv12 I__1800 (
            .O(N__8883),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    LocalMux I__1799 (
            .O(N__8876),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    CascadeMux I__1798 (
            .O(N__8869),
            .I(N__8863));
    InMux I__1797 (
            .O(N__8868),
            .I(N__8860));
    InMux I__1796 (
            .O(N__8867),
            .I(N__8857));
    InMux I__1795 (
            .O(N__8866),
            .I(N__8853));
    InMux I__1794 (
            .O(N__8863),
            .I(N__8850));
    LocalMux I__1793 (
            .O(N__8860),
            .I(N__8847));
    LocalMux I__1792 (
            .O(N__8857),
            .I(N__8844));
    InMux I__1791 (
            .O(N__8856),
            .I(N__8841));
    LocalMux I__1790 (
            .O(N__8853),
            .I(N__8838));
    LocalMux I__1789 (
            .O(N__8850),
            .I(N__8834));
    Span4Mux_v I__1788 (
            .O(N__8847),
            .I(N__8831));
    Span4Mux_v I__1787 (
            .O(N__8844),
            .I(N__8826));
    LocalMux I__1786 (
            .O(N__8841),
            .I(N__8826));
    Span4Mux_v I__1785 (
            .O(N__8838),
            .I(N__8823));
    InMux I__1784 (
            .O(N__8837),
            .I(N__8820));
    Span4Mux_v I__1783 (
            .O(N__8834),
            .I(N__8817));
    Span4Mux_v I__1782 (
            .O(N__8831),
            .I(N__8814));
    Span4Mux_v I__1781 (
            .O(N__8826),
            .I(N__8811));
    Sp12to4 I__1780 (
            .O(N__8823),
            .I(N__8806));
    LocalMux I__1779 (
            .O(N__8820),
            .I(N__8806));
    Sp12to4 I__1778 (
            .O(N__8817),
            .I(N__8799));
    Sp12to4 I__1777 (
            .O(N__8814),
            .I(N__8799));
    Sp12to4 I__1776 (
            .O(N__8811),
            .I(N__8799));
    Span12Mux_h I__1775 (
            .O(N__8806),
            .I(N__8796));
    Span12Mux_h I__1774 (
            .O(N__8799),
            .I(N__8793));
    Span12Mux_v I__1773 (
            .O(N__8796),
            .I(N__8790));
    Span12Mux_v I__1772 (
            .O(N__8793),
            .I(N__8787));
    Odrv12 I__1771 (
            .O(N__8790),
            .I(RnW_c));
    Odrv12 I__1770 (
            .O(N__8787),
            .I(RnW_c));
    InMux I__1769 (
            .O(N__8782),
            .I(N__8779));
    LocalMux I__1768 (
            .O(N__8779),
            .I(N__8774));
    InMux I__1767 (
            .O(N__8778),
            .I(N__8771));
    InMux I__1766 (
            .O(N__8777),
            .I(N__8765));
    Span4Mux_h I__1765 (
            .O(N__8774),
            .I(N__8762));
    LocalMux I__1764 (
            .O(N__8771),
            .I(N__8759));
    InMux I__1763 (
            .O(N__8770),
            .I(N__8752));
    InMux I__1762 (
            .O(N__8769),
            .I(N__8752));
    InMux I__1761 (
            .O(N__8768),
            .I(N__8752));
    LocalMux I__1760 (
            .O(N__8765),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    Odrv4 I__1759 (
            .O(N__8762),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    Odrv12 I__1758 (
            .O(N__8759),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    LocalMux I__1757 (
            .O(N__8752),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    CascadeMux I__1756 (
            .O(N__8743),
            .I(N__8739));
    InMux I__1755 (
            .O(N__8742),
            .I(N__8736));
    InMux I__1754 (
            .O(N__8739),
            .I(N__8733));
    LocalMux I__1753 (
            .O(N__8736),
            .I(N__8730));
    LocalMux I__1752 (
            .O(N__8733),
            .I(N__8727));
    Span4Mux_v I__1751 (
            .O(N__8730),
            .I(N__8723));
    Span4Mux_v I__1750 (
            .O(N__8727),
            .I(N__8720));
    InMux I__1749 (
            .O(N__8726),
            .I(N__8717));
    Odrv4 I__1748 (
            .O(N__8723),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn));
    Odrv4 I__1747 (
            .O(N__8720),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn));
    LocalMux I__1746 (
            .O(N__8717),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn));
    InMux I__1745 (
            .O(N__8710),
            .I(N__8707));
    LocalMux I__1744 (
            .O(N__8707),
            .I(N__8704));
    Sp12to4 I__1743 (
            .O(N__8704),
            .I(N__8701));
    Span12Mux_v I__1742 (
            .O(N__8701),
            .I(N__8698));
    Span12Mux_h I__1741 (
            .O(N__8698),
            .I(N__8695));
    Odrv12 I__1740 (
            .O(N__8695),
            .I(TACKn_in));
    CascadeMux I__1739 (
            .O(N__8692),
            .I(N__8689));
    InMux I__1738 (
            .O(N__8689),
            .I(N__8685));
    InMux I__1737 (
            .O(N__8688),
            .I(N__8682));
    LocalMux I__1736 (
            .O(N__8685),
            .I(N__8677));
    LocalMux I__1735 (
            .O(N__8682),
            .I(N__8677));
    Odrv12 I__1734 (
            .O(N__8677),
            .I(U409_ADDRESS_DECODE_un1_RAMSPACEn));
    SRMux I__1733 (
            .O(N__8674),
            .I(N__8670));
    SRMux I__1732 (
            .O(N__8673),
            .I(N__8667));
    LocalMux I__1731 (
            .O(N__8670),
            .I(N__8663));
    LocalMux I__1730 (
            .O(N__8667),
            .I(N__8660));
    SRMux I__1729 (
            .O(N__8666),
            .I(N__8657));
    Span4Mux_v I__1728 (
            .O(N__8663),
            .I(N__8651));
    Span4Mux_h I__1727 (
            .O(N__8660),
            .I(N__8651));
    LocalMux I__1726 (
            .O(N__8657),
            .I(N__8648));
    SRMux I__1725 (
            .O(N__8656),
            .I(N__8645));
    Odrv4 I__1724 (
            .O(N__8651),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    Odrv4 I__1723 (
            .O(N__8648),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    LocalMux I__1722 (
            .O(N__8645),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    IoInMux I__1721 (
            .O(N__8638),
            .I(N__8635));
    LocalMux I__1720 (
            .O(N__8635),
            .I(N__8632));
    Span4Mux_s2_v I__1719 (
            .O(N__8632),
            .I(N__8629));
    Span4Mux_v I__1718 (
            .O(N__8629),
            .I(N__8626));
    Odrv4 I__1717 (
            .O(N__8626),
            .I(GB_BUFFER_CLK40_IN_c_g_THRU_CO));
    CascadeMux I__1716 (
            .O(N__8623),
            .I(N__8616));
    InMux I__1715 (
            .O(N__8622),
            .I(N__8609));
    InMux I__1714 (
            .O(N__8621),
            .I(N__8609));
    InMux I__1713 (
            .O(N__8620),
            .I(N__8609));
    InMux I__1712 (
            .O(N__8619),
            .I(N__8604));
    InMux I__1711 (
            .O(N__8616),
            .I(N__8604));
    LocalMux I__1710 (
            .O(N__8609),
            .I(N_23));
    LocalMux I__1709 (
            .O(N__8604),
            .I(N_23));
    CascadeMux I__1708 (
            .O(N__8599),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ));
    CascadeMux I__1707 (
            .O(N__8596),
            .I(N__8592));
    CascadeMux I__1706 (
            .O(N__8595),
            .I(N__8587));
    InMux I__1705 (
            .O(N__8592),
            .I(N__8579));
    InMux I__1704 (
            .O(N__8591),
            .I(N__8579));
    InMux I__1703 (
            .O(N__8590),
            .I(N__8579));
    InMux I__1702 (
            .O(N__8587),
            .I(N__8574));
    InMux I__1701 (
            .O(N__8586),
            .I(N__8574));
    LocalMux I__1700 (
            .O(N__8579),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_3));
    LocalMux I__1699 (
            .O(N__8574),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_3));
    InMux I__1698 (
            .O(N__8569),
            .I(N__8560));
    InMux I__1697 (
            .O(N__8568),
            .I(N__8560));
    InMux I__1696 (
            .O(N__8567),
            .I(N__8553));
    InMux I__1695 (
            .O(N__8566),
            .I(N__8553));
    InMux I__1694 (
            .O(N__8565),
            .I(N__8553));
    LocalMux I__1693 (
            .O(N__8560),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_0));
    LocalMux I__1692 (
            .O(N__8553),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_0));
    InMux I__1691 (
            .O(N__8548),
            .I(N__8545));
    LocalMux I__1690 (
            .O(N__8545),
            .I(N__8539));
    InMux I__1689 (
            .O(N__8544),
            .I(N__8536));
    InMux I__1688 (
            .O(N__8543),
            .I(N__8533));
    InMux I__1687 (
            .O(N__8542),
            .I(N__8529));
    Span4Mux_h I__1686 (
            .O(N__8539),
            .I(N__8524));
    LocalMux I__1685 (
            .O(N__8536),
            .I(N__8524));
    LocalMux I__1684 (
            .O(N__8533),
            .I(N__8521));
    InMux I__1683 (
            .O(N__8532),
            .I(N__8518));
    LocalMux I__1682 (
            .O(N__8529),
            .I(N__8515));
    Span4Mux_v I__1681 (
            .O(N__8524),
            .I(N__8508));
    Span4Mux_v I__1680 (
            .O(N__8521),
            .I(N__8508));
    LocalMux I__1679 (
            .O(N__8518),
            .I(N__8508));
    Odrv12 I__1678 (
            .O(N__8515),
            .I(\U409_ADDRESS_DECODE.CIA_SPACE_4 ));
    Odrv4 I__1677 (
            .O(N__8508),
            .I(\U409_ADDRESS_DECODE.CIA_SPACE_4 ));
    CascadeMux I__1676 (
            .O(N__8503),
            .I(N__8500));
    InMux I__1675 (
            .O(N__8500),
            .I(N__8497));
    LocalMux I__1674 (
            .O(N__8497),
            .I(N__8492));
    InMux I__1673 (
            .O(N__8496),
            .I(N__8489));
    CascadeMux I__1672 (
            .O(N__8495),
            .I(N__8486));
    Span4Mux_v I__1671 (
            .O(N__8492),
            .I(N__8481));
    LocalMux I__1670 (
            .O(N__8489),
            .I(N__8481));
    InMux I__1669 (
            .O(N__8486),
            .I(N__8478));
    Span4Mux_h I__1668 (
            .O(N__8481),
            .I(N__8474));
    LocalMux I__1667 (
            .O(N__8478),
            .I(N__8471));
    InMux I__1666 (
            .O(N__8477),
            .I(N__8468));
    Span4Mux_v I__1665 (
            .O(N__8474),
            .I(N__8463));
    Span4Mux_v I__1664 (
            .O(N__8471),
            .I(N__8463));
    LocalMux I__1663 (
            .O(N__8468),
            .I(N__8460));
    Odrv4 I__1662 (
            .O(N__8463),
            .I(\U409_ADDRESS_DECODE.CIA_SPACE_5 ));
    Odrv12 I__1661 (
            .O(N__8460),
            .I(\U409_ADDRESS_DECODE.CIA_SPACE_5 ));
    InMux I__1660 (
            .O(N__8455),
            .I(N__8451));
    InMux I__1659 (
            .O(N__8454),
            .I(N__8448));
    LocalMux I__1658 (
            .O(N__8451),
            .I(LIDE_BASE_4));
    LocalMux I__1657 (
            .O(N__8448),
            .I(LIDE_BASE_4));
    CascadeMux I__1656 (
            .O(N__8443),
            .I(N__8440));
    InMux I__1655 (
            .O(N__8440),
            .I(N__8436));
    InMux I__1654 (
            .O(N__8439),
            .I(N__8433));
    LocalMux I__1653 (
            .O(N__8436),
            .I(LIDE_BASE_3));
    LocalMux I__1652 (
            .O(N__8433),
            .I(LIDE_BASE_3));
    InMux I__1651 (
            .O(N__8428),
            .I(N__8425));
    LocalMux I__1650 (
            .O(N__8425),
            .I(\U409_ADDRESS_DECODE.ATA_SPACE_1Z0Z_0 ));
    InMux I__1649 (
            .O(N__8422),
            .I(N__8418));
    InMux I__1648 (
            .O(N__8421),
            .I(N__8414));
    LocalMux I__1647 (
            .O(N__8418),
            .I(N__8410));
    InMux I__1646 (
            .O(N__8417),
            .I(N__8407));
    LocalMux I__1645 (
            .O(N__8414),
            .I(N__8404));
    InMux I__1644 (
            .O(N__8413),
            .I(N__8401));
    Span4Mux_v I__1643 (
            .O(N__8410),
            .I(N__8398));
    LocalMux I__1642 (
            .O(N__8407),
            .I(N__8391));
    Span4Mux_v I__1641 (
            .O(N__8404),
            .I(N__8391));
    LocalMux I__1640 (
            .O(N__8401),
            .I(N__8391));
    Span4Mux_h I__1639 (
            .O(N__8398),
            .I(N__8385));
    Span4Mux_v I__1638 (
            .O(N__8391),
            .I(N__8385));
    InMux I__1637 (
            .O(N__8390),
            .I(N__8382));
    Odrv4 I__1636 (
            .O(N__8385),
            .I(AUTOCONFIG_SPACE));
    LocalMux I__1635 (
            .O(N__8382),
            .I(AUTOCONFIG_SPACE));
    IoInMux I__1634 (
            .O(N__8377),
            .I(N__8374));
    LocalMux I__1633 (
            .O(N__8374),
            .I(N__8371));
    Span12Mux_s7_v I__1632 (
            .O(N__8371),
            .I(N__8368));
    Span12Mux_v I__1631 (
            .O(N__8368),
            .I(N__8365));
    Odrv12 I__1630 (
            .O(N__8365),
            .I(BUFENn_c));
    CascadeMux I__1629 (
            .O(N__8362),
            .I(N__8359));
    InMux I__1628 (
            .O(N__8359),
            .I(N__8352));
    InMux I__1627 (
            .O(N__8358),
            .I(N__8352));
    InMux I__1626 (
            .O(N__8357),
            .I(N__8349));
    LocalMux I__1625 (
            .O(N__8352),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0 ));
    LocalMux I__1624 (
            .O(N__8349),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0 ));
    InMux I__1623 (
            .O(N__8344),
            .I(N__8339));
    InMux I__1622 (
            .O(N__8343),
            .I(N__8334));
    InMux I__1621 (
            .O(N__8342),
            .I(N__8334));
    LocalMux I__1620 (
            .O(N__8339),
            .I(\U409_ADDRESS_DECODE.ATA_ENZ0 ));
    LocalMux I__1619 (
            .O(N__8334),
            .I(\U409_ADDRESS_DECODE.ATA_ENZ0 ));
    IoInMux I__1618 (
            .O(N__8329),
            .I(N__8326));
    LocalMux I__1617 (
            .O(N__8326),
            .I(N__8323));
    IoSpan4Mux I__1616 (
            .O(N__8323),
            .I(N__8320));
    Sp12to4 I__1615 (
            .O(N__8320),
            .I(N__8317));
    Span12Mux_s7_h I__1614 (
            .O(N__8317),
            .I(N__8314));
    Odrv12 I__1613 (
            .O(N__8314),
            .I(U409_ADDRESS_DECODE_un1_ATA_ENn_i));
    CascadeMux I__1612 (
            .O(N__8311),
            .I(N__8305));
    InMux I__1611 (
            .O(N__8310),
            .I(N__8302));
    InMux I__1610 (
            .O(N__8309),
            .I(N__8299));
    InMux I__1609 (
            .O(N__8308),
            .I(N__8294));
    InMux I__1608 (
            .O(N__8305),
            .I(N__8294));
    LocalMux I__1607 (
            .O(N__8302),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_7));
    LocalMux I__1606 (
            .O(N__8299),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_7));
    LocalMux I__1605 (
            .O(N__8294),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_7));
    CascadeMux I__1604 (
            .O(N__8287),
            .I(\U409_ADDRESS_DECODE.m27Z0Z_3_cascade_ ));
    InMux I__1603 (
            .O(N__8284),
            .I(N__8278));
    InMux I__1602 (
            .O(N__8283),
            .I(N__8278));
    LocalMux I__1601 (
            .O(N__8278),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ));
    CascadeMux I__1600 (
            .O(N__8275),
            .I(N__8270));
    InMux I__1599 (
            .O(N__8274),
            .I(N__8264));
    InMux I__1598 (
            .O(N__8273),
            .I(N__8264));
    InMux I__1597 (
            .O(N__8270),
            .I(N__8259));
    InMux I__1596 (
            .O(N__8269),
            .I(N__8259));
    LocalMux I__1595 (
            .O(N__8264),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_4));
    LocalMux I__1594 (
            .O(N__8259),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_4));
    InMux I__1593 (
            .O(N__8254),
            .I(N__8251));
    LocalMux I__1592 (
            .O(N__8251),
            .I(U409_ADDRESS_DECODE_m33_1));
    CascadeMux I__1591 (
            .O(N__8248),
            .I(U409_ADDRESS_DECODE_m33_1_cascade_));
    InMux I__1590 (
            .O(N__8245),
            .I(N__8239));
    InMux I__1589 (
            .O(N__8244),
            .I(N__8236));
    InMux I__1588 (
            .O(N__8243),
            .I(N__8231));
    InMux I__1587 (
            .O(N__8242),
            .I(N__8231));
    LocalMux I__1586 (
            .O(N__8239),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_5));
    LocalMux I__1585 (
            .O(N__8236),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_5));
    LocalMux I__1584 (
            .O(N__8231),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_5));
    InMux I__1583 (
            .O(N__8224),
            .I(N__8218));
    InMux I__1582 (
            .O(N__8223),
            .I(N__8211));
    InMux I__1581 (
            .O(N__8222),
            .I(N__8211));
    InMux I__1580 (
            .O(N__8221),
            .I(N__8211));
    LocalMux I__1579 (
            .O(N__8218),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_1));
    LocalMux I__1578 (
            .O(N__8211),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_1));
    CascadeMux I__1577 (
            .O(N__8206),
            .I(N__8202));
    InMux I__1576 (
            .O(N__8205),
            .I(N__8199));
    InMux I__1575 (
            .O(N__8202),
            .I(N__8196));
    LocalMux I__1574 (
            .O(N__8199),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c2 ));
    LocalMux I__1573 (
            .O(N__8196),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c2 ));
    InMux I__1572 (
            .O(N__8191),
            .I(N__8184));
    InMux I__1571 (
            .O(N__8190),
            .I(N__8181));
    InMux I__1570 (
            .O(N__8189),
            .I(N__8178));
    InMux I__1569 (
            .O(N__8188),
            .I(N__8173));
    InMux I__1568 (
            .O(N__8187),
            .I(N__8173));
    LocalMux I__1567 (
            .O(N__8184),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_2));
    LocalMux I__1566 (
            .O(N__8181),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_2));
    LocalMux I__1565 (
            .O(N__8178),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_2));
    LocalMux I__1564 (
            .O(N__8173),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_2));
    CascadeMux I__1563 (
            .O(N__8164),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c2_cascade_ ));
    InMux I__1562 (
            .O(N__8161),
            .I(N__8155));
    InMux I__1561 (
            .O(N__8160),
            .I(N__8155));
    LocalMux I__1560 (
            .O(N__8155),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ));
    CascadeMux I__1559 (
            .O(N__8152),
            .I(N__8149));
    InMux I__1558 (
            .O(N__8149),
            .I(N__8144));
    InMux I__1557 (
            .O(N__8148),
            .I(N__8139));
    InMux I__1556 (
            .O(N__8147),
            .I(N__8139));
    LocalMux I__1555 (
            .O(N__8144),
            .I(N__8134));
    LocalMux I__1554 (
            .O(N__8139),
            .I(N__8131));
    CascadeMux I__1553 (
            .O(N__8138),
            .I(N__8128));
    CascadeMux I__1552 (
            .O(N__8137),
            .I(N__8125));
    Span4Mux_v I__1551 (
            .O(N__8134),
            .I(N__8120));
    Span4Mux_v I__1550 (
            .O(N__8131),
            .I(N__8120));
    InMux I__1549 (
            .O(N__8128),
            .I(N__8115));
    InMux I__1548 (
            .O(N__8125),
            .I(N__8115));
    Sp12to4 I__1547 (
            .O(N__8120),
            .I(N__8110));
    LocalMux I__1546 (
            .O(N__8115),
            .I(N__8110));
    Span12Mux_h I__1545 (
            .O(N__8110),
            .I(N__8107));
    Span12Mux_v I__1544 (
            .O(N__8107),
            .I(N__8104));
    Odrv12 I__1543 (
            .O(N__8104),
            .I(D_in_5));
    InMux I__1542 (
            .O(N__8101),
            .I(N__8098));
    LocalMux I__1541 (
            .O(N__8098),
            .I(N__8094));
    CascadeMux I__1540 (
            .O(N__8097),
            .I(N__8091));
    Span4Mux_v I__1539 (
            .O(N__8094),
            .I(N__8088));
    InMux I__1538 (
            .O(N__8091),
            .I(N__8085));
    Odrv4 I__1537 (
            .O(N__8088),
            .I(BRIDGE_BASE_1));
    LocalMux I__1536 (
            .O(N__8085),
            .I(BRIDGE_BASE_1));
    CascadeMux I__1535 (
            .O(N__8080),
            .I(N__8077));
    InMux I__1534 (
            .O(N__8077),
            .I(N__8073));
    InMux I__1533 (
            .O(N__8076),
            .I(N__8070));
    LocalMux I__1532 (
            .O(N__8073),
            .I(N__8067));
    LocalMux I__1531 (
            .O(N__8070),
            .I(LIDE_BASE_7));
    Odrv12 I__1530 (
            .O(N__8067),
            .I(LIDE_BASE_7));
    CascadeMux I__1529 (
            .O(N__8062),
            .I(N__8058));
    CascadeMux I__1528 (
            .O(N__8061),
            .I(N__8055));
    InMux I__1527 (
            .O(N__8058),
            .I(N__8052));
    InMux I__1526 (
            .O(N__8055),
            .I(N__8049));
    LocalMux I__1525 (
            .O(N__8052),
            .I(N__8043));
    LocalMux I__1524 (
            .O(N__8049),
            .I(N__8040));
    InMux I__1523 (
            .O(N__8048),
            .I(N__8033));
    InMux I__1522 (
            .O(N__8047),
            .I(N__8033));
    InMux I__1521 (
            .O(N__8046),
            .I(N__8033));
    Span4Mux_v I__1520 (
            .O(N__8043),
            .I(N__8030));
    Span4Mux_h I__1519 (
            .O(N__8040),
            .I(N__8025));
    LocalMux I__1518 (
            .O(N__8033),
            .I(N__8025));
    Span4Mux_h I__1517 (
            .O(N__8030),
            .I(N__8020));
    Span4Mux_v I__1516 (
            .O(N__8025),
            .I(N__8020));
    Sp12to4 I__1515 (
            .O(N__8020),
            .I(N__8017));
    Odrv12 I__1514 (
            .O(N__8017),
            .I(D_in_7));
    InMux I__1513 (
            .O(N__8014),
            .I(N__8008));
    InMux I__1512 (
            .O(N__8013),
            .I(N__8003));
    InMux I__1511 (
            .O(N__8012),
            .I(N__8003));
    InMux I__1510 (
            .O(N__8011),
            .I(N__8000));
    LocalMux I__1509 (
            .O(N__8008),
            .I(\U409_AUTOCONFIG.BRIDGE_CONF_RNID7FUZ0Z1 ));
    LocalMux I__1508 (
            .O(N__8003),
            .I(\U409_AUTOCONFIG.BRIDGE_CONF_RNID7FUZ0Z1 ));
    LocalMux I__1507 (
            .O(N__8000),
            .I(\U409_AUTOCONFIG.BRIDGE_CONF_RNID7FUZ0Z1 ));
    CascadeMux I__1506 (
            .O(N__7993),
            .I(N__7990));
    InMux I__1505 (
            .O(N__7990),
            .I(N__7986));
    CascadeMux I__1504 (
            .O(N__7989),
            .I(N__7983));
    LocalMux I__1503 (
            .O(N__7986),
            .I(N__7980));
    InMux I__1502 (
            .O(N__7983),
            .I(N__7977));
    Odrv4 I__1501 (
            .O(N__7980),
            .I(BRIDGE_BASE_3));
    LocalMux I__1500 (
            .O(N__7977),
            .I(BRIDGE_BASE_3));
    InMux I__1499 (
            .O(N__7972),
            .I(N__7964));
    InMux I__1498 (
            .O(N__7971),
            .I(N__7964));
    InMux I__1497 (
            .O(N__7970),
            .I(N__7959));
    InMux I__1496 (
            .O(N__7969),
            .I(N__7959));
    LocalMux I__1495 (
            .O(N__7964),
            .I(\U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2Z0Z_1 ));
    LocalMux I__1494 (
            .O(N__7959),
            .I(\U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2Z0Z_1 ));
    CascadeMux I__1493 (
            .O(N__7954),
            .I(N__7949));
    CascadeMux I__1492 (
            .O(N__7953),
            .I(N__7946));
    InMux I__1491 (
            .O(N__7952),
            .I(N__7943));
    InMux I__1490 (
            .O(N__7949),
            .I(N__7940));
    InMux I__1489 (
            .O(N__7946),
            .I(N__7937));
    LocalMux I__1488 (
            .O(N__7943),
            .I(N__7930));
    LocalMux I__1487 (
            .O(N__7940),
            .I(N__7930));
    LocalMux I__1486 (
            .O(N__7937),
            .I(N__7930));
    Span4Mux_v I__1485 (
            .O(N__7930),
            .I(N__7927));
    Sp12to4 I__1484 (
            .O(N__7927),
            .I(N__7924));
    Span12Mux_h I__1483 (
            .O(N__7924),
            .I(N__7921));
    Odrv12 I__1482 (
            .O(N__7921),
            .I(D_in_4));
    CascadeMux I__1481 (
            .O(N__7918),
            .I(N__7914));
    CascadeMux I__1480 (
            .O(N__7917),
            .I(N__7911));
    InMux I__1479 (
            .O(N__7914),
            .I(N__7891));
    InMux I__1478 (
            .O(N__7911),
            .I(N__7891));
    InMux I__1477 (
            .O(N__7910),
            .I(N__7891));
    InMux I__1476 (
            .O(N__7909),
            .I(N__7891));
    InMux I__1475 (
            .O(N__7908),
            .I(N__7891));
    InMux I__1474 (
            .O(N__7907),
            .I(N__7891));
    InMux I__1473 (
            .O(N__7906),
            .I(N__7881));
    InMux I__1472 (
            .O(N__7905),
            .I(N__7881));
    InMux I__1471 (
            .O(N__7904),
            .I(N__7881));
    LocalMux I__1470 (
            .O(N__7891),
            .I(N__7878));
    InMux I__1469 (
            .O(N__7890),
            .I(N__7866));
    InMux I__1468 (
            .O(N__7889),
            .I(N__7866));
    InMux I__1467 (
            .O(N__7888),
            .I(N__7866));
    LocalMux I__1466 (
            .O(N__7881),
            .I(N__7862));
    Span4Mux_v I__1465 (
            .O(N__7878),
            .I(N__7859));
    InMux I__1464 (
            .O(N__7877),
            .I(N__7854));
    InMux I__1463 (
            .O(N__7876),
            .I(N__7854));
    InMux I__1462 (
            .O(N__7875),
            .I(N__7847));
    InMux I__1461 (
            .O(N__7874),
            .I(N__7847));
    InMux I__1460 (
            .O(N__7873),
            .I(N__7847));
    LocalMux I__1459 (
            .O(N__7866),
            .I(N__7844));
    InMux I__1458 (
            .O(N__7865),
            .I(N__7841));
    Span4Mux_v I__1457 (
            .O(N__7862),
            .I(N__7832));
    Span4Mux_h I__1456 (
            .O(N__7859),
            .I(N__7832));
    LocalMux I__1455 (
            .O(N__7854),
            .I(N__7832));
    LocalMux I__1454 (
            .O(N__7847),
            .I(N__7832));
    Odrv4 I__1453 (
            .O(N__7844),
            .I(un1_AUTOCONFIG_SPACE));
    LocalMux I__1452 (
            .O(N__7841),
            .I(un1_AUTOCONFIG_SPACE));
    Odrv4 I__1451 (
            .O(N__7832),
            .I(un1_AUTOCONFIG_SPACE));
    CascadeMux I__1450 (
            .O(N__7825),
            .I(N_71_mux_cascade_));
    CascadeMux I__1449 (
            .O(N__7822),
            .I(N_23_cascade_));
    InMux I__1448 (
            .O(N__7819),
            .I(N__7816));
    LocalMux I__1447 (
            .O(N__7816),
            .I(\U409_ADDRESS_DECODE.m33Z0Z_3 ));
    InMux I__1446 (
            .O(N__7813),
            .I(N__7810));
    LocalMux I__1445 (
            .O(N__7810),
            .I(N__7806));
    InMux I__1444 (
            .O(N__7809),
            .I(N__7802));
    Span4Mux_v I__1443 (
            .O(N__7806),
            .I(N__7799));
    InMux I__1442 (
            .O(N__7805),
            .I(N__7794));
    LocalMux I__1441 (
            .O(N__7802),
            .I(N__7791));
    Sp12to4 I__1440 (
            .O(N__7799),
            .I(N__7788));
    InMux I__1439 (
            .O(N__7798),
            .I(N__7783));
    InMux I__1438 (
            .O(N__7797),
            .I(N__7783));
    LocalMux I__1437 (
            .O(N__7794),
            .I(N__7780));
    Span4Mux_v I__1436 (
            .O(N__7791),
            .I(N__7777));
    Span12Mux_h I__1435 (
            .O(N__7788),
            .I(N__7774));
    LocalMux I__1434 (
            .O(N__7783),
            .I(N__7771));
    Sp12to4 I__1433 (
            .O(N__7780),
            .I(N__7768));
    Span4Mux_v I__1432 (
            .O(N__7777),
            .I(N__7765));
    Span12Mux_v I__1431 (
            .O(N__7774),
            .I(N__7762));
    Span12Mux_v I__1430 (
            .O(N__7771),
            .I(N__7759));
    Span12Mux_v I__1429 (
            .O(N__7768),
            .I(N__7754));
    Sp12to4 I__1428 (
            .O(N__7765),
            .I(N__7754));
    Odrv12 I__1427 (
            .O(N__7762),
            .I(A_c_18));
    Odrv12 I__1426 (
            .O(N__7759),
            .I(A_c_18));
    Odrv12 I__1425 (
            .O(N__7754),
            .I(A_c_18));
    InMux I__1424 (
            .O(N__7747),
            .I(N__7743));
    InMux I__1423 (
            .O(N__7746),
            .I(N__7740));
    LocalMux I__1422 (
            .O(N__7743),
            .I(LIDE_BASE_1));
    LocalMux I__1421 (
            .O(N__7740),
            .I(LIDE_BASE_1));
    InMux I__1420 (
            .O(N__7735),
            .I(N__7729));
    InMux I__1419 (
            .O(N__7734),
            .I(N__7724));
    InMux I__1418 (
            .O(N__7733),
            .I(N__7724));
    CascadeMux I__1417 (
            .O(N__7732),
            .I(N__7720));
    LocalMux I__1416 (
            .O(N__7729),
            .I(N__7717));
    LocalMux I__1415 (
            .O(N__7724),
            .I(N__7714));
    InMux I__1414 (
            .O(N__7723),
            .I(N__7711));
    InMux I__1413 (
            .O(N__7720),
            .I(N__7707));
    Span4Mux_v I__1412 (
            .O(N__7717),
            .I(N__7704));
    Span4Mux_v I__1411 (
            .O(N__7714),
            .I(N__7701));
    LocalMux I__1410 (
            .O(N__7711),
            .I(N__7698));
    InMux I__1409 (
            .O(N__7710),
            .I(N__7695));
    LocalMux I__1408 (
            .O(N__7707),
            .I(N__7692));
    Span4Mux_v I__1407 (
            .O(N__7704),
            .I(N__7689));
    Sp12to4 I__1406 (
            .O(N__7701),
            .I(N__7686));
    Span4Mux_h I__1405 (
            .O(N__7698),
            .I(N__7681));
    LocalMux I__1404 (
            .O(N__7695),
            .I(N__7681));
    Span12Mux_v I__1403 (
            .O(N__7692),
            .I(N__7678));
    Span4Mux_v I__1402 (
            .O(N__7689),
            .I(N__7675));
    Span12Mux_h I__1401 (
            .O(N__7686),
            .I(N__7670));
    Sp12to4 I__1400 (
            .O(N__7681),
            .I(N__7670));
    Span12Mux_h I__1399 (
            .O(N__7678),
            .I(N__7667));
    Sp12to4 I__1398 (
            .O(N__7675),
            .I(N__7662));
    Span12Mux_v I__1397 (
            .O(N__7670),
            .I(N__7662));
    Odrv12 I__1396 (
            .O(N__7667),
            .I(A_c_17));
    Odrv12 I__1395 (
            .O(N__7662),
            .I(A_c_17));
    CascadeMux I__1394 (
            .O(N__7657),
            .I(N__7654));
    InMux I__1393 (
            .O(N__7654),
            .I(N__7650));
    InMux I__1392 (
            .O(N__7653),
            .I(N__7647));
    LocalMux I__1391 (
            .O(N__7650),
            .I(LIDE_BASE_2));
    LocalMux I__1390 (
            .O(N__7647),
            .I(LIDE_BASE_2));
    CascadeMux I__1389 (
            .O(N__7642),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_0_cascade_ ));
    CascadeMux I__1388 (
            .O(N__7639),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_ ));
    CascadeMux I__1387 (
            .O(N__7636),
            .I(N__7632));
    InMux I__1386 (
            .O(N__7635),
            .I(N__7626));
    InMux I__1385 (
            .O(N__7632),
            .I(N__7626));
    InMux I__1384 (
            .O(N__7631),
            .I(N__7621));
    LocalMux I__1383 (
            .O(N__7626),
            .I(N__7617));
    InMux I__1382 (
            .O(N__7625),
            .I(N__7614));
    InMux I__1381 (
            .O(N__7624),
            .I(N__7609));
    LocalMux I__1380 (
            .O(N__7621),
            .I(N__7605));
    InMux I__1379 (
            .O(N__7620),
            .I(N__7602));
    Span4Mux_h I__1378 (
            .O(N__7617),
            .I(N__7597));
    LocalMux I__1377 (
            .O(N__7614),
            .I(N__7597));
    InMux I__1376 (
            .O(N__7613),
            .I(N__7594));
    InMux I__1375 (
            .O(N__7612),
            .I(N__7591));
    LocalMux I__1374 (
            .O(N__7609),
            .I(N__7588));
    InMux I__1373 (
            .O(N__7608),
            .I(N__7585));
    Odrv12 I__1372 (
            .O(N__7605),
            .I(CONFIGURED));
    LocalMux I__1371 (
            .O(N__7602),
            .I(CONFIGURED));
    Odrv4 I__1370 (
            .O(N__7597),
            .I(CONFIGURED));
    LocalMux I__1369 (
            .O(N__7594),
            .I(CONFIGURED));
    LocalMux I__1368 (
            .O(N__7591),
            .I(CONFIGURED));
    Odrv4 I__1367 (
            .O(N__7588),
            .I(CONFIGURED));
    LocalMux I__1366 (
            .O(N__7585),
            .I(CONFIGURED));
    InMux I__1365 (
            .O(N__7570),
            .I(N__7567));
    LocalMux I__1364 (
            .O(N__7567),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3 ));
    CascadeMux I__1363 (
            .O(N__7564),
            .I(N__7561));
    InMux I__1362 (
            .O(N__7561),
            .I(N__7557));
    InMux I__1361 (
            .O(N__7560),
            .I(N__7554));
    LocalMux I__1360 (
            .O(N__7557),
            .I(LIDE_BASE_6));
    LocalMux I__1359 (
            .O(N__7554),
            .I(LIDE_BASE_6));
    InMux I__1358 (
            .O(N__7549),
            .I(N__7545));
    InMux I__1357 (
            .O(N__7548),
            .I(N__7542));
    LocalMux I__1356 (
            .O(N__7545),
            .I(LIDE_BASE_5));
    LocalMux I__1355 (
            .O(N__7542),
            .I(LIDE_BASE_5));
    InMux I__1354 (
            .O(N__7537),
            .I(N__7534));
    LocalMux I__1353 (
            .O(N__7534),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2 ));
    InMux I__1352 (
            .O(N__7531),
            .I(N__7526));
    InMux I__1351 (
            .O(N__7530),
            .I(N__7521));
    InMux I__1350 (
            .O(N__7529),
            .I(N__7521));
    LocalMux I__1349 (
            .O(N__7526),
            .I(\U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1Z0Z_0 ));
    LocalMux I__1348 (
            .O(N__7521),
            .I(\U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1Z0Z_0 ));
    InMux I__1347 (
            .O(N__7516),
            .I(N__7513));
    LocalMux I__1346 (
            .O(N__7513),
            .I(N__7509));
    CascadeMux I__1345 (
            .O(N__7512),
            .I(N__7506));
    Span4Mux_v I__1344 (
            .O(N__7509),
            .I(N__7503));
    InMux I__1343 (
            .O(N__7506),
            .I(N__7500));
    Odrv4 I__1342 (
            .O(N__7503),
            .I(BRIDGE_BASE_5));
    LocalMux I__1341 (
            .O(N__7500),
            .I(BRIDGE_BASE_5));
    InMux I__1340 (
            .O(N__7495),
            .I(N__7490));
    InMux I__1339 (
            .O(N__7494),
            .I(N__7485));
    InMux I__1338 (
            .O(N__7493),
            .I(N__7485));
    LocalMux I__1337 (
            .O(N__7490),
            .I(N__7482));
    LocalMux I__1336 (
            .O(N__7485),
            .I(\U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2Z0Z_0 ));
    Odrv4 I__1335 (
            .O(N__7482),
            .I(\U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2Z0Z_0 ));
    InMux I__1334 (
            .O(N__7477),
            .I(N__7474));
    LocalMux I__1333 (
            .O(N__7474),
            .I(N__7471));
    Span4Mux_v I__1332 (
            .O(N__7471),
            .I(N__7468));
    Span4Mux_h I__1331 (
            .O(N__7468),
            .I(N__7464));
    InMux I__1330 (
            .O(N__7467),
            .I(N__7461));
    Odrv4 I__1329 (
            .O(N__7464),
            .I(\U409_AUTOCONFIG.un1_AZ0Z_13 ));
    LocalMux I__1328 (
            .O(N__7461),
            .I(\U409_AUTOCONFIG.un1_AZ0Z_13 ));
    InMux I__1327 (
            .O(N__7456),
            .I(N__7452));
    InMux I__1326 (
            .O(N__7455),
            .I(N__7445));
    LocalMux I__1325 (
            .O(N__7452),
            .I(N__7442));
    InMux I__1324 (
            .O(N__7451),
            .I(N__7439));
    CascadeMux I__1323 (
            .O(N__7450),
            .I(N__7432));
    InMux I__1322 (
            .O(N__7449),
            .I(N__7429));
    InMux I__1321 (
            .O(N__7448),
            .I(N__7424));
    LocalMux I__1320 (
            .O(N__7445),
            .I(N__7417));
    Span4Mux_v I__1319 (
            .O(N__7442),
            .I(N__7417));
    LocalMux I__1318 (
            .O(N__7439),
            .I(N__7417));
    InMux I__1317 (
            .O(N__7438),
            .I(N__7408));
    InMux I__1316 (
            .O(N__7437),
            .I(N__7408));
    InMux I__1315 (
            .O(N__7436),
            .I(N__7408));
    InMux I__1314 (
            .O(N__7435),
            .I(N__7408));
    InMux I__1313 (
            .O(N__7432),
            .I(N__7403));
    LocalMux I__1312 (
            .O(N__7429),
            .I(N__7400));
    InMux I__1311 (
            .O(N__7428),
            .I(N__7397));
    InMux I__1310 (
            .O(N__7427),
            .I(N__7394));
    LocalMux I__1309 (
            .O(N__7424),
            .I(N__7387));
    Span4Mux_v I__1308 (
            .O(N__7417),
            .I(N__7387));
    LocalMux I__1307 (
            .O(N__7408),
            .I(N__7387));
    InMux I__1306 (
            .O(N__7407),
            .I(N__7384));
    InMux I__1305 (
            .O(N__7406),
            .I(N__7381));
    LocalMux I__1304 (
            .O(N__7403),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    Odrv12 I__1303 (
            .O(N__7400),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    LocalMux I__1302 (
            .O(N__7397),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    LocalMux I__1301 (
            .O(N__7394),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    Odrv4 I__1300 (
            .O(N__7387),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    LocalMux I__1299 (
            .O(N__7384),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    LocalMux I__1298 (
            .O(N__7381),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    InMux I__1297 (
            .O(N__7366),
            .I(N__7363));
    LocalMux I__1296 (
            .O(N__7363),
            .I(\U409_CIA.un1_CIA_CLK_COUNT_3_2 ));
    InMux I__1295 (
            .O(N__7360),
            .I(N__7354));
    InMux I__1294 (
            .O(N__7359),
            .I(N__7351));
    InMux I__1293 (
            .O(N__7358),
            .I(N__7346));
    InMux I__1292 (
            .O(N__7357),
            .I(N__7346));
    LocalMux I__1291 (
            .O(N__7354),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1290 (
            .O(N__7351),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1289 (
            .O(N__7346),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    CascadeMux I__1288 (
            .O(N__7339),
            .I(N__7333));
    InMux I__1287 (
            .O(N__7338),
            .I(N__7330));
    InMux I__1286 (
            .O(N__7337),
            .I(N__7327));
    InMux I__1285 (
            .O(N__7336),
            .I(N__7324));
    InMux I__1284 (
            .O(N__7333),
            .I(N__7321));
    LocalMux I__1283 (
            .O(N__7330),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1282 (
            .O(N__7327),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1281 (
            .O(N__7324),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1280 (
            .O(N__7321),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    CascadeMux I__1279 (
            .O(N__7312),
            .I(N__7308));
    InMux I__1278 (
            .O(N__7311),
            .I(N__7303));
    InMux I__1277 (
            .O(N__7308),
            .I(N__7300));
    InMux I__1276 (
            .O(N__7307),
            .I(N__7297));
    InMux I__1275 (
            .O(N__7306),
            .I(N__7294));
    LocalMux I__1274 (
            .O(N__7303),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__1273 (
            .O(N__7300),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__1272 (
            .O(N__7297),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__1271 (
            .O(N__7294),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    InMux I__1270 (
            .O(N__7285),
            .I(N__7279));
    InMux I__1269 (
            .O(N__7284),
            .I(N__7276));
    InMux I__1268 (
            .O(N__7283),
            .I(N__7271));
    InMux I__1267 (
            .O(N__7282),
            .I(N__7271));
    LocalMux I__1266 (
            .O(N__7279),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1265 (
            .O(N__7276),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1264 (
            .O(N__7271),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    CascadeMux I__1263 (
            .O(N__7264),
            .I(\U409_CIA.CIA_CLK_COUNT11_3_cascade_ ));
    InMux I__1262 (
            .O(N__7261),
            .I(N__7255));
    InMux I__1261 (
            .O(N__7260),
            .I(N__7255));
    LocalMux I__1260 (
            .O(N__7255),
            .I(\U409_CIA.CIA_CLK_COUNT11 ));
    InMux I__1259 (
            .O(N__7252),
            .I(N__7242));
    InMux I__1258 (
            .O(N__7251),
            .I(N__7242));
    InMux I__1257 (
            .O(N__7250),
            .I(N__7233));
    InMux I__1256 (
            .O(N__7249),
            .I(N__7233));
    InMux I__1255 (
            .O(N__7248),
            .I(N__7233));
    InMux I__1254 (
            .O(N__7247),
            .I(N__7233));
    LocalMux I__1253 (
            .O(N__7242),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1252 (
            .O(N__7233),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    CascadeMux I__1251 (
            .O(N__7228),
            .I(N__7221));
    CascadeMux I__1250 (
            .O(N__7227),
            .I(N__7218));
    CascadeMux I__1249 (
            .O(N__7226),
            .I(N__7215));
    InMux I__1248 (
            .O(N__7225),
            .I(N__7211));
    InMux I__1247 (
            .O(N__7224),
            .I(N__7206));
    InMux I__1246 (
            .O(N__7221),
            .I(N__7206));
    InMux I__1245 (
            .O(N__7218),
            .I(N__7199));
    InMux I__1244 (
            .O(N__7215),
            .I(N__7199));
    InMux I__1243 (
            .O(N__7214),
            .I(N__7199));
    LocalMux I__1242 (
            .O(N__7211),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1241 (
            .O(N__7206),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1240 (
            .O(N__7199),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    CascadeMux I__1239 (
            .O(N__7192),
            .I(N__7188));
    InMux I__1238 (
            .O(N__7191),
            .I(N__7182));
    InMux I__1237 (
            .O(N__7188),
            .I(N__7182));
    InMux I__1236 (
            .O(N__7187),
            .I(N__7179));
    LocalMux I__1235 (
            .O(N__7182),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    LocalMux I__1234 (
            .O(N__7179),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    InMux I__1233 (
            .O(N__7174),
            .I(N__7167));
    InMux I__1232 (
            .O(N__7173),
            .I(N__7167));
    InMux I__1231 (
            .O(N__7172),
            .I(N__7164));
    LocalMux I__1230 (
            .O(N__7167),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__1229 (
            .O(N__7164),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    InMux I__1228 (
            .O(N__7159),
            .I(N__7155));
    InMux I__1227 (
            .O(N__7158),
            .I(N__7152));
    LocalMux I__1226 (
            .O(N__7155),
            .I(\U409_CIA.CLK_CIA6_4 ));
    LocalMux I__1225 (
            .O(N__7152),
            .I(\U409_CIA.CLK_CIA6_4 ));
    CascadeMux I__1224 (
            .O(N__7147),
            .I(\U409_ADDRESS_DECODE.N_77_mux_cascade_ ));
    IoInMux I__1223 (
            .O(N__7144),
            .I(N__7141));
    LocalMux I__1222 (
            .O(N__7141),
            .I(N__7138));
    IoSpan4Mux I__1221 (
            .O(N__7138),
            .I(N__7135));
    Span4Mux_s3_h I__1220 (
            .O(N__7135),
            .I(N__7132));
    Sp12to4 I__1219 (
            .O(N__7132),
            .I(N__7129));
    Span12Mux_s8_h I__1218 (
            .O(N__7129),
            .I(N__7126));
    Odrv12 I__1217 (
            .O(N__7126),
            .I(N_22_0_i));
    InMux I__1216 (
            .O(N__7123),
            .I(N__7120));
    LocalMux I__1215 (
            .O(N__7120),
            .I(N__7117));
    Span4Mux_h I__1214 (
            .O(N__7117),
            .I(N__7113));
    InMux I__1213 (
            .O(N__7116),
            .I(N__7110));
    Span4Mux_v I__1212 (
            .O(N__7113),
            .I(N__7107));
    LocalMux I__1211 (
            .O(N__7110),
            .I(N__7104));
    Odrv4 I__1210 (
            .O(N__7107),
            .I(U409_ADDRESS_DECODE_un1_RTC_ENn));
    Odrv4 I__1209 (
            .O(N__7104),
            .I(U409_ADDRESS_DECODE_un1_RTC_ENn));
    InMux I__1208 (
            .O(N__7099),
            .I(N__7096));
    LocalMux I__1207 (
            .O(N__7096),
            .I(N__7093));
    Span4Mux_h I__1206 (
            .O(N__7093),
            .I(N__7090));
    Span4Mux_v I__1205 (
            .O(N__7090),
            .I(N__7087));
    Odrv4 I__1204 (
            .O(N__7087),
            .I(\U409_ADDRESS_DECODE.PORTSIZE_2 ));
    InMux I__1203 (
            .O(N__7084),
            .I(N__7078));
    InMux I__1202 (
            .O(N__7083),
            .I(N__7078));
    LocalMux I__1201 (
            .O(N__7078),
            .I(BRIDGE_BASE_7));
    InMux I__1200 (
            .O(N__7075),
            .I(N__7070));
    InMux I__1199 (
            .O(N__7074),
            .I(N__7066));
    InMux I__1198 (
            .O(N__7073),
            .I(N__7063));
    LocalMux I__1197 (
            .O(N__7070),
            .I(N__7060));
    InMux I__1196 (
            .O(N__7069),
            .I(N__7057));
    LocalMux I__1195 (
            .O(N__7066),
            .I(N__7052));
    LocalMux I__1194 (
            .O(N__7063),
            .I(N__7052));
    Span4Mux_v I__1193 (
            .O(N__7060),
            .I(N__7049));
    LocalMux I__1192 (
            .O(N__7057),
            .I(N__7046));
    Span4Mux_v I__1191 (
            .O(N__7052),
            .I(N__7041));
    Span4Mux_h I__1190 (
            .O(N__7049),
            .I(N__7036));
    Span4Mux_v I__1189 (
            .O(N__7046),
            .I(N__7036));
    InMux I__1188 (
            .O(N__7045),
            .I(N__7033));
    InMux I__1187 (
            .O(N__7044),
            .I(N__7030));
    Sp12to4 I__1186 (
            .O(N__7041),
            .I(N__7021));
    Sp12to4 I__1185 (
            .O(N__7036),
            .I(N__7021));
    LocalMux I__1184 (
            .O(N__7033),
            .I(N__7021));
    LocalMux I__1183 (
            .O(N__7030),
            .I(N__7021));
    Odrv12 I__1182 (
            .O(N__7021),
            .I(A_c_7));
    InMux I__1181 (
            .O(N__7018),
            .I(N__7013));
    InMux I__1180 (
            .O(N__7017),
            .I(N__7010));
    InMux I__1179 (
            .O(N__7016),
            .I(N__7007));
    LocalMux I__1178 (
            .O(N__7013),
            .I(N__7004));
    LocalMux I__1177 (
            .O(N__7010),
            .I(N__6998));
    LocalMux I__1176 (
            .O(N__7007),
            .I(N__6998));
    Span4Mux_v I__1175 (
            .O(N__7004),
            .I(N__6994));
    InMux I__1174 (
            .O(N__7003),
            .I(N__6991));
    Span4Mux_v I__1173 (
            .O(N__6998),
            .I(N__6988));
    InMux I__1172 (
            .O(N__6997),
            .I(N__6985));
    Sp12to4 I__1171 (
            .O(N__6994),
            .I(N__6976));
    LocalMux I__1170 (
            .O(N__6991),
            .I(N__6976));
    Sp12to4 I__1169 (
            .O(N__6988),
            .I(N__6976));
    LocalMux I__1168 (
            .O(N__6985),
            .I(N__6976));
    Span12Mux_h I__1167 (
            .O(N__6976),
            .I(N__6973));
    Odrv12 I__1166 (
            .O(N__6973),
            .I(A_c_5));
    CascadeMux I__1165 (
            .O(N__6970),
            .I(N__6967));
    InMux I__1164 (
            .O(N__6967),
            .I(N__6964));
    LocalMux I__1163 (
            .O(N__6964),
            .I(N__6961));
    Span4Mux_h I__1162 (
            .O(N__6961),
            .I(N__6958));
    Odrv4 I__1161 (
            .O(N__6958),
            .I(\U409_AUTOCONFIG.un1_STATE_6Z0Z_1 ));
    InMux I__1160 (
            .O(N__6955),
            .I(N__6950));
    InMux I__1159 (
            .O(N__6954),
            .I(N__6945));
    InMux I__1158 (
            .O(N__6953),
            .I(N__6945));
    LocalMux I__1157 (
            .O(N__6950),
            .I(\U409_AUTOCONFIG.un1_STATE_6_0 ));
    LocalMux I__1156 (
            .O(N__6945),
            .I(\U409_AUTOCONFIG.un1_STATE_6_0 ));
    CascadeMux I__1155 (
            .O(N__6940),
            .I(N__6935));
    CascadeMux I__1154 (
            .O(N__6939),
            .I(N__6929));
    CascadeMux I__1153 (
            .O(N__6938),
            .I(N__6924));
    InMux I__1152 (
            .O(N__6935),
            .I(N__6916));
    InMux I__1151 (
            .O(N__6934),
            .I(N__6916));
    CascadeMux I__1150 (
            .O(N__6933),
            .I(N__6913));
    InMux I__1149 (
            .O(N__6932),
            .I(N__6904));
    InMux I__1148 (
            .O(N__6929),
            .I(N__6904));
    InMux I__1147 (
            .O(N__6928),
            .I(N__6904));
    InMux I__1146 (
            .O(N__6927),
            .I(N__6901));
    InMux I__1145 (
            .O(N__6924),
            .I(N__6895));
    InMux I__1144 (
            .O(N__6923),
            .I(N__6895));
    CascadeMux I__1143 (
            .O(N__6922),
            .I(N__6891));
    CascadeMux I__1142 (
            .O(N__6921),
            .I(N__6888));
    LocalMux I__1141 (
            .O(N__6916),
            .I(N__6882));
    InMux I__1140 (
            .O(N__6913),
            .I(N__6879));
    InMux I__1139 (
            .O(N__6912),
            .I(N__6876));
    InMux I__1138 (
            .O(N__6911),
            .I(N__6873));
    LocalMux I__1137 (
            .O(N__6904),
            .I(N__6868));
    LocalMux I__1136 (
            .O(N__6901),
            .I(N__6868));
    InMux I__1135 (
            .O(N__6900),
            .I(N__6865));
    LocalMux I__1134 (
            .O(N__6895),
            .I(N__6861));
    InMux I__1133 (
            .O(N__6894),
            .I(N__6854));
    InMux I__1132 (
            .O(N__6891),
            .I(N__6854));
    InMux I__1131 (
            .O(N__6888),
            .I(N__6854));
    CascadeMux I__1130 (
            .O(N__6887),
            .I(N__6851));
    CascadeMux I__1129 (
            .O(N__6886),
            .I(N__6846));
    CascadeMux I__1128 (
            .O(N__6885),
            .I(N__6843));
    Span4Mux_v I__1127 (
            .O(N__6882),
            .I(N__6838));
    LocalMux I__1126 (
            .O(N__6879),
            .I(N__6838));
    LocalMux I__1125 (
            .O(N__6876),
            .I(N__6835));
    LocalMux I__1124 (
            .O(N__6873),
            .I(N__6832));
    Span4Mux_v I__1123 (
            .O(N__6868),
            .I(N__6829));
    LocalMux I__1122 (
            .O(N__6865),
            .I(N__6826));
    InMux I__1121 (
            .O(N__6864),
            .I(N__6823));
    Span4Mux_v I__1120 (
            .O(N__6861),
            .I(N__6818));
    LocalMux I__1119 (
            .O(N__6854),
            .I(N__6818));
    InMux I__1118 (
            .O(N__6851),
            .I(N__6813));
    InMux I__1117 (
            .O(N__6850),
            .I(N__6813));
    InMux I__1116 (
            .O(N__6849),
            .I(N__6806));
    InMux I__1115 (
            .O(N__6846),
            .I(N__6806));
    InMux I__1114 (
            .O(N__6843),
            .I(N__6806));
    Span4Mux_v I__1113 (
            .O(N__6838),
            .I(N__6803));
    Span4Mux_v I__1112 (
            .O(N__6835),
            .I(N__6798));
    Span4Mux_v I__1111 (
            .O(N__6832),
            .I(N__6798));
    Span4Mux_h I__1110 (
            .O(N__6829),
            .I(N__6793));
    Span4Mux_v I__1109 (
            .O(N__6826),
            .I(N__6793));
    LocalMux I__1108 (
            .O(N__6823),
            .I(N__6784));
    Sp12to4 I__1107 (
            .O(N__6818),
            .I(N__6784));
    LocalMux I__1106 (
            .O(N__6813),
            .I(N__6784));
    LocalMux I__1105 (
            .O(N__6806),
            .I(N__6784));
    Sp12to4 I__1104 (
            .O(N__6803),
            .I(N__6779));
    Sp12to4 I__1103 (
            .O(N__6798),
            .I(N__6779));
    Span4Mux_h I__1102 (
            .O(N__6793),
            .I(N__6776));
    Span12Mux_h I__1101 (
            .O(N__6784),
            .I(N__6773));
    Span12Mux_h I__1100 (
            .O(N__6779),
            .I(N__6768));
    Sp12to4 I__1099 (
            .O(N__6776),
            .I(N__6768));
    Span12Mux_v I__1098 (
            .O(N__6773),
            .I(N__6765));
    Span12Mux_v I__1097 (
            .O(N__6768),
            .I(N__6762));
    Odrv12 I__1096 (
            .O(N__6765),
            .I(A_c_1));
    Odrv12 I__1095 (
            .O(N__6762),
            .I(A_c_1));
    CascadeMux I__1094 (
            .O(N__6757),
            .I(\U409_AUTOCONFIG.un1_STATE_6_0_cascade_ ));
    CascadeMux I__1093 (
            .O(N__6754),
            .I(N__6749));
    InMux I__1092 (
            .O(N__6753),
            .I(N__6746));
    CascadeMux I__1091 (
            .O(N__6752),
            .I(N__6741));
    InMux I__1090 (
            .O(N__6749),
            .I(N__6738));
    LocalMux I__1089 (
            .O(N__6746),
            .I(N__6735));
    InMux I__1088 (
            .O(N__6745),
            .I(N__6728));
    InMux I__1087 (
            .O(N__6744),
            .I(N__6728));
    InMux I__1086 (
            .O(N__6741),
            .I(N__6728));
    LocalMux I__1085 (
            .O(N__6738),
            .I(N__6725));
    Span4Mux_h I__1084 (
            .O(N__6735),
            .I(N__6722));
    LocalMux I__1083 (
            .O(N__6728),
            .I(N__6719));
    Span4Mux_v I__1082 (
            .O(N__6725),
            .I(N__6716));
    Span4Mux_v I__1081 (
            .O(N__6722),
            .I(N__6713));
    Span4Mux_h I__1080 (
            .O(N__6719),
            .I(N__6710));
    Sp12to4 I__1079 (
            .O(N__6716),
            .I(N__6707));
    Sp12to4 I__1078 (
            .O(N__6713),
            .I(N__6702));
    Sp12to4 I__1077 (
            .O(N__6710),
            .I(N__6702));
    Span12Mux_h I__1076 (
            .O(N__6707),
            .I(N__6699));
    Span12Mux_v I__1075 (
            .O(N__6702),
            .I(N__6696));
    Odrv12 I__1074 (
            .O(N__6699),
            .I(D_in_6));
    Odrv12 I__1073 (
            .O(N__6696),
            .I(D_in_6));
    CascadeMux I__1072 (
            .O(N__6691),
            .I(\U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1Z0Z_0_cascade_ ));
    CascadeMux I__1071 (
            .O(N__6688),
            .I(N__6685));
    InMux I__1070 (
            .O(N__6685),
            .I(N__6679));
    InMux I__1069 (
            .O(N__6684),
            .I(N__6679));
    LocalMux I__1068 (
            .O(N__6679),
            .I(BRIDGE_BASE_6));
    InMux I__1067 (
            .O(N__6676),
            .I(N__6673));
    LocalMux I__1066 (
            .O(N__6673),
            .I(N__6669));
    InMux I__1065 (
            .O(N__6672),
            .I(N__6666));
    Span4Mux_h I__1064 (
            .O(N__6669),
            .I(N__6661));
    LocalMux I__1063 (
            .O(N__6666),
            .I(N__6661));
    Odrv4 I__1062 (
            .O(N__6661),
            .I(CIA_SPACE));
    CascadeMux I__1061 (
            .O(N__6658),
            .I(\U409_CIA.VMA_RNOZ0Z_0_cascade_ ));
    CascadeMux I__1060 (
            .O(N__6655),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENn_2_cascade_ ));
    IoInMux I__1059 (
            .O(N__6652),
            .I(N__6649));
    LocalMux I__1058 (
            .O(N__6649),
            .I(N__6646));
    IoSpan4Mux I__1057 (
            .O(N__6646),
            .I(N__6643));
    Span4Mux_s2_v I__1056 (
            .O(N__6643),
            .I(N__6640));
    Span4Mux_h I__1055 (
            .O(N__6640),
            .I(N__6637));
    Sp12to4 I__1054 (
            .O(N__6637),
            .I(N__6634));
    Span12Mux_v I__1053 (
            .O(N__6634),
            .I(N__6631));
    Odrv12 I__1052 (
            .O(N__6631),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn_i));
    InMux I__1051 (
            .O(N__6628),
            .I(N__6625));
    LocalMux I__1050 (
            .O(N__6625),
            .I(N__6621));
    InMux I__1049 (
            .O(N__6624),
            .I(N__6618));
    Span4Mux_h I__1048 (
            .O(N__6621),
            .I(N__6614));
    LocalMux I__1047 (
            .O(N__6618),
            .I(N__6611));
    InMux I__1046 (
            .O(N__6617),
            .I(N__6608));
    Odrv4 I__1045 (
            .O(N__6614),
            .I(\U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1 ));
    Odrv4 I__1044 (
            .O(N__6611),
            .I(\U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1 ));
    LocalMux I__1043 (
            .O(N__6608),
            .I(\U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1 ));
    InMux I__1042 (
            .O(N__6601),
            .I(N__6595));
    InMux I__1041 (
            .O(N__6600),
            .I(N__6595));
    LocalMux I__1040 (
            .O(N__6595),
            .I(BRIDGE_BASE_0));
    InMux I__1039 (
            .O(N__6592),
            .I(N__6589));
    LocalMux I__1038 (
            .O(N__6589),
            .I(N__6586));
    Odrv4 I__1037 (
            .O(N__6586),
            .I(\U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_4 ));
    InMux I__1036 (
            .O(N__6583),
            .I(N__6580));
    LocalMux I__1035 (
            .O(N__6580),
            .I(N__6577));
    Odrv4 I__1034 (
            .O(N__6577),
            .I(\U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_3 ));
    CascadeMux I__1033 (
            .O(N__6574),
            .I(\U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_1_cascade_ ));
    InMux I__1032 (
            .O(N__6571),
            .I(N__6568));
    LocalMux I__1031 (
            .O(N__6568),
            .I(\U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_2 ));
    IoInMux I__1030 (
            .O(N__6565),
            .I(N__6562));
    LocalMux I__1029 (
            .O(N__6562),
            .I(N__6559));
    IoSpan4Mux I__1028 (
            .O(N__6559),
            .I(N__6556));
    Sp12to4 I__1027 (
            .O(N__6556),
            .I(N__6553));
    Span12Mux_s7_h I__1026 (
            .O(N__6553),
            .I(N__6550));
    Span12Mux_h I__1025 (
            .O(N__6550),
            .I(N__6547));
    Odrv12 I__1024 (
            .O(N__6547),
            .I(U409_ADDRESS_DECODE_un1_BREG_ENn_i));
    InMux I__1023 (
            .O(N__6544),
            .I(N__6540));
    InMux I__1022 (
            .O(N__6543),
            .I(N__6536));
    LocalMux I__1021 (
            .O(N__6540),
            .I(N__6530));
    InMux I__1020 (
            .O(N__6539),
            .I(N__6527));
    LocalMux I__1019 (
            .O(N__6536),
            .I(N__6524));
    InMux I__1018 (
            .O(N__6535),
            .I(N__6519));
    InMux I__1017 (
            .O(N__6534),
            .I(N__6519));
    InMux I__1016 (
            .O(N__6533),
            .I(N__6515));
    Span4Mux_v I__1015 (
            .O(N__6530),
            .I(N__6506));
    LocalMux I__1014 (
            .O(N__6527),
            .I(N__6506));
    Span4Mux_h I__1013 (
            .O(N__6524),
            .I(N__6506));
    LocalMux I__1012 (
            .O(N__6519),
            .I(N__6506));
    InMux I__1011 (
            .O(N__6518),
            .I(N__6503));
    LocalMux I__1010 (
            .O(N__6515),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    Odrv4 I__1009 (
            .O(N__6506),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    LocalMux I__1008 (
            .O(N__6503),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    InMux I__1007 (
            .O(N__6496),
            .I(N__6493));
    LocalMux I__1006 (
            .O(N__6493),
            .I(N__6490));
    Odrv4 I__1005 (
            .O(N__6490),
            .I(\U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_0 ));
    InMux I__1004 (
            .O(N__6487),
            .I(N__6484));
    LocalMux I__1003 (
            .O(N__6484),
            .I(N__6480));
    InMux I__1002 (
            .O(N__6483),
            .I(N__6477));
    Odrv4 I__1001 (
            .O(N__6480),
            .I(BRIDGE_BASE_4));
    LocalMux I__1000 (
            .O(N__6477),
            .I(BRIDGE_BASE_4));
    InMux I__999 (
            .O(N__6472),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ));
    InMux I__998 (
            .O(N__6469),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ));
    InMux I__997 (
            .O(N__6466),
            .I(N__6463));
    LocalMux I__996 (
            .O(N__6463),
            .I(\U409_CIA.CLK_CIA6_3 ));
    InMux I__995 (
            .O(N__6460),
            .I(N__6457));
    LocalMux I__994 (
            .O(N__6457),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0 ));
    IoInMux I__993 (
            .O(N__6454),
            .I(N__6451));
    LocalMux I__992 (
            .O(N__6451),
            .I(N__6448));
    IoSpan4Mux I__991 (
            .O(N__6448),
            .I(N__6445));
    Sp12to4 I__990 (
            .O(N__6445),
            .I(N__6442));
    Span12Mux_s7_h I__989 (
            .O(N__6442),
            .I(N__6439));
    Span12Mux_h I__988 (
            .O(N__6439),
            .I(N__6436));
    Odrv12 I__987 (
            .O(N__6436),
            .I(U409_ADDRESS_DECODE_un1_RTC_ENn_i));
    CascadeMux I__986 (
            .O(N__6433),
            .I(N__6430));
    InMux I__985 (
            .O(N__6430),
            .I(N__6426));
    InMux I__984 (
            .O(N__6429),
            .I(N__6423));
    LocalMux I__983 (
            .O(N__6426),
            .I(BRIDGE_BASE_2));
    LocalMux I__982 (
            .O(N__6423),
            .I(BRIDGE_BASE_2));
    InMux I__981 (
            .O(N__6418),
            .I(N__6415));
    LocalMux I__980 (
            .O(N__6415),
            .I(\U409_AUTOCONFIG.AC_STARTZ0 ));
    InMux I__979 (
            .O(N__6412),
            .I(N__6409));
    LocalMux I__978 (
            .O(N__6409),
            .I(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_a3_0 ));
    CascadeMux I__977 (
            .O(N__6406),
            .I(\U409_CIA.CLK_CIA_r_1_0_cascade_ ));
    InMux I__976 (
            .O(N__6403),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ));
    InMux I__975 (
            .O(N__6400),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ));
    InMux I__974 (
            .O(N__6397),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ));
    InMux I__973 (
            .O(N__6394),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ));
    InMux I__972 (
            .O(N__6391),
            .I(N__6388));
    LocalMux I__971 (
            .O(N__6388),
            .I(\U409_AUTOCONFIG.PR_OUTZ0Z_0 ));
    CascadeMux I__970 (
            .O(N__6385),
            .I(\U409_AUTOCONFIG.LIDE_OUT_RNI5BMPZ0Z_0_cascade_ ));
    InMux I__969 (
            .O(N__6382),
            .I(N__6375));
    InMux I__968 (
            .O(N__6381),
            .I(N__6375));
    InMux I__967 (
            .O(N__6380),
            .I(N__6372));
    LocalMux I__966 (
            .O(N__6375),
            .I(\U409_AUTOCONFIG.D_OUT_sm0_0 ));
    LocalMux I__965 (
            .O(N__6372),
            .I(\U409_AUTOCONFIG.D_OUT_sm0_0 ));
    IoInMux I__964 (
            .O(N__6367),
            .I(N__6364));
    LocalMux I__963 (
            .O(N__6364),
            .I(N__6361));
    IoSpan4Mux I__962 (
            .O(N__6361),
            .I(N__6358));
    Sp12to4 I__961 (
            .O(N__6358),
            .I(N__6355));
    Span12Mux_s7_v I__960 (
            .O(N__6355),
            .I(N__6352));
    Odrv12 I__959 (
            .O(N__6352),
            .I(D_OUT_0));
    InMux I__958 (
            .O(N__6349),
            .I(N__6345));
    InMux I__957 (
            .O(N__6348),
            .I(N__6342));
    LocalMux I__956 (
            .O(N__6345),
            .I(\U409_AUTOCONFIG.N_90 ));
    LocalMux I__955 (
            .O(N__6342),
            .I(\U409_AUTOCONFIG.N_90 ));
    InMux I__954 (
            .O(N__6337),
            .I(N__6334));
    LocalMux I__953 (
            .O(N__6334),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ));
    InMux I__952 (
            .O(N__6331),
            .I(N__6328));
    LocalMux I__951 (
            .O(N__6328),
            .I(\U409_AUTOCONFIG.N_98 ));
    InMux I__950 (
            .O(N__6325),
            .I(N__6322));
    LocalMux I__949 (
            .O(N__6322),
            .I(N__6319));
    Span12Mux_h I__948 (
            .O(N__6319),
            .I(N__6316));
    Span12Mux_v I__947 (
            .O(N__6316),
            .I(N__6313));
    Odrv12 I__946 (
            .O(N__6313),
            .I(CPUCONFn_c));
    CascadeMux I__945 (
            .O(N__6310),
            .I(\U409_AUTOCONFIG.STATE4_cascade_ ));
    InMux I__944 (
            .O(N__6307),
            .I(N__6303));
    InMux I__943 (
            .O(N__6306),
            .I(N__6300));
    LocalMux I__942 (
            .O(N__6303),
            .I(N__6295));
    LocalMux I__941 (
            .O(N__6300),
            .I(N__6295));
    Span4Mux_v I__940 (
            .O(N__6295),
            .I(N__6292));
    Odrv4 I__939 (
            .O(N__6292),
            .I(\U409_AUTOCONFIG.N_104 ));
    CascadeMux I__938 (
            .O(N__6289),
            .I(\U409_AUTOCONFIG.N_103_cascade_ ));
    InMux I__937 (
            .O(N__6286),
            .I(N__6283));
    LocalMux I__936 (
            .O(N__6283),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ));
    CEMux I__935 (
            .O(N__6280),
            .I(N__6275));
    CEMux I__934 (
            .O(N__6279),
            .I(N__6272));
    CEMux I__933 (
            .O(N__6278),
            .I(N__6269));
    LocalMux I__932 (
            .O(N__6275),
            .I(N__6264));
    LocalMux I__931 (
            .O(N__6272),
            .I(N__6261));
    LocalMux I__930 (
            .O(N__6269),
            .I(N__6258));
    CEMux I__929 (
            .O(N__6268),
            .I(N__6255));
    CEMux I__928 (
            .O(N__6267),
            .I(N__6252));
    Span4Mux_v I__927 (
            .O(N__6264),
            .I(N__6249));
    Span4Mux_h I__926 (
            .O(N__6261),
            .I(N__6246));
    Span4Mux_h I__925 (
            .O(N__6258),
            .I(N__6243));
    LocalMux I__924 (
            .O(N__6255),
            .I(N__6240));
    LocalMux I__923 (
            .O(N__6252),
            .I(N__6237));
    Odrv4 I__922 (
            .O(N__6249),
            .I(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i ));
    Odrv4 I__921 (
            .O(N__6246),
            .I(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i ));
    Odrv4 I__920 (
            .O(N__6243),
            .I(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i ));
    Odrv4 I__919 (
            .O(N__6240),
            .I(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i ));
    Odrv4 I__918 (
            .O(N__6237),
            .I(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i ));
    InMux I__917 (
            .O(N__6226),
            .I(N__6205));
    InMux I__916 (
            .O(N__6225),
            .I(N__6205));
    InMux I__915 (
            .O(N__6224),
            .I(N__6202));
    InMux I__914 (
            .O(N__6223),
            .I(N__6199));
    InMux I__913 (
            .O(N__6222),
            .I(N__6196));
    InMux I__912 (
            .O(N__6221),
            .I(N__6187));
    InMux I__911 (
            .O(N__6220),
            .I(N__6187));
    InMux I__910 (
            .O(N__6219),
            .I(N__6187));
    InMux I__909 (
            .O(N__6218),
            .I(N__6187));
    InMux I__908 (
            .O(N__6217),
            .I(N__6182));
    InMux I__907 (
            .O(N__6216),
            .I(N__6182));
    InMux I__906 (
            .O(N__6215),
            .I(N__6177));
    InMux I__905 (
            .O(N__6214),
            .I(N__6177));
    InMux I__904 (
            .O(N__6213),
            .I(N__6174));
    InMux I__903 (
            .O(N__6212),
            .I(N__6169));
    InMux I__902 (
            .O(N__6211),
            .I(N__6169));
    InMux I__901 (
            .O(N__6210),
            .I(N__6166));
    LocalMux I__900 (
            .O(N__6205),
            .I(N__6161));
    LocalMux I__899 (
            .O(N__6202),
            .I(N__6161));
    LocalMux I__898 (
            .O(N__6199),
            .I(N__6156));
    LocalMux I__897 (
            .O(N__6196),
            .I(N__6156));
    LocalMux I__896 (
            .O(N__6187),
            .I(N__6143));
    LocalMux I__895 (
            .O(N__6182),
            .I(N__6143));
    LocalMux I__894 (
            .O(N__6177),
            .I(N__6143));
    LocalMux I__893 (
            .O(N__6174),
            .I(N__6143));
    LocalMux I__892 (
            .O(N__6169),
            .I(N__6143));
    LocalMux I__891 (
            .O(N__6166),
            .I(N__6143));
    Span4Mux_v I__890 (
            .O(N__6161),
            .I(N__6139));
    Span4Mux_v I__889 (
            .O(N__6156),
            .I(N__6136));
    Span4Mux_v I__888 (
            .O(N__6143),
            .I(N__6133));
    InMux I__887 (
            .O(N__6142),
            .I(N__6130));
    Sp12to4 I__886 (
            .O(N__6139),
            .I(N__6121));
    Sp12to4 I__885 (
            .O(N__6136),
            .I(N__6121));
    Sp12to4 I__884 (
            .O(N__6133),
            .I(N__6121));
    LocalMux I__883 (
            .O(N__6130),
            .I(N__6121));
    Odrv12 I__882 (
            .O(N__6121),
            .I(A_c_4));
    CascadeMux I__881 (
            .O(N__6118),
            .I(N__6113));
    CascadeMux I__880 (
            .O(N__6117),
            .I(N__6107));
    InMux I__879 (
            .O(N__6116),
            .I(N__6100));
    InMux I__878 (
            .O(N__6113),
            .I(N__6100));
    InMux I__877 (
            .O(N__6112),
            .I(N__6095));
    InMux I__876 (
            .O(N__6111),
            .I(N__6095));
    InMux I__875 (
            .O(N__6110),
            .I(N__6092));
    InMux I__874 (
            .O(N__6107),
            .I(N__6088));
    InMux I__873 (
            .O(N__6106),
            .I(N__6085));
    CascadeMux I__872 (
            .O(N__6105),
            .I(N__6081));
    LocalMux I__871 (
            .O(N__6100),
            .I(N__6073));
    LocalMux I__870 (
            .O(N__6095),
            .I(N__6073));
    LocalMux I__869 (
            .O(N__6092),
            .I(N__6073));
    InMux I__868 (
            .O(N__6091),
            .I(N__6070));
    LocalMux I__867 (
            .O(N__6088),
            .I(N__6067));
    LocalMux I__866 (
            .O(N__6085),
            .I(N__6064));
    InMux I__865 (
            .O(N__6084),
            .I(N__6061));
    InMux I__864 (
            .O(N__6081),
            .I(N__6058));
    CascadeMux I__863 (
            .O(N__6080),
            .I(N__6055));
    Span4Mux_v I__862 (
            .O(N__6073),
            .I(N__6052));
    LocalMux I__861 (
            .O(N__6070),
            .I(N__6046));
    Span4Mux_h I__860 (
            .O(N__6067),
            .I(N__6036));
    Span4Mux_v I__859 (
            .O(N__6064),
            .I(N__6036));
    LocalMux I__858 (
            .O(N__6061),
            .I(N__6036));
    LocalMux I__857 (
            .O(N__6058),
            .I(N__6036));
    InMux I__856 (
            .O(N__6055),
            .I(N__6033));
    Span4Mux_h I__855 (
            .O(N__6052),
            .I(N__6030));
    InMux I__854 (
            .O(N__6051),
            .I(N__6023));
    InMux I__853 (
            .O(N__6050),
            .I(N__6023));
    InMux I__852 (
            .O(N__6049),
            .I(N__6023));
    Span4Mux_v I__851 (
            .O(N__6046),
            .I(N__6020));
    InMux I__850 (
            .O(N__6045),
            .I(N__6017));
    Span4Mux_v I__849 (
            .O(N__6036),
            .I(N__6014));
    LocalMux I__848 (
            .O(N__6033),
            .I(N__6011));
    Sp12to4 I__847 (
            .O(N__6030),
            .I(N__6002));
    LocalMux I__846 (
            .O(N__6023),
            .I(N__6002));
    Sp12to4 I__845 (
            .O(N__6020),
            .I(N__6002));
    LocalMux I__844 (
            .O(N__6017),
            .I(N__6002));
    Span4Mux_h I__843 (
            .O(N__6014),
            .I(N__5997));
    Span4Mux_v I__842 (
            .O(N__6011),
            .I(N__5997));
    Span12Mux_h I__841 (
            .O(N__6002),
            .I(N__5994));
    Span4Mux_h I__840 (
            .O(N__5997),
            .I(N__5991));
    Span12Mux_v I__839 (
            .O(N__5994),
            .I(N__5988));
    Sp12to4 I__838 (
            .O(N__5991),
            .I(N__5985));
    Odrv12 I__837 (
            .O(N__5988),
            .I(A_c_2));
    Odrv12 I__836 (
            .O(N__5985),
            .I(A_c_2));
    InMux I__835 (
            .O(N__5980),
            .I(N__5972));
    InMux I__834 (
            .O(N__5979),
            .I(N__5972));
    InMux I__833 (
            .O(N__5978),
            .I(N__5969));
    CascadeMux I__832 (
            .O(N__5977),
            .I(N__5965));
    LocalMux I__831 (
            .O(N__5972),
            .I(N__5957));
    LocalMux I__830 (
            .O(N__5969),
            .I(N__5954));
    InMux I__829 (
            .O(N__5968),
            .I(N__5951));
    InMux I__828 (
            .O(N__5965),
            .I(N__5947));
    InMux I__827 (
            .O(N__5964),
            .I(N__5940));
    InMux I__826 (
            .O(N__5963),
            .I(N__5940));
    InMux I__825 (
            .O(N__5962),
            .I(N__5940));
    CascadeMux I__824 (
            .O(N__5961),
            .I(N__5936));
    CascadeMux I__823 (
            .O(N__5960),
            .I(N__5932));
    Span4Mux_v I__822 (
            .O(N__5957),
            .I(N__5928));
    Span4Mux_v I__821 (
            .O(N__5954),
            .I(N__5925));
    LocalMux I__820 (
            .O(N__5951),
            .I(N__5922));
    InMux I__819 (
            .O(N__5950),
            .I(N__5919));
    LocalMux I__818 (
            .O(N__5947),
            .I(N__5914));
    LocalMux I__817 (
            .O(N__5940),
            .I(N__5914));
    InMux I__816 (
            .O(N__5939),
            .I(N__5911));
    InMux I__815 (
            .O(N__5936),
            .I(N__5902));
    InMux I__814 (
            .O(N__5935),
            .I(N__5902));
    InMux I__813 (
            .O(N__5932),
            .I(N__5902));
    InMux I__812 (
            .O(N__5931),
            .I(N__5902));
    Odrv4 I__811 (
            .O(N__5928),
            .I(\U409_AUTOCONFIG.N_109 ));
    Odrv4 I__810 (
            .O(N__5925),
            .I(\U409_AUTOCONFIG.N_109 ));
    Odrv4 I__809 (
            .O(N__5922),
            .I(\U409_AUTOCONFIG.N_109 ));
    LocalMux I__808 (
            .O(N__5919),
            .I(\U409_AUTOCONFIG.N_109 ));
    Odrv4 I__807 (
            .O(N__5914),
            .I(\U409_AUTOCONFIG.N_109 ));
    LocalMux I__806 (
            .O(N__5911),
            .I(\U409_AUTOCONFIG.N_109 ));
    LocalMux I__805 (
            .O(N__5902),
            .I(\U409_AUTOCONFIG.N_109 ));
    CascadeMux I__804 (
            .O(N__5887),
            .I(N__5883));
    InMux I__803 (
            .O(N__5886),
            .I(N__5878));
    InMux I__802 (
            .O(N__5883),
            .I(N__5878));
    LocalMux I__801 (
            .O(N__5878),
            .I(N__5875));
    Odrv4 I__800 (
            .O(N__5875),
            .I(\U409_AUTOCONFIG.N_115 ));
    CascadeMux I__799 (
            .O(N__5872),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0_cascade_ ));
    InMux I__798 (
            .O(N__5869),
            .I(N__5866));
    LocalMux I__797 (
            .O(N__5866),
            .I(N__5862));
    InMux I__796 (
            .O(N__5865),
            .I(N__5859));
    Span4Mux_v I__795 (
            .O(N__5862),
            .I(N__5856));
    LocalMux I__794 (
            .O(N__5859),
            .I(N__5853));
    Odrv4 I__793 (
            .O(N__5856),
            .I(\U409_AUTOCONFIG.N_119 ));
    Odrv4 I__792 (
            .O(N__5853),
            .I(\U409_AUTOCONFIG.N_119 ));
    InMux I__791 (
            .O(N__5848),
            .I(N__5845));
    LocalMux I__790 (
            .O(N__5845),
            .I(N__5842));
    Odrv4 I__789 (
            .O(N__5842),
            .I(\U409_AUTOCONFIG.PR_OUTZ0Z_3 ));
    CascadeMux I__788 (
            .O(N__5839),
            .I(\U409_AUTOCONFIG.D_OUT_sm0_0_cascade_ ));
    IoInMux I__787 (
            .O(N__5836),
            .I(N__5833));
    LocalMux I__786 (
            .O(N__5833),
            .I(N__5830));
    Span4Mux_s1_v I__785 (
            .O(N__5830),
            .I(N__5827));
    Span4Mux_v I__784 (
            .O(N__5827),
            .I(N__5824));
    Span4Mux_v I__783 (
            .O(N__5824),
            .I(N__5821));
    Span4Mux_v I__782 (
            .O(N__5821),
            .I(N__5818));
    Odrv4 I__781 (
            .O(N__5818),
            .I(D_OUT_3));
    InMux I__780 (
            .O(N__5815),
            .I(N__5812));
    LocalMux I__779 (
            .O(N__5812),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ));
    InMux I__778 (
            .O(N__5809),
            .I(N__5806));
    LocalMux I__777 (
            .O(N__5806),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ));
    InMux I__776 (
            .O(N__5803),
            .I(N__5800));
    LocalMux I__775 (
            .O(N__5800),
            .I(\U409_AUTOCONFIG.LIDE_OUT_RNIBHMPZ0Z_3 ));
    InMux I__774 (
            .O(N__5797),
            .I(N__5794));
    LocalMux I__773 (
            .O(N__5794),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_0 ));
    CascadeMux I__772 (
            .O(N__5791),
            .I(\U409_AUTOCONFIG.PR_OUT_cnst_i_i_0_2_cascade_ ));
    InMux I__771 (
            .O(N__5788),
            .I(N__5785));
    LocalMux I__770 (
            .O(N__5785),
            .I(N__5782));
    Span4Mux_v I__769 (
            .O(N__5782),
            .I(N__5779));
    Odrv4 I__768 (
            .O(N__5779),
            .I(\U409_AUTOCONFIG.PR_OUTZ0Z_2 ));
    IoInMux I__767 (
            .O(N__5776),
            .I(N__5773));
    LocalMux I__766 (
            .O(N__5773),
            .I(N__5770));
    Span4Mux_s3_v I__765 (
            .O(N__5770),
            .I(N__5767));
    Sp12to4 I__764 (
            .O(N__5767),
            .I(N__5764));
    Span12Mux_h I__763 (
            .O(N__5764),
            .I(N__5761));
    Span12Mux_v I__762 (
            .O(N__5761),
            .I(N__5758));
    Odrv12 I__761 (
            .O(N__5758),
            .I(PORTSIZE_0_i));
    CascadeMux I__760 (
            .O(N__5755),
            .I(N__5751));
    CascadeMux I__759 (
            .O(N__5754),
            .I(N__5748));
    InMux I__758 (
            .O(N__5751),
            .I(N__5744));
    InMux I__757 (
            .O(N__5748),
            .I(N__5741));
    InMux I__756 (
            .O(N__5747),
            .I(N__5738));
    LocalMux I__755 (
            .O(N__5744),
            .I(N__5731));
    LocalMux I__754 (
            .O(N__5741),
            .I(N__5731));
    LocalMux I__753 (
            .O(N__5738),
            .I(N__5727));
    InMux I__752 (
            .O(N__5737),
            .I(N__5724));
    InMux I__751 (
            .O(N__5736),
            .I(N__5721));
    Span4Mux_v I__750 (
            .O(N__5731),
            .I(N__5718));
    InMux I__749 (
            .O(N__5730),
            .I(N__5715));
    Span4Mux_h I__748 (
            .O(N__5727),
            .I(N__5708));
    LocalMux I__747 (
            .O(N__5724),
            .I(N__5708));
    LocalMux I__746 (
            .O(N__5721),
            .I(N__5708));
    Sp12to4 I__745 (
            .O(N__5718),
            .I(N__5705));
    LocalMux I__744 (
            .O(N__5715),
            .I(N__5702));
    Sp12to4 I__743 (
            .O(N__5708),
            .I(N__5699));
    Span12Mux_h I__742 (
            .O(N__5705),
            .I(N__5694));
    Span12Mux_v I__741 (
            .O(N__5702),
            .I(N__5694));
    Span12Mux_v I__740 (
            .O(N__5699),
            .I(N__5691));
    Span12Mux_v I__739 (
            .O(N__5694),
            .I(N__5688));
    Odrv12 I__738 (
            .O(N__5691),
            .I(A_c_3));
    Odrv12 I__737 (
            .O(N__5688),
            .I(A_c_3));
    InMux I__736 (
            .O(N__5683),
            .I(N__5679));
    InMux I__735 (
            .O(N__5682),
            .I(N__5676));
    LocalMux I__734 (
            .O(N__5679),
            .I(N__5671));
    LocalMux I__733 (
            .O(N__5676),
            .I(N__5666));
    InMux I__732 (
            .O(N__5675),
            .I(N__5661));
    InMux I__731 (
            .O(N__5674),
            .I(N__5661));
    Span4Mux_v I__730 (
            .O(N__5671),
            .I(N__5658));
    InMux I__729 (
            .O(N__5670),
            .I(N__5655));
    InMux I__728 (
            .O(N__5669),
            .I(N__5652));
    Span4Mux_v I__727 (
            .O(N__5666),
            .I(N__5649));
    LocalMux I__726 (
            .O(N__5661),
            .I(N__5640));
    Sp12to4 I__725 (
            .O(N__5658),
            .I(N__5640));
    LocalMux I__724 (
            .O(N__5655),
            .I(N__5640));
    LocalMux I__723 (
            .O(N__5652),
            .I(N__5640));
    Span4Mux_h I__722 (
            .O(N__5649),
            .I(N__5637));
    Odrv12 I__721 (
            .O(N__5640),
            .I(A_c_6));
    Odrv4 I__720 (
            .O(N__5637),
            .I(A_c_6));
    CascadeMux I__719 (
            .O(N__5632),
            .I(\U409_AUTOCONFIG.N_109_cascade_ ));
    CascadeMux I__718 (
            .O(N__5629),
            .I(N__5625));
    InMux I__717 (
            .O(N__5628),
            .I(N__5620));
    InMux I__716 (
            .O(N__5625),
            .I(N__5620));
    LocalMux I__715 (
            .O(N__5620),
            .I(\U409_AUTOCONFIG.N_117 ));
    InMux I__714 (
            .O(N__5617),
            .I(N__5614));
    LocalMux I__713 (
            .O(N__5614),
            .I(N__5610));
    InMux I__712 (
            .O(N__5613),
            .I(N__5607));
    Odrv12 I__711 (
            .O(N__5610),
            .I(\U409_AUTOCONFIG.N_113 ));
    LocalMux I__710 (
            .O(N__5607),
            .I(\U409_AUTOCONFIG.N_113 ));
    InMux I__709 (
            .O(N__5602),
            .I(N__5599));
    LocalMux I__708 (
            .O(N__5599),
            .I(N__5596));
    Span4Mux_v I__707 (
            .O(N__5596),
            .I(N__5593));
    Sp12to4 I__706 (
            .O(N__5593),
            .I(N__5590));
    Span12Mux_h I__705 (
            .O(N__5590),
            .I(N__5587));
    Span12Mux_h I__704 (
            .O(N__5587),
            .I(N__5584));
    Span12Mux_v I__703 (
            .O(N__5584),
            .I(N__5581));
    Odrv12 I__702 (
            .O(N__5581),
            .I(AUTOBOOT_c));
    InMux I__701 (
            .O(N__5578),
            .I(N__5575));
    LocalMux I__700 (
            .O(N__5575),
            .I(N__5572));
    Odrv12 I__699 (
            .O(N__5572),
            .I(\U409_AUTOCONFIG.N_101 ));
    InMux I__698 (
            .O(N__5569),
            .I(N__5566));
    LocalMux I__697 (
            .O(N__5566),
            .I(\U409_AUTOCONFIG.PR_OUTZ0Z_1 ));
    InMux I__696 (
            .O(N__5563),
            .I(N__5560));
    LocalMux I__695 (
            .O(N__5560),
            .I(\U409_AUTOCONFIG.N_91 ));
    CascadeMux I__694 (
            .O(N__5557),
            .I(\U409_AUTOCONFIG.N_91_cascade_ ));
    InMux I__693 (
            .O(N__5554),
            .I(N__5551));
    LocalMux I__692 (
            .O(N__5551),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2 ));
    InMux I__691 (
            .O(N__5548),
            .I(N__5542));
    InMux I__690 (
            .O(N__5547),
            .I(N__5542));
    LocalMux I__689 (
            .O(N__5542),
            .I(\U409_AUTOCONFIG.N_216_3 ));
    CascadeMux I__688 (
            .O(N__5539),
            .I(\U409_AUTOCONFIG.LIDE_OUT_7_i_0_1_cascade_ ));
    InMux I__687 (
            .O(N__5536),
            .I(N__5533));
    LocalMux I__686 (
            .O(N__5533),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ));
    InMux I__685 (
            .O(N__5530),
            .I(N__5527));
    LocalMux I__684 (
            .O(N__5527),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ));
    InMux I__683 (
            .O(N__5524),
            .I(N__5521));
    LocalMux I__682 (
            .O(N__5521),
            .I(N__5518));
    Odrv4 I__681 (
            .O(N__5518),
            .I(\U409_AUTOCONFIG.LIDE_OUT_RNI7DMPZ0Z_1 ));
    InMux I__680 (
            .O(N__5515),
            .I(N__5511));
    CascadeMux I__679 (
            .O(N__5514),
            .I(N__5508));
    LocalMux I__678 (
            .O(N__5511),
            .I(N__5505));
    InMux I__677 (
            .O(N__5508),
            .I(N__5502));
    Odrv4 I__676 (
            .O(N__5505),
            .I(\U409_AUTOCONFIG.N_116 ));
    LocalMux I__675 (
            .O(N__5502),
            .I(\U409_AUTOCONFIG.N_116 ));
    InMux I__674 (
            .O(N__5497),
            .I(N__5494));
    LocalMux I__673 (
            .O(N__5494),
            .I(N__5489));
    InMux I__672 (
            .O(N__5493),
            .I(N__5486));
    InMux I__671 (
            .O(N__5492),
            .I(N__5483));
    Odrv4 I__670 (
            .O(N__5489),
            .I(\U409_AUTOCONFIG.N_89 ));
    LocalMux I__669 (
            .O(N__5486),
            .I(\U409_AUTOCONFIG.N_89 ));
    LocalMux I__668 (
            .O(N__5483),
            .I(\U409_AUTOCONFIG.N_89 ));
    InMux I__667 (
            .O(N__5476),
            .I(N__5473));
    LocalMux I__666 (
            .O(N__5473),
            .I(N__5470));
    Odrv4 I__665 (
            .O(N__5470),
            .I(U409_ADDRESS_DECODE_AUTOVECTOR_8));
    CascadeMux I__664 (
            .O(N__5467),
            .I(N__5464));
    InMux I__663 (
            .O(N__5464),
            .I(N__5461));
    LocalMux I__662 (
            .O(N__5461),
            .I(N__5458));
    Span4Mux_h I__661 (
            .O(N__5458),
            .I(N__5455));
    Span4Mux_v I__660 (
            .O(N__5455),
            .I(N__5452));
    Odrv4 I__659 (
            .O(N__5452),
            .I(U409_ADDRESS_DECODE_AUTOVECTOR_9));
    InMux I__658 (
            .O(N__5449),
            .I(N__5446));
    LocalMux I__657 (
            .O(N__5446),
            .I(U409_ADDRESS_DECODE_AUTOVECTOR_10));
    InMux I__656 (
            .O(N__5443),
            .I(N__5440));
    LocalMux I__655 (
            .O(N__5440),
            .I(\U409_AUTOCONFIG.N_99 ));
    CascadeMux I__654 (
            .O(N__5437),
            .I(N__5434));
    InMux I__653 (
            .O(N__5434),
            .I(N__5431));
    LocalMux I__652 (
            .O(N__5431),
            .I(N__5428));
    Odrv4 I__651 (
            .O(N__5428),
            .I(\U409_AUTOCONFIG.N_100 ));
    CascadeMux I__650 (
            .O(N__5425),
            .I(\U409_AUTOCONFIG.LIDE_OUT_RNI9FMPZ0Z_2_cascade_ ));
    IoInMux I__649 (
            .O(N__5422),
            .I(N__5419));
    LocalMux I__648 (
            .O(N__5419),
            .I(N__5416));
    Span4Mux_s2_v I__647 (
            .O(N__5416),
            .I(N__5413));
    Span4Mux_v I__646 (
            .O(N__5413),
            .I(N__5410));
    Span4Mux_v I__645 (
            .O(N__5410),
            .I(N__5407));
    Odrv4 I__644 (
            .O(N__5407),
            .I(D_OUT_2));
    IoInMux I__643 (
            .O(N__5404),
            .I(N__5401));
    LocalMux I__642 (
            .O(N__5401),
            .I(N__5398));
    Span4Mux_s1_v I__641 (
            .O(N__5398),
            .I(N__5395));
    Span4Mux_v I__640 (
            .O(N__5395),
            .I(N__5392));
    Span4Mux_v I__639 (
            .O(N__5392),
            .I(N__5389));
    Odrv4 I__638 (
            .O(N__5389),
            .I(D_OUT_1));
    InMux I__637 (
            .O(N__5386),
            .I(N__5383));
    LocalMux I__636 (
            .O(N__5383),
            .I(\U409_AUTOCONFIG.N_111 ));
    CascadeMux I__635 (
            .O(N__5380),
            .I(\U409_AUTOCONFIG.N_105_cascade_ ));
    InMux I__634 (
            .O(N__5377),
            .I(N__5374));
    LocalMux I__633 (
            .O(N__5374),
            .I(N__5370));
    InMux I__632 (
            .O(N__5373),
            .I(N__5367));
    Odrv4 I__631 (
            .O(N__5370),
            .I(PRO_BASE_1));
    LocalMux I__630 (
            .O(N__5367),
            .I(PRO_BASE_1));
    CascadeMux I__629 (
            .O(N__5362),
            .I(\U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1_cascade_ ));
    InMux I__628 (
            .O(N__5359),
            .I(N__5350));
    InMux I__627 (
            .O(N__5358),
            .I(N__5350));
    InMux I__626 (
            .O(N__5357),
            .I(N__5350));
    LocalMux I__625 (
            .O(N__5350),
            .I(\U409_AUTOCONFIG.CONFIGENn_1_sqmuxa ));
    InMux I__624 (
            .O(N__5347),
            .I(N__5344));
    LocalMux I__623 (
            .O(N__5344),
            .I(N__5341));
    Odrv4 I__622 (
            .O(N__5341),
            .I(\U409_AUTOCONFIG.LIDE_OUT_7_i_a4_0_0 ));
    CascadeMux I__621 (
            .O(N__5338),
            .I(\U409_AUTOCONFIG.N_216_3_cascade_ ));
    InMux I__620 (
            .O(N__5335),
            .I(N__5332));
    LocalMux I__619 (
            .O(N__5332),
            .I(\U409_AUTOCONFIG.N_108 ));
    CascadeMux I__618 (
            .O(N__5329),
            .I(\U409_AUTOCONFIG.N_108_cascade_ ));
    InMux I__617 (
            .O(N__5326),
            .I(N__5323));
    LocalMux I__616 (
            .O(N__5323),
            .I(\U409_ADDRESS_DECODE.N_59 ));
    CascadeMux I__615 (
            .O(N__5320),
            .I(\U409_ADDRESS_DECODE.N_59_cascade_ ));
    InMux I__614 (
            .O(N__5317),
            .I(N__5314));
    LocalMux I__613 (
            .O(N__5314),
            .I(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7 ));
    InMux I__612 (
            .O(N__5311),
            .I(N__5308));
    LocalMux I__611 (
            .O(N__5308),
            .I(N__5305));
    Span4Mux_v I__610 (
            .O(N__5305),
            .I(N__5301));
    InMux I__609 (
            .O(N__5304),
            .I(N__5298));
    Span4Mux_v I__608 (
            .O(N__5301),
            .I(N__5293));
    LocalMux I__607 (
            .O(N__5298),
            .I(N__5293));
    Span4Mux_h I__606 (
            .O(N__5293),
            .I(N__5290));
    Sp12to4 I__605 (
            .O(N__5290),
            .I(N__5287));
    Odrv12 I__604 (
            .O(N__5287),
            .I(TT_c_1));
    InMux I__603 (
            .O(N__5284),
            .I(N__5281));
    LocalMux I__602 (
            .O(N__5281),
            .I(N__5278));
    Span4Mux_v I__601 (
            .O(N__5278),
            .I(N__5274));
    InMux I__600 (
            .O(N__5277),
            .I(N__5271));
    Span4Mux_h I__599 (
            .O(N__5274),
            .I(N__5268));
    LocalMux I__598 (
            .O(N__5271),
            .I(N__5265));
    Sp12to4 I__597 (
            .O(N__5268),
            .I(N__5260));
    Span12Mux_h I__596 (
            .O(N__5265),
            .I(N__5260));
    Odrv12 I__595 (
            .O(N__5260),
            .I(TT_c_0));
    CascadeMux I__594 (
            .O(N__5257),
            .I(N__5254));
    InMux I__593 (
            .O(N__5254),
            .I(N__5251));
    LocalMux I__592 (
            .O(N__5251),
            .I(N__5248));
    Span4Mux_v I__591 (
            .O(N__5248),
            .I(N__5245));
    Span4Mux_v I__590 (
            .O(N__5245),
            .I(N__5242));
    IoSpan4Mux I__589 (
            .O(N__5242),
            .I(N__5239));
    Odrv4 I__588 (
            .O(N__5239),
            .I(TM_c_2));
    IoInMux I__587 (
            .O(N__5236),
            .I(N__5233));
    LocalMux I__586 (
            .O(N__5233),
            .I(N__5228));
    IoInMux I__585 (
            .O(N__5232),
            .I(N__5225));
    IoInMux I__584 (
            .O(N__5231),
            .I(N__5222));
    IoSpan4Mux I__583 (
            .O(N__5228),
            .I(N__5214));
    LocalMux I__582 (
            .O(N__5225),
            .I(N__5214));
    LocalMux I__581 (
            .O(N__5222),
            .I(N__5214));
    IoInMux I__580 (
            .O(N__5221),
            .I(N__5211));
    IoSpan4Mux I__579 (
            .O(N__5214),
            .I(N__5208));
    LocalMux I__578 (
            .O(N__5211),
            .I(N__5205));
    Span4Mux_s3_v I__577 (
            .O(N__5208),
            .I(N__5200));
    Span4Mux_s3_v I__576 (
            .O(N__5205),
            .I(N__5200));
    Span4Mux_v I__575 (
            .O(N__5200),
            .I(N__5197));
    Odrv4 I__574 (
            .O(N__5197),
            .I(D_1_i));
    IoInMux I__573 (
            .O(N__5194),
            .I(N__5191));
    LocalMux I__572 (
            .O(N__5191),
            .I(N__5188));
    Span4Mux_s1_v I__571 (
            .O(N__5188),
            .I(N__5185));
    Sp12to4 I__570 (
            .O(N__5185),
            .I(N__5181));
    CascadeMux I__569 (
            .O(N__5184),
            .I(N__5178));
    Span12Mux_h I__568 (
            .O(N__5181),
            .I(N__5175));
    InMux I__567 (
            .O(N__5178),
            .I(N__5172));
    Odrv12 I__566 (
            .O(N__5175),
            .I(CONFIGENn_c));
    LocalMux I__565 (
            .O(N__5172),
            .I(CONFIGENn_c));
    InMux I__564 (
            .O(N__5167),
            .I(N__5163));
    InMux I__563 (
            .O(N__5166),
            .I(N__5160));
    LocalMux I__562 (
            .O(N__5163),
            .I(PRO_BASE_2));
    LocalMux I__561 (
            .O(N__5160),
            .I(PRO_BASE_2));
    InMux I__560 (
            .O(N__5155),
            .I(N__5151));
    InMux I__559 (
            .O(N__5154),
            .I(N__5148));
    LocalMux I__558 (
            .O(N__5151),
            .I(PRO_BASE_0));
    LocalMux I__557 (
            .O(N__5148),
            .I(PRO_BASE_0));
    IoInMux I__556 (
            .O(N__5143),
            .I(N__5140));
    LocalMux I__555 (
            .O(N__5140),
            .I(N__5137));
    Span4Mux_s0_v I__554 (
            .O(N__5137),
            .I(N__5134));
    Sp12to4 I__553 (
            .O(N__5134),
            .I(N__5131));
    Span12Mux_h I__552 (
            .O(N__5131),
            .I(N__5128));
    Span12Mux_v I__551 (
            .O(N__5128),
            .I(N__5125));
    Odrv12 I__550 (
            .O(N__5125),
            .I(U409_ADDRESS_DECODE_un1_BPRO_ENn_i));
    InMux I__549 (
            .O(N__5122),
            .I(N__5117));
    InMux I__548 (
            .O(N__5121),
            .I(N__5114));
    InMux I__547 (
            .O(N__5120),
            .I(N__5111));
    LocalMux I__546 (
            .O(N__5117),
            .I(N__5108));
    LocalMux I__545 (
            .O(N__5114),
            .I(N__5103));
    LocalMux I__544 (
            .O(N__5111),
            .I(N__5103));
    Sp12to4 I__543 (
            .O(N__5108),
            .I(N__5100));
    Sp12to4 I__542 (
            .O(N__5103),
            .I(N__5097));
    Span12Mux_v I__541 (
            .O(N__5100),
            .I(N__5094));
    Span12Mux_v I__540 (
            .O(N__5097),
            .I(N__5091));
    Odrv12 I__539 (
            .O(N__5094),
            .I(A_c_29));
    Odrv12 I__538 (
            .O(N__5091),
            .I(A_c_29));
    CascadeMux I__537 (
            .O(N__5086),
            .I(\U409_ADDRESS_DECODE.N_26_cascade_ ));
    InMux I__536 (
            .O(N__5083),
            .I(N__5080));
    LocalMux I__535 (
            .O(N__5080),
            .I(\U409_ADDRESS_DECODE.m54Z0Z_1 ));
    InMux I__534 (
            .O(N__5077),
            .I(N__5074));
    LocalMux I__533 (
            .O(N__5074),
            .I(N__5071));
    Span4Mux_h I__532 (
            .O(N__5071),
            .I(N__5068));
    Odrv4 I__531 (
            .O(N__5068),
            .I(\U409_AUTOCONFIG.un1_A_13Z0Z_3 ));
    InMux I__530 (
            .O(N__5065),
            .I(N__5062));
    LocalMux I__529 (
            .O(N__5062),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a4_0_0Z0Z_0 ));
    InMux I__528 (
            .O(N__5059),
            .I(N__5056));
    LocalMux I__527 (
            .O(N__5056),
            .I(N__5052));
    InMux I__526 (
            .O(N__5055),
            .I(N__5049));
    Span4Mux_v I__525 (
            .O(N__5052),
            .I(N__5044));
    LocalMux I__524 (
            .O(N__5049),
            .I(N__5044));
    Span4Mux_h I__523 (
            .O(N__5044),
            .I(N__5040));
    InMux I__522 (
            .O(N__5043),
            .I(N__5037));
    Span4Mux_v I__521 (
            .O(N__5040),
            .I(N__5032));
    LocalMux I__520 (
            .O(N__5037),
            .I(N__5032));
    Span4Mux_h I__519 (
            .O(N__5032),
            .I(N__5029));
    Span4Mux_v I__518 (
            .O(N__5029),
            .I(N__5026));
    Odrv4 I__517 (
            .O(N__5026),
            .I(A_c_30));
    InMux I__516 (
            .O(N__5023),
            .I(N__5019));
    CascadeMux I__515 (
            .O(N__5022),
            .I(N__5016));
    LocalMux I__514 (
            .O(N__5019),
            .I(N__5013));
    InMux I__513 (
            .O(N__5016),
            .I(N__5009));
    Span4Mux_h I__512 (
            .O(N__5013),
            .I(N__5006));
    InMux I__511 (
            .O(N__5012),
            .I(N__5003));
    LocalMux I__510 (
            .O(N__5009),
            .I(N__5000));
    Span4Mux_v I__509 (
            .O(N__5006),
            .I(N__4995));
    LocalMux I__508 (
            .O(N__5003),
            .I(N__4995));
    Span12Mux_h I__507 (
            .O(N__5000),
            .I(N__4992));
    Span4Mux_h I__506 (
            .O(N__4995),
            .I(N__4989));
    Span12Mux_v I__505 (
            .O(N__4992),
            .I(N__4986));
    Span4Mux_v I__504 (
            .O(N__4989),
            .I(N__4983));
    Odrv12 I__503 (
            .O(N__4986),
            .I(A_c_31));
    Odrv4 I__502 (
            .O(N__4983),
            .I(A_c_31));
    InMux I__501 (
            .O(N__4978),
            .I(N__4975));
    LocalMux I__500 (
            .O(N__4975),
            .I(\U409_ADDRESS_DECODE.m12Z0Z_5 ));
    CascadeMux I__499 (
            .O(N__4972),
            .I(\U409_ADDRESS_DECODE.m12Z0Z_0_cascade_ ));
    InMux I__498 (
            .O(N__4969),
            .I(N__4966));
    LocalMux I__497 (
            .O(N__4966),
            .I(\U409_AUTOCONFIG.un1_A_13Z0Z_1 ));
    CascadeMux I__496 (
            .O(N__4963),
            .I(N__4960));
    InMux I__495 (
            .O(N__4960),
            .I(N__4956));
    InMux I__494 (
            .O(N__4959),
            .I(N__4953));
    LocalMux I__493 (
            .O(N__4956),
            .I(N__4950));
    LocalMux I__492 (
            .O(N__4953),
            .I(N__4947));
    Sp12to4 I__491 (
            .O(N__4950),
            .I(N__4944));
    Span4Mux_v I__490 (
            .O(N__4947),
            .I(N__4941));
    Span12Mux_v I__489 (
            .O(N__4944),
            .I(N__4938));
    Span4Mux_h I__488 (
            .O(N__4941),
            .I(N__4935));
    Odrv12 I__487 (
            .O(N__4938),
            .I(A_c_25));
    Odrv4 I__486 (
            .O(N__4935),
            .I(A_c_25));
    CascadeMux I__485 (
            .O(N__4930),
            .I(N__4927));
    InMux I__484 (
            .O(N__4927),
            .I(N__4923));
    InMux I__483 (
            .O(N__4926),
            .I(N__4920));
    LocalMux I__482 (
            .O(N__4923),
            .I(N__4917));
    LocalMux I__481 (
            .O(N__4920),
            .I(N__4914));
    Span4Mux_v I__480 (
            .O(N__4917),
            .I(N__4911));
    Sp12to4 I__479 (
            .O(N__4914),
            .I(N__4908));
    Span4Mux_v I__478 (
            .O(N__4911),
            .I(N__4905));
    Span12Mux_v I__477 (
            .O(N__4908),
            .I(N__4902));
    Span4Mux_h I__476 (
            .O(N__4905),
            .I(N__4899));
    Odrv12 I__475 (
            .O(N__4902),
            .I(A_c_24));
    Odrv4 I__474 (
            .O(N__4899),
            .I(A_c_24));
    InMux I__473 (
            .O(N__4894),
            .I(N__4891));
    LocalMux I__472 (
            .O(N__4891),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_3 ));
    CascadeMux I__471 (
            .O(N__4888),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4_cascade_ ));
    InMux I__470 (
            .O(N__4885),
            .I(N__4879));
    InMux I__469 (
            .O(N__4884),
            .I(N__4879));
    LocalMux I__468 (
            .O(N__4879),
            .I(N__4876));
    Span4Mux_v I__467 (
            .O(N__4876),
            .I(N__4873));
    Sp12to4 I__466 (
            .O(N__4873),
            .I(N__4870));
    Odrv12 I__465 (
            .O(N__4870),
            .I(A_c_27));
    CascadeMux I__464 (
            .O(N__4867),
            .I(N__4863));
    InMux I__463 (
            .O(N__4866),
            .I(N__4860));
    InMux I__462 (
            .O(N__4863),
            .I(N__4857));
    LocalMux I__461 (
            .O(N__4860),
            .I(N__4854));
    LocalMux I__460 (
            .O(N__4857),
            .I(N__4851));
    Span4Mux_v I__459 (
            .O(N__4854),
            .I(N__4846));
    Span4Mux_v I__458 (
            .O(N__4851),
            .I(N__4846));
    Span4Mux_v I__457 (
            .O(N__4846),
            .I(N__4843));
    Span4Mux_v I__456 (
            .O(N__4843),
            .I(N__4840));
    Span4Mux_h I__455 (
            .O(N__4840),
            .I(N__4837));
    Odrv4 I__454 (
            .O(N__4837),
            .I(A_c_28));
    InMux I__453 (
            .O(N__4834),
            .I(N__4830));
    InMux I__452 (
            .O(N__4833),
            .I(N__4827));
    LocalMux I__451 (
            .O(N__4830),
            .I(N__4824));
    LocalMux I__450 (
            .O(N__4827),
            .I(N__4821));
    Span4Mux_v I__449 (
            .O(N__4824),
            .I(N__4818));
    Span4Mux_v I__448 (
            .O(N__4821),
            .I(N__4815));
    Span4Mux_v I__447 (
            .O(N__4818),
            .I(N__4812));
    Span4Mux_v I__446 (
            .O(N__4815),
            .I(N__4809));
    Span4Mux_h I__445 (
            .O(N__4812),
            .I(N__4806));
    Span4Mux_h I__444 (
            .O(N__4809),
            .I(N__4803));
    Odrv4 I__443 (
            .O(N__4806),
            .I(A_c_26));
    Odrv4 I__442 (
            .O(N__4803),
            .I(A_c_26));
    IoInMux I__441 (
            .O(N__4798),
            .I(N__4795));
    LocalMux I__440 (
            .O(N__4795),
            .I(N__4792));
    IoSpan4Mux I__439 (
            .O(N__4792),
            .I(N__4789));
    Sp12to4 I__438 (
            .O(N__4789),
            .I(N__4786));
    Span12Mux_s1_h I__437 (
            .O(N__4786),
            .I(N__4783));
    Span12Mux_v I__436 (
            .O(N__4783),
            .I(N__4780));
    Odrv12 I__435 (
            .O(N__4780),
            .I(PPIO_c));
    IoInMux I__434 (
            .O(N__4777),
            .I(N__4774));
    LocalMux I__433 (
            .O(N__4774),
            .I(N__4771));
    Span12Mux_s2_h I__432 (
            .O(N__4771),
            .I(N__4768));
    Span12Mux_v I__431 (
            .O(N__4768),
            .I(N__4765));
    Odrv12 I__430 (
            .O(N__4765),
            .I(SPIO_c));
    ClkMux I__429 (
            .O(N__4762),
            .I(N__4723));
    ClkMux I__428 (
            .O(N__4761),
            .I(N__4723));
    ClkMux I__427 (
            .O(N__4760),
            .I(N__4723));
    ClkMux I__426 (
            .O(N__4759),
            .I(N__4723));
    ClkMux I__425 (
            .O(N__4758),
            .I(N__4723));
    ClkMux I__424 (
            .O(N__4757),
            .I(N__4723));
    ClkMux I__423 (
            .O(N__4756),
            .I(N__4723));
    ClkMux I__422 (
            .O(N__4755),
            .I(N__4723));
    ClkMux I__421 (
            .O(N__4754),
            .I(N__4723));
    ClkMux I__420 (
            .O(N__4753),
            .I(N__4723));
    ClkMux I__419 (
            .O(N__4752),
            .I(N__4723));
    ClkMux I__418 (
            .O(N__4751),
            .I(N__4723));
    ClkMux I__417 (
            .O(N__4750),
            .I(N__4723));
    GlobalMux I__416 (
            .O(N__4723),
            .I(CLK80_OUT));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .I(N__4762));
    INV \INVU409_TRANSFER_ACK.LASTCLK_1C  (
            .O(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .I(N__4760));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .I(N__4758));
    INV \INVU409_TRANSFER_ACK.CIA_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .I(N__4755));
    INV \INVU409_TRANSFER_ACK.ROMENnC  (
            .O(\INVU409_TRANSFER_ACK.ROMENnC_net ),
            .I(N__4757));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .I(N__4754));
    INV \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC  (
            .O(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .I(N__4753));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net ),
            .I(N__4751));
    INV \INVU409_TRANSFER_ACK.TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .I(N__4750));
    INV \INVU409_AUTOCONFIG.AC_TACKC  (
            .O(\INVU409_AUTOCONFIG.AC_TACKC_net ),
            .I(N__11161));
    INV \INVU409_AUTOCONFIG.STATE_1C  (
            .O(\INVU409_AUTOCONFIG.STATE_1C_net ),
            .I(N__11165));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_EN_nerC  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_EN_nerC_net ),
            .I(N__4752));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net ),
            .I(N__4759));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .I(N__4756));
    INV \INVU409_AUTOCONFIG.BRIDGE_BASE_5C  (
            .O(\INVU409_AUTOCONFIG.BRIDGE_BASE_5C_net ),
            .I(N__11171));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .I(N__4761));
    INV \INVU409_AUTOCONFIG.BRIDGE_BASE_4C  (
            .O(\INVU409_AUTOCONFIG.BRIDGE_BASE_4C_net ),
            .I(N__11170));
    INV \INVU409_AUTOCONFIG.BRIDGE_BASE_0C  (
            .O(\INVU409_AUTOCONFIG.BRIDGE_BASE_0C_net ),
            .I(N__11174));
    INV \INVU409_AUTOCONFIG.LIDE_BASE_1C  (
            .O(\INVU409_AUTOCONFIG.LIDE_BASE_1C_net ),
            .I(N__11181));
    INV \INVU409_AUTOCONFIG.LIDE_OUT_2C  (
            .O(\INVU409_AUTOCONFIG.LIDE_OUT_2C_net ),
            .I(N__11173));
    INV \INVU409_AUTOCONFIG.BRIDGE_OUT_3C  (
            .O(\INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net ),
            .I(N__11180));
    INV \INVU409_AUTOCONFIG.BRIDGE_OUT_1C  (
            .O(\INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net ),
            .I(N__11172));
    INV \INVU409_AUTOCONFIG.PR_OUT_1C  (
            .O(\INVU409_AUTOCONFIG.PR_OUT_1C_net ),
            .I(N__11179));
    INV \INVU409_AUTOCONFIG.LIDE_OUT_0C  (
            .O(\INVU409_AUTOCONFIG.LIDE_OUT_0C_net ),
            .I(N__11182));
    INV \INVU409_AUTOCONFIG.LIDE_CONFC  (
            .O(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .I(N__11183));
    INV \INVU409_AUTOCONFIG.CONFIGENnC  (
            .O(\INVU409_AUTOCONFIG.CONFIGENnC_net ),
            .I(N__11187));
    defparam IN_MUX_bfv_14_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_6_0_));
    defparam IN_MUX_bfv_14_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_7_0_ (
            .carryinitin(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .carryinitout(bfn_14_7_0_));
    defparam IN_MUX_bfv_17_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_5_0_));
    defparam IN_MUX_bfv_17_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_6_0_ (
            .carryinitin(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .carryinitout(bfn_17_6_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_12_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__9538),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.m12_5_LC_1_15_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.m12_5_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.m12_5_LC_1_15_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.m12_5_LC_1_15_4  (
            .in0(N__4885),
            .in1(N__5043),
            .in2(N__4930),
            .in3(N__4866),
            .lcout(\U409_ADDRESS_DECODE.m12Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_1_15_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_1_15_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_1_15_6  (
            .in0(N__4884),
            .in1(N__5120),
            .in2(N__4867),
            .in3(N__4833),
            .lcout(U409_ADDRESS_DECODE_AUTOVECTOR_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_13_1_LC_2_10_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_13_1_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_13_1_LC_2_10_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_AUTOCONFIG.un1_A_13_1_LC_2_10_7  (
            .in0(N__5730),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5682),
            .lcout(\U409_AUTOCONFIG.un1_A_13Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.m12_0_LC_2_15_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.m12_0_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.m12_0_LC_2_15_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_ADDRESS_DECODE.m12_0_LC_2_15_1  (
            .in0(N__4834),
            .in1(N__11809),
            .in2(_gnd_net_),
            .in3(N__5121),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.m12Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.m12_LC_2_15_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.m12_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.m12_LC_2_15_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_ADDRESS_DECODE.m12_LC_2_15_2  (
            .in0(N__5012),
            .in1(N__4978),
            .in2(N__4972),
            .in3(N__4959),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACE ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_3_7_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_3_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_3_7_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_3_7_6  (
            .in0(N__7735),
            .in1(N__9974),
            .in2(N__9283),
            .in3(N__7805),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACE_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.m1_LC_3_9_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.m1_LC_3_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.m1_LC_3_9_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.m1_LC_3_9_7  (
            .in0(N__10174),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9915),
            .lcout(\U409_ADDRESS_DECODE.N_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_13_3_LC_3_10_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_13_3_LC_3_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_13_3_LC_3_10_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_AUTOCONFIG.un1_A_13_3_LC_3_10_5  (
            .in0(N__6900),
            .in1(N__7044),
            .in2(N__6080),
            .in3(N__4969),
            .lcout(\U409_AUTOCONFIG.un1_A_13Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_3_11_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_3_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_3_11_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_3_11_4  (
            .in0(N__9082),
            .in1(N__8477),
            .in2(N__4963),
            .in3(N__4926),
            .lcout(U409_ADDRESS_DECODE_AUTOVECTOR_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_3_LC_5_5_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_3_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_3_LC_5_5_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_3_LC_5_5_0  (
            .in0(N__7710),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7809),
            .lcout(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_4_LC_5_6_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_4_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_4_LC_5_6_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_4_LC_5_6_0  (
            .in0(N__9092),
            .in1(N__9698),
            .in2(N__10018),
            .in3(N__10100),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_5_6_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_5_6_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_5_6_1  (
            .in0(N__4894),
            .in1(N__9375),
            .in2(N__4888),
            .in3(N__9284),
            .lcout(AUTOCONFIG_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.m13_LC_5_7_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.m13_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.m13_LC_5_7_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.m13_LC_5_7_0  (
            .in0(N__9352),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10194),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACE_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BPRO_ENn_i_LC_5_7_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BPRO_ENn_i_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BPRO_ENn_i_LC_5_7_5 .LUT_INIT=16'b0111110111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BPRO_ENn_i_LC_5_7_5  (
            .in0(N__5083),
            .in1(N__5167),
            .in2(N__5022),
            .in3(N__7631),
            .lcout(U409_ADDRESS_DECODE_un1_BPRO_ENn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.m47_LC_5_8_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.m47_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.m47_LC_5_8_0 .LUT_INIT=16'b0111011110111011;
    LogicCell40 \U409_ADDRESS_DECODE.m47_LC_5_8_0  (
            .in0(N__5122),
            .in1(N__11876),
            .in2(_gnd_net_),
            .in3(N__5155),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.N_26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.m54_1_LC_5_8_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.m54_1_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.m54_1_LC_5_8_1 .LUT_INIT=16'b0000101000000101;
    LogicCell40 \U409_ADDRESS_DECODE.m54_1_LC_5_8_1  (
            .in0(N__5059),
            .in1(_gnd_net_),
            .in2(N__5086),
            .in3(N__5377),
            .lcout(\U409_ADDRESS_DECODE.m54Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_13_LC_5_9_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_13_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_13_LC_5_9_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U409_AUTOCONFIG.un1_A_13_LC_5_9_0  (
            .in0(N__6223),
            .in1(N__7017),
            .in2(_gnd_net_),
            .in3(N__5077),
            .lcout(\U409_AUTOCONFIG.un1_AZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a4_0_0_LC_5_10_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a4_0_0_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a4_0_0_LC_5_10_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a4_0_0_LC_5_10_0  (
            .in0(N__5065),
            .in1(N__5747),
            .in2(N__5514),
            .in3(N__6911),
            .lcout(\U409_AUTOCONFIG.N_104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a4_0_0_0_LC_5_10_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a4_0_0_0_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a4_0_0_0_LC_5_10_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a4_0_0_0_LC_5_10_3  (
            .in0(N__7016),
            .in1(N__7045),
            .in2(_gnd_net_),
            .in3(N__5683),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a4_0_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_1_3_LC_5_10_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_1_3_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_1_3_LC_5_10_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_1_3_LC_5_10_7  (
            .in0(N__6222),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6091),
            .lcout(\U409_AUTOCONFIG.N_116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_0_LC_5_11_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_0_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_0_LC_5_11_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_10_0_LC_5_11_3  (
            .in0(N__5055),
            .in1(N__5317),
            .in2(_gnd_net_),
            .in3(N__5023),
            .lcout(U409_ADDRESS_DECODE_AUTOVECTOR_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_3_0_LC_5_11_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_3_0_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_3_0_LC_5_11_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_3_0_LC_5_11_5  (
            .in0(N__7069),
            .in1(N__5669),
            .in2(_gnd_net_),
            .in3(N__5736),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_7_i_a4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_5_11_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_5_11_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_LC_5_11_6  (
            .in0(N__9867),
            .in1(N__5326),
            .in2(N__8495),
            .in3(N__8542),
            .lcout(CIA_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.m3_LC_5_12_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.m3_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.m3_LC_5_12_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_ADDRESS_DECODE.m3_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(N__9683),
            .in2(_gnd_net_),
            .in3(N__10045),
            .lcout(\U409_ADDRESS_DECODE.N_59 ),
            .ltout(\U409_ADDRESS_DECODE.N_59_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_5_12_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_5_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_5_12_2  (
            .in0(N__5311),
            .in1(N__5284),
            .in2(N__5320),
            .in3(N__11883),
            .lcout(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.m41_LC_5_17_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.m41_LC_5_17_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.m41_LC_5_17_7 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_ADDRESS_DECODE.m41_LC_5_17_7  (
            .in0(N__5304),
            .in1(N__5277),
            .in2(N__5257),
            .in3(N__11887),
            .lcout(\U409_ADDRESS_DECODE.N_58_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_6_6_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_6_6_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_ADDRESS_DECODE.D_1_i_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__8390),
            .in2(_gnd_net_),
            .in3(N__8868),
            .lcout(D_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_6_7_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_6_7_1 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_6_7_1 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_AUTOCONFIG.CONFIGENn_LC_6_7_1  (
            .in0(N__7456),
            .in1(N__6533),
            .in2(N__5184),
            .in3(N__6624),
            .lcout(CONFIGENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.CONFIGENnC_net ),
            .ce(),
            .sr(N__11395));
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_6_8_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_6_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_6_8_1 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_LC_6_8_1  (
            .in0(N__7449),
            .in1(N__6539),
            .in2(_gnd_net_),
            .in3(N__6617),
            .lcout(\U409_AUTOCONFIG.LIDE_CONFZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .ce(),
            .sr(N__11394));
    defparam \U409_AUTOCONFIG.PRO_BASE_2_LC_6_8_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PRO_BASE_2_LC_6_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.PRO_BASE_2_LC_6_8_3 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U409_AUTOCONFIG.PRO_BASE_2_LC_6_8_3  (
            .in0(N__5359),
            .in1(N__7906),
            .in2(N__8062),
            .in3(N__5166),
            .lcout(PRO_BASE_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .ce(),
            .sr(N__11394));
    defparam \U409_AUTOCONFIG.PRO_BASE_0_LC_6_8_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PRO_BASE_0_LC_6_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.PRO_BASE_0_LC_6_8_6 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U409_AUTOCONFIG.PRO_BASE_0_LC_6_8_6  (
            .in0(N__7904),
            .in1(N__5154),
            .in2(N__8152),
            .in3(N__5357),
            .lcout(PRO_BASE_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .ce(),
            .sr(N__11394));
    defparam \U409_AUTOCONFIG.PRO_BASE_1_LC_6_8_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PRO_BASE_1_LC_6_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.PRO_BASE_1_LC_6_8_7 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U409_AUTOCONFIG.PRO_BASE_1_LC_6_8_7  (
            .in0(N__5358),
            .in1(N__7905),
            .in2(N__6754),
            .in3(N__5373),
            .lcout(PRO_BASE_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .ce(),
            .sr(N__11394));
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_1_1_LC_6_9_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_1_1_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_1_1_LC_6_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_RNO_1_1_LC_6_9_0  (
            .in0(_gnd_net_),
            .in1(N__5980),
            .in2(_gnd_net_),
            .in3(N__6849),
            .lcout(\U409_AUTOCONFIG.N_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_6_9_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_6_9_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_6_9_1  (
            .in0(N__5979),
            .in1(N__6215),
            .in2(N__6886),
            .in3(N__6112),
            .lcout(\U409_AUTOCONFIG.N_100 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNIDEFO1_0_LC_6_9_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNIDEFO1_0_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNIDEFO1_0_LC_6_9_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNIDEFO1_0_LC_6_9_4  (
            .in0(N__7467),
            .in1(N__8904),
            .in2(_gnd_net_),
            .in3(N__8778),
            .lcout(\U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1 ),
            .ltout(\U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_LC_6_9_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_LC_6_9_5 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_LC_6_9_5  (
            .in0(_gnd_net_),
            .in1(N__7451),
            .in2(N__5362),
            .in3(N__6518),
            .lcout(\U409_AUTOCONFIG.CONFIGENn_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_6_9_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_6_9_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_6_9_7  (
            .in0(N__5347),
            .in1(N__6111),
            .in2(N__6885),
            .in3(N__6214),
            .lcout(\U409_AUTOCONFIG.N_99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_14_2_0_a2_LC_6_10_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_14_2_0_a2_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_14_2_0_a2_LC_6_10_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_AUTOCONFIG.un1_A_14_2_0_a2_LC_6_10_3  (
            .in0(N__6213),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6110),
            .lcout(\U409_AUTOCONFIG.N_216_3 ),
            .ltout(\U409_AUTOCONFIG.N_216_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_o4_2_LC_6_10_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_o4_2_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_o4_2_LC_6_10_4 .LUT_INIT=16'b0011001110110011;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_cnst_i_i_o4_2_LC_6_10_4  (
            .in0(N__5335),
            .in1(N__11875),
            .in2(N__5338),
            .in3(N__6912),
            .lcout(\U409_AUTOCONFIG.N_89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_2_3_LC_6_11_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_2_3_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_2_3_LC_6_11_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_2_3_LC_6_11_3  (
            .in0(N__6997),
            .in1(N__7073),
            .in2(_gnd_net_),
            .in3(N__5670),
            .lcout(\U409_AUTOCONFIG.N_108 ),
            .ltout(\U409_AUTOCONFIG.N_108_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_3_LC_6_11_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_3_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_3_LC_6_11_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_3_LC_6_11_4  (
            .in0(N__6210),
            .in1(N__5737),
            .in2(N__5329),
            .in3(N__6045),
            .lcout(\U409_AUTOCONFIG.N_119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_AUTOVECTOR_LC_6_11_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_AUTOVECTOR_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_AUTOVECTOR_LC_6_11_7 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \U409_TRANSFER_ACK.un1_AUTOVECTOR_LC_6_11_7  (
            .in0(N__5476),
            .in1(N__7123),
            .in2(N__5467),
            .in3(N__5449),
            .lcout(\U409_TRANSFER_ACK.un1_AUTOVECTOR_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_7_8_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_7_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_7_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_0_LC_7_8_0  (
            .in0(N__5563),
            .in1(N__5443),
            .in2(N__5437),
            .in3(N__5578),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_0C_net ),
            .ce(N__6279),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI9FMP_2_LC_7_8_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI9FMP_2_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI9FMP_2_LC_7_8_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNI9FMP_2_LC_7_8_1  (
            .in0(N__7448),
            .in1(N__6337),
            .in2(_gnd_net_),
            .in3(N__5554),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.LIDE_OUT_RNI9FMPZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_RNIVV912_2_LC_7_8_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_RNIVV912_2_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_RNIVV912_2_LC_7_8_2 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_RNIVV912_2_LC_7_8_2  (
            .in0(N__5788),
            .in1(N__6382),
            .in2(N__5425),
            .in3(N__7635),
            .lcout(D_OUT_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_RNISS912_1_LC_7_8_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_RNISS912_1_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_RNISS912_1_LC_7_8_3 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_RNISS912_1_LC_7_8_3  (
            .in0(N__6381),
            .in1(N__5569),
            .in2(N__7636),
            .in3(N__5524),
            .lcout(D_OUT_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_0_LC_7_8_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_0_LC_7_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.PR_OUT_0_LC_7_8_4 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_0_LC_7_8_4  (
            .in0(N__5497),
            .in1(N__6307),
            .in2(N__5977),
            .in3(N__5617),
            .lcout(\U409_AUTOCONFIG.PR_OUTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_0C_net ),
            .ce(N__6279),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_0_o2_2_LC_7_9_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_0_o2_2_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_0_o2_2_LC_7_9_1 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_7_0_o2_2_LC_7_9_1  (
            .in0(N__5962),
            .in1(N__6218),
            .in2(N__6118),
            .in3(N__5865),
            .lcout(\U409_AUTOCONFIG.N_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_0_1_LC_7_9_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_0_1_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_0_1_LC_7_9_2 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_RNO_0_1_LC_7_9_2  (
            .in0(N__6221),
            .in1(N__6116),
            .in2(_gnd_net_),
            .in3(N__5964),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.N_105_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_1_LC_7_9_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_1_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.PR_OUT_1_LC_7_9_3 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_1_LC_7_9_3  (
            .in0(N__5386),
            .in1(N__6220),
            .in2(N__5380),
            .in3(N__5493),
            .lcout(\U409_AUTOCONFIG.PR_OUTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.PR_OUT_1C_net ),
            .ce(N__6268),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_i_o4_0_LC_7_9_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_i_o4_0_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_i_o4_0_LC_7_9_4 .LUT_INIT=16'b0111001100110011;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_7_i_o4_0_LC_7_9_4  (
            .in0(N__6219),
            .in1(N__11852),
            .in2(N__6887),
            .in3(N__5963),
            .lcout(\U409_AUTOCONFIG.N_91 ),
            .ltout(\U409_AUTOCONFIG.N_91_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_7_9_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_7_9_5 .LUT_INIT=16'b0000110100001101;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_7_9_5  (
            .in0(N__6348),
            .in1(N__6850),
            .in2(N__5557),
            .in3(_gnd_net_),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.PR_OUT_1C_net ),
            .ce(N__6268),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_7_10_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_7_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_7_10_0 .LUT_INIT=16'b0000001000001010;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_7_10_0  (
            .in0(N__11853),
            .in1(N__5547),
            .in2(N__5629),
            .in3(N__5931),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net ),
            .ce(N__6280),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_7_10_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_7_10_1 .LUT_INIT=16'b0010000001100000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_7_10_1  (
            .in0(N__5548),
            .in1(N__6928),
            .in2(N__5960),
            .in3(N__5613),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.LIDE_OUT_7_i_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_7_10_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_7_10_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_7_10_2 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_1_LC_7_10_2  (
            .in0(N__11854),
            .in1(_gnd_net_),
            .in2(N__5539),
            .in3(_gnd_net_),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net ),
            .ce(N__6280),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI7DMP_1_LC_7_10_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI7DMP_1_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI7DMP_1_LC_7_10_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNI7DMP_1_LC_7_10_3  (
            .in0(N__7455),
            .in1(N__5536),
            .in2(_gnd_net_),
            .in3(N__5530),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_RNI7DMPZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_3_LC_7_10_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_3_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.PR_OUT_3_LC_7_10_4 .LUT_INIT=16'b0000001010101010;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_3_LC_7_10_4  (
            .in0(N__11855),
            .in1(N__5515),
            .in2(N__6939),
            .in3(N__5935),
            .lcout(\U409_AUTOCONFIG.PR_OUTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net ),
            .ce(N__6280),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_0_2_LC_7_10_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_0_2_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_0_2_LC_7_10_5 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_RNO_0_2_LC_7_10_5  (
            .in0(N__6217),
            .in1(N__6932),
            .in2(N__5961),
            .in3(N__5492),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.PR_OUT_cnst_i_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_2_LC_7_10_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_2_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.PR_OUT_2_LC_7_10_6 .LUT_INIT=16'b0000010100001111;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_2_LC_7_10_6  (
            .in0(N__5628),
            .in1(_gnd_net_),
            .in2(N__5791),
            .in3(N__6216),
            .lcout(\U409_AUTOCONFIG.PR_OUTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net ),
            .ce(N__6280),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNIOGLSO_LC_7_11_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNIOGLSO_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNIOGLSO_LC_7_11_0 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_RNIOGLSO_LC_7_11_0  (
            .in0(N__7099),
            .in1(N__6672),
            .in2(_gnd_net_),
            .in3(N__8421),
            .lcout(PORTSIZE_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_STATE_6_1_LC_7_11_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_STATE_6_1_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_STATE_6_1_LC_7_11_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_AUTOCONFIG.un1_STATE_6_1_LC_7_11_1  (
            .in0(N__5675),
            .in1(N__6212),
            .in2(N__5755),
            .in3(N__6051),
            .lcout(\U409_AUTOCONFIG.un1_STATE_6Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_0_3_LC_7_11_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_0_3_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_0_3_LC_7_11_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_0_3_LC_7_11_4  (
            .in0(N__7074),
            .in1(N__7003),
            .in2(N__5754),
            .in3(N__5674),
            .lcout(\U409_AUTOCONFIG.N_109 ),
            .ltout(\U409_AUTOCONFIG.N_109_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_1_LC_7_11_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_1_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_1_LC_7_11_5 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_1_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(N__6049),
            .in2(N__5632),
            .in3(N__6927),
            .lcout(\U409_AUTOCONFIG.N_117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_i_a2_0_0_LC_7_11_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_i_a2_0_0_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_i_a2_0_0_LC_7_11_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_7_i_a2_0_0_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(N__6211),
            .in2(_gnd_net_),
            .in3(N__6050),
            .lcout(\U409_AUTOCONFIG.N_113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_7_12_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_7_12_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_7_12_3  (
            .in0(N__5602),
            .in1(N__6142),
            .in2(N__6105),
            .in3(N__5939),
            .lcout(\U409_AUTOCONFIG.N_101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BREG_ENn_4_LC_8_6_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BREG_ENn_4_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BREG_ENn_4_LC_8_6_7 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BREG_ENn_4_LC_8_6_7  (
            .in0(N__7516),
            .in1(N__9744),
            .in2(_gnd_net_),
            .in3(N__6496),
            .lcout(\U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_0_LC_8_7_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_0_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_0_LC_8_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_0_LC_8_7_3  (
            .in0(N__10107),
            .in1(N__9913),
            .in2(N__10005),
            .in3(N__7798),
            .lcout(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0 ),
            .ltout(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_8_7_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_8_7_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_8_7_4  (
            .in0(N__8532),
            .in1(N__9729),
            .in2(N__5872),
            .in3(N__7734),
            .lcout(U409_ADDRESS_DECODE_un1_RTC_ENn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BREG_ENn_2_LC_8_7_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BREG_ENn_2_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BREG_ENn_2_LC_8_7_6 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BREG_ENn_2_LC_8_7_6  (
            .in0(N__7797),
            .in1(N__7733),
            .in2(N__6433),
            .in3(N__8101),
            .lcout(\U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_LC_8_7_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_LC_8_7_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_LC_8_7_7  (
            .in0(_gnd_net_),
            .in1(N__8867),
            .in2(_gnd_net_),
            .in3(N__8413),
            .lcout(un1_AUTOCONFIG_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_8_8_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_8_8_0 .LUT_INIT=16'b0000100000001010;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_8_8_0  (
            .in0(N__11848),
            .in1(N__6934),
            .in2(N__5887),
            .in3(N__5869),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net ),
            .ce(N__6278),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_8_8_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_8_8_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_3_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__11849),
            .in2(_gnd_net_),
            .in3(N__5886),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net ),
            .ce(N__6278),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIH4AI_LC_8_8_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIH4AI_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIH4AI_LC_8_8_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNIH4AI_LC_8_8_2  (
            .in0(N__6535),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7436),
            .lcout(\U409_AUTOCONFIG.D_OUT_sm0_0 ),
            .ltout(\U409_AUTOCONFIG.D_OUT_sm0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_RNI23A12_3_LC_8_8_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_RNI23A12_3_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_RNI23A12_3_LC_8_8_3 .LUT_INIT=16'b1111101011001010;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_RNI23A12_3_LC_8_8_3  (
            .in0(N__5803),
            .in1(N__5848),
            .in2(N__5839),
            .in3(N__7625),
            .lcout(D_OUT_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIBHMP_3_LC_8_8_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIBHMP_3_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIBHMP_3_LC_8_8_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNIBHMP_3_LC_8_8_4  (
            .in0(N__5815),
            .in1(N__5809),
            .in2(_gnd_net_),
            .in3(N__7438),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_RNIBHMPZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI5BMP_0_LC_8_8_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI5BMP_0_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI5BMP_0_LC_8_8_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNI5BMP_0_LC_8_8_5  (
            .in0(N__7437),
            .in1(N__5797),
            .in2(_gnd_net_),
            .in3(N__6286),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.LIDE_OUT_RNI5BMPZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_RNIPP912_0_LC_8_8_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_RNIPP912_0_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_RNIPP912_0_LC_8_8_6 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_RNIPP912_0_LC_8_8_6  (
            .in0(N__6391),
            .in1(N__7620),
            .in2(N__6385),
            .in3(N__6380),
            .lcout(D_OUT_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_0_LC_8_8_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_0_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_0_LC_8_8_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_0_LC_8_8_7  (
            .in0(N__7435),
            .in1(N__6534),
            .in2(N__6940),
            .in3(N__6955),
            .lcout(\U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_8_9_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_8_9_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_8_9_0 .LUT_INIT=16'b0101000100000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_2_LC_8_9_0  (
            .in0(N__6331),
            .in1(N__6349),
            .in2(N__6922),
            .in3(N__11850),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_2C_net ),
            .ce(N__6267),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_8_9_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_8_9_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_8_9_3  (
            .in0(N__6226),
            .in1(N__5978),
            .in2(N__6117),
            .in3(N__6894),
            .lcout(\U409_AUTOCONFIG.N_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_START_RNI04BC_LC_8_9_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_START_RNI04BC_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.AC_START_RNI04BC_LC_8_9_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U409_AUTOCONFIG.AC_START_RNI04BC_LC_8_9_4  (
            .in0(N__6325),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6418),
            .lcout(\U409_AUTOCONFIG.STATE4 ),
            .ltout(\U409_AUTOCONFIG.STATE4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNI10V92_1_LC_8_9_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNI10V92_1_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNI10V92_1_LC_8_9_5 .LUT_INIT=16'b0101010111010101;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNI10V92_1_LC_8_9_5  (
            .in0(N__11851),
            .in1(N__6412),
            .in2(N__6310),
            .in3(N__8905),
            .lcout(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_8_9_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_8_9_6 .LUT_INIT=16'b0000100100000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_8_9_6  (
            .in0(N__6106),
            .in1(N__6225),
            .in2(N__6921),
            .in3(N__5968),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.N_103_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_8_9_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_8_9_7 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_8_9_7  (
            .in0(N__6306),
            .in1(_gnd_net_),
            .in2(N__6289),
            .in3(N__11837),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_2C_net ),
            .ce(N__6267),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_0_a2_3_LC_8_10_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_0_a2_3_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_0_a2_3_LC_8_10_2 .LUT_INIT=16'b1001000000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_7_0_a2_3_LC_8_10_2  (
            .in0(N__6224),
            .in1(N__6084),
            .in2(N__6933),
            .in3(N__5950),
            .lcout(\U409_AUTOCONFIG.N_115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_START_LC_8_10_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_START_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.AC_START_LC_8_10_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U409_AUTOCONFIG.AC_START_LC_8_10_3  (
            .in0(N__7624),
            .in1(N__10394),
            .in2(_gnd_net_),
            .in3(N__8417),
            .lcout(\U409_AUTOCONFIG.AC_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11169),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNIJFAU_0_LC_8_10_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNIJFAU_0_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNIJFAU_0_LC_8_10_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNIJFAU_0_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(N__8856),
            .in2(_gnd_net_),
            .in3(N__8782),
            .lcout(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_8_11_2 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_8_11_2 .LUT_INIT=16'b0000001000010000;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_1_LC_8_11_2  (
            .in0(N__7311),
            .in1(N__7360),
            .in2(N__11573),
            .in3(N__7285),
            .lcout(),
            .ltout(\U409_CIA.CLK_CIA_r_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_LC_8_11_3 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_LC_8_11_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CLK_CIA_LC_8_11_3 .LUT_INIT=16'b1010101001101010;
    LogicCell40 \U409_CIA.CLK_CIA_LC_8_11_3  (
            .in0(N__11566),
            .in1(N__6466),
            .in2(N__6406),
            .in3(N__7338),
            .lcout(CLK_CIA_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12844),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_8_12_0 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_8_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(N__7251),
            .in2(N__7228),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_8_12_1 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_8_12_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_8_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_2_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(N__7359),
            .in2(_gnd_net_),
            .in3(N__6403),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .clk(N__12846),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_8_12_2 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_8_12_2 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_8_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_3_LC_8_12_2  (
            .in0(N__7260),
            .in1(N__7306),
            .in2(_gnd_net_),
            .in3(N__6400),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .clk(N__12846),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_8_12_3 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_8_12_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_8_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_4_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__7284),
            .in2(_gnd_net_),
            .in3(N__6397),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .clk(N__12846),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_8_12_4 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_8_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_5_LC_8_12_4  (
            .in0(N__7261),
            .in1(N__7336),
            .in2(_gnd_net_),
            .in3(N__6394),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .clk(N__12846),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_8_12_5 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_8_12_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_8_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_6_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(N__7174),
            .in2(_gnd_net_),
            .in3(N__6472),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ),
            .clk(N__12846),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_8_12_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_8_12_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_7_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(N__7191),
            .in2(_gnd_net_),
            .in3(N__6469),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12846),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_8_12_7 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_8_12_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_0_LC_8_12_7  (
            .in0(N__7252),
            .in1(N__7173),
            .in2(N__7192),
            .in3(N__7224),
            .lcout(\U409_CIA.CLK_CIA6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BREG_ENn_3_LC_9_6_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BREG_ENn_3_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BREG_ENn_3_LC_9_6_4 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BREG_ENn_3_LC_9_6_4  (
            .in0(N__10016),
            .in1(N__10108),
            .in2(N__7993),
            .in3(N__6487),
            .lcout(\U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_9_6_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_9_6_7 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_9_6_7  (
            .in0(N__8543),
            .in1(N__6460),
            .in2(N__9760),
            .in3(N__7723),
            .lcout(U409_ADDRESS_DECODE_un1_RTC_ENn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_1_LC_9_7_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_1_LC_9_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_1_LC_9_7_1 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_1_LC_9_7_1  (
            .in0(N__7874),
            .in1(N__7493),
            .in2(N__8137),
            .in3(N__7747),
            .lcout(LIDE_BASE_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_1C_net ),
            .ce(),
            .sr(N__11393));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_9_7_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_9_7_3 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_9_7_3  (
            .in0(N__7873),
            .in1(N__6429),
            .in2(N__6752),
            .in3(N__8014),
            .lcout(BRIDGE_BASE_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_1C_net ),
            .ce(),
            .sr(N__11393));
    defparam \U409_AUTOCONFIG.LIDE_BASE_2_LC_9_7_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_2_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_2_LC_9_7_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_2_LC_9_7_4  (
            .in0(N__7494),
            .in1(N__7875),
            .in2(N__7657),
            .in3(N__6744),
            .lcout(LIDE_BASE_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_1C_net ),
            .ce(),
            .sr(N__11393));
    defparam \U409_AUTOCONFIG.LIDE_BASE_5_LC_9_7_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_5_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_5_LC_9_7_5 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_5_LC_9_7_5  (
            .in0(N__7971),
            .in1(N__7876),
            .in2(N__8138),
            .in3(N__7549),
            .lcout(LIDE_BASE_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_1C_net ),
            .ce(),
            .sr(N__11393));
    defparam \U409_AUTOCONFIG.LIDE_BASE_6_LC_9_7_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_6_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_6_LC_9_7_6 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_6_LC_9_7_6  (
            .in0(N__7877),
            .in1(N__7972),
            .in2(N__7564),
            .in3(N__6745),
            .lcout(LIDE_BASE_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_1C_net ),
            .ce(),
            .sr(N__11393));
    defparam \U409_AUTOCONFIG.CONFIGURED_LC_9_7_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.CONFIGURED_LC_9_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.CONFIGURED_LC_9_7_7 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \U409_AUTOCONFIG.CONFIGURED_LC_9_7_7  (
            .in0(N__6544),
            .in1(N__6628),
            .in2(N__7450),
            .in3(N__7612),
            .lcout(CONFIGURED),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_1C_net ),
            .ce(),
            .sr(N__11393));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_9_8_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_9_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_9_8_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_9_8_0  (
            .in0(N__7865),
            .in1(N__6600),
            .in2(N__7953),
            .in3(N__8011),
            .lcout(BRIDGE_BASE_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_0C_net ),
            .ce(),
            .sr(N__11392));
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1_LC_9_8_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1_LC_9_8_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1_LC_9_8_1  (
            .in0(N__6923),
            .in1(N__7406),
            .in2(_gnd_net_),
            .in3(N__6953),
            .lcout(\U409_AUTOCONFIG.BRIDGE_CONF_RNID7FUZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BREG_ENn_1_LC_9_8_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BREG_ENn_1_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BREG_ENn_1_LC_9_8_2 .LUT_INIT=16'b1000000000001000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BREG_ENn_1_LC_9_8_2  (
            .in0(N__7613),
            .in1(N__9395),
            .in2(N__9301),
            .in3(N__6601),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BREG_ENn_i_LC_9_8_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BREG_ENn_i_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BREG_ENn_i_LC_9_8_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BREG_ENn_i_LC_9_8_3  (
            .in0(N__6592),
            .in1(N__6583),
            .in2(N__6574),
            .in3(N__6571),
            .lcout(U409_ADDRESS_DECODE_un1_BREG_ENn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_1_LC_9_8_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_1_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_1_LC_9_8_7 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_1_LC_9_8_7  (
            .in0(N__7407),
            .in1(N__6543),
            .in2(N__6938),
            .in3(N__6954),
            .lcout(\U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BREG_ENn_0_LC_9_9_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BREG_ENn_0_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BREG_ENn_0_LC_9_9_2 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BREG_ENn_0_LC_9_9_2  (
            .in0(N__9899),
            .in1(N__10209),
            .in2(N__6688),
            .in3(N__7084),
            .lcout(\U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_4_LC_9_9_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_4_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_4_LC_9_9_3 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_4_LC_9_9_3  (
            .in0(N__7888),
            .in1(N__6483),
            .in2(N__7954),
            .in3(N__7529),
            .lcout(BRIDGE_BASE_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_4C_net ),
            .ce(),
            .sr(N__11388));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_7_LC_9_9_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_7_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_7_LC_9_9_4 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_7_LC_9_9_4  (
            .in0(N__7530),
            .in1(N__7890),
            .in2(N__8061),
            .in3(N__7083),
            .lcout(BRIDGE_BASE_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_4C_net ),
            .ce(),
            .sr(N__11388));
    defparam \U409_AUTOCONFIG.STATE_RNIU6QK1_0_LC_9_9_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNIU6QK1_0_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNIU6QK1_0_LC_9_9_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNIU6QK1_0_LC_9_9_5  (
            .in0(N__7075),
            .in1(N__7018),
            .in2(N__6970),
            .in3(N__8920),
            .lcout(\U409_AUTOCONFIG.un1_STATE_6_0 ),
            .ltout(\U409_AUTOCONFIG.un1_STATE_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1_0_LC_9_9_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1_0_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1_0_LC_9_9_6 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1_0_LC_9_9_6  (
            .in0(N__6864),
            .in1(_gnd_net_),
            .in2(N__6757),
            .in3(N__7427),
            .lcout(\U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1Z0Z_0 ),
            .ltout(\U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_6_LC_9_9_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_6_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_6_LC_9_9_7 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_6_LC_9_9_7  (
            .in0(N__7889),
            .in1(N__6753),
            .in2(N__6691),
            .in3(N__6684),
            .lcout(BRIDGE_BASE_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_4C_net ),
            .ce(),
            .sr(N__11388));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_9_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_9_10_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_9_10_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__8205),
            .in2(_gnd_net_),
            .in3(N__8191),
            .lcout(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__8673));
    defparam \U409_CIA.VMA_RNO_0_LC_9_11_3 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_0_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_0_LC_9_11_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_CIA.VMA_RNO_0_LC_9_11_3  (
            .in0(N__7366),
            .in1(N__7337),
            .in2(N__7312),
            .in3(N__7159),
            .lcout(),
            .ltout(\U409_CIA.VMA_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_LC_9_11_4 .C_ON=1'b0;
    defparam \U409_CIA.VMA_LC_9_11_4 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.VMA_LC_9_11_4 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \U409_CIA.VMA_LC_9_11_4  (
            .in0(N__6676),
            .in1(N__10904),
            .in2(N__6658),
            .in3(N__7225),
            .lcout(\U409_CIA.VMAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12843),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_0_0_0_LC_9_11_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_0_0_0_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_0_0_0_LC_9_11_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_0_a3_0_0_0_LC_9_11_6  (
            .in0(N__9895),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10090),
            .lcout(\U409_ADDRESS_DECODE.un1_RTC_ENn_2 ),
            .ltout(\U409_ADDRESS_DECODE.un1_RTC_ENn_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_9_11_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_9_11_7 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_9_11_7  (
            .in0(N__8496),
            .in1(N__8544),
            .in2(N__6655),
            .in3(N__9708),
            .lcout(U409_ADDRESS_DECODE_un1_REGSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_1_LC_9_12_1 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_1_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_1_LC_9_12_1 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \U409_CIA.VMA_RNO_1_LC_9_12_1  (
            .in0(N__7248),
            .in1(N__7282),
            .in2(N__7226),
            .in3(N__7358),
            .lcout(\U409_CIA.un1_CIA_CLK_COUNT_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIGOMD1_2_LC_9_12_2 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIGOMD1_2_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIGOMD1_2_LC_9_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIGOMD1_2_LC_9_12_2  (
            .in0(N__7357),
            .in1(N__7214),
            .in2(N__7339),
            .in3(N__7247),
            .lcout(),
            .ltout(\U409_CIA.CIA_CLK_COUNT11_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNICTDR2_3_LC_9_12_3 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNICTDR2_3_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNICTDR2_3_LC_9_12_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNICTDR2_3_LC_9_12_3  (
            .in0(N__7307),
            .in1(N__7283),
            .in2(N__7264),
            .in3(N__7158),
            .lcout(\U409_CIA.CIA_CLK_COUNT11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_9_12_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_9_12_4 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_9_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_0_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7249),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12845),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_9_12_5 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_9_12_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_9_12_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_1_LC_9_12_5  (
            .in0(N__7250),
            .in1(_gnd_net_),
            .in2(N__7227),
            .in3(_gnd_net_),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12845),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_9_12_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_9_12_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(N__7187),
            .in2(_gnd_net_),
            .in3(N__7172),
            .lcout(\U409_CIA.CLK_CIA6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.m20_LC_10_6_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.m20_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.m20_LC_10_6_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_ADDRESS_DECODE.m20_LC_10_6_5  (
            .in0(N__9398),
            .in1(N__9758),
            .in2(N__9100),
            .in3(N__10017),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.N_77_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.N_22_0_i_LC_10_6_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.N_22_0_i_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.N_22_0_i_LC_10_6_6 .LUT_INIT=16'b1100111111001111;
    LogicCell40 \U409_ADDRESS_DECODE.N_22_0_i_LC_10_6_6  (
            .in0(_gnd_net_),
            .in1(N__10111),
            .in2(N__7147),
            .in3(_gnd_net_),
            .lcout(N_22_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNIO8F0F_LC_10_7_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNIO8F0F_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNIO8F0F_LC_10_7_0 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_RNIO8F0F_LC_10_7_0  (
            .in0(N__7116),
            .in1(N__8357),
            .in2(N__8743),
            .in3(N__8343),
            .lcout(\U409_ADDRESS_DECODE.PORTSIZE_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_0_LC_10_7_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_0_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_0_LC_10_7_2 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_0_LC_10_7_2  (
            .in0(N__7813),
            .in1(N__7746),
            .in2(N__7732),
            .in3(N__7653),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_LC_10_7_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_LC_10_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_LC_10_7_3  (
            .in0(N__7570),
            .in1(N__7537),
            .in2(N__7642),
            .in3(N__8428),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACEZ0 ),
            .ltout(\U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_LC_10_7_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_LC_10_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_LC_10_7_4 .LUT_INIT=16'b1010101000100000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_LC_10_7_4  (
            .in0(N__11815),
            .in1(N__8866),
            .in2(N__7639),
            .in3(N__8342),
            .lcout(\U409_ADDRESS_DECODE.ATA_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11175),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_10_7_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_10_7_6 .LUT_INIT=16'b1000001000000000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_10_7_6  (
            .in0(N__9396),
            .in1(N__10214),
            .in2(N__8080),
            .in3(N__7608),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_10_7_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_10_7_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_10_7_7 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_10_7_7  (
            .in0(N__9914),
            .in1(N__7560),
            .in2(N__9754),
            .in3(N__7548),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_5_LC_10_8_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_5_LC_10_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_5_LC_10_8_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_5_LC_10_8_0  (
            .in0(N__8148),
            .in1(N__7909),
            .in2(N__7512),
            .in3(N__7531),
            .lcout(BRIDGE_BASE_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_5C_net ),
            .ce(),
            .sr(N__11389));
    defparam \U409_AUTOCONFIG.LIDE_BASE_3_LC_10_8_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_3_LC_10_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_3_LC_10_8_1 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_3_LC_10_8_1  (
            .in0(N__7910),
            .in1(N__7495),
            .in2(N__8443),
            .in3(N__8047),
            .lcout(LIDE_BASE_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_5C_net ),
            .ce(),
            .sr(N__11389));
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_LC_10_8_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_LC_10_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_LC_10_8_2 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_CONF_LC_10_8_2  (
            .in0(N__7477),
            .in1(N__7428),
            .in2(_gnd_net_),
            .in3(N__8919),
            .lcout(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_5C_net ),
            .ce(),
            .sr(N__11389));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_10_8_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_10_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_10_8_4 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_10_8_4  (
            .in0(N__8147),
            .in1(N__8012),
            .in2(N__8097),
            .in3(N__7907),
            .lcout(BRIDGE_BASE_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_5C_net ),
            .ce(),
            .sr(N__11389));
    defparam \U409_AUTOCONFIG.LIDE_BASE_7_LC_10_8_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_7_LC_10_8_5 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_7_LC_10_8_5 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_7_LC_10_8_5  (
            .in0(N__7970),
            .in1(N__8048),
            .in2(N__7918),
            .in3(N__8076),
            .lcout(LIDE_BASE_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_5C_net ),
            .ce(),
            .sr(N__11389));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_10_8_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_10_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_10_8_6 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_10_8_6  (
            .in0(N__8046),
            .in1(N__8013),
            .in2(N__7989),
            .in3(N__7908),
            .lcout(BRIDGE_BASE_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_5C_net ),
            .ce(),
            .sr(N__11389));
    defparam \U409_AUTOCONFIG.LIDE_BASE_4_LC_10_8_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_4_LC_10_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_4_LC_10_8_7 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_4_LC_10_8_7  (
            .in0(N__7969),
            .in1(N__7952),
            .in2(N__7917),
            .in3(N__8455),
            .lcout(LIDE_BASE_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_5C_net ),
            .ce(),
            .sr(N__11389));
    defparam \U409_ADDRESS_DECODE.m33_LC_10_9_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.m33_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.m33_LC_10_9_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.m33_LC_10_9_0  (
            .in0(N__8242),
            .in1(N__8565),
            .in2(N__8311),
            .in3(N__7819),
            .lcout(N_71_mux),
            .ltout(N_71_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.m38_LC_10_9_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.m38_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.m38_LC_10_9_1 .LUT_INIT=16'b0001110100111111;
    LogicCell40 \U409_ADDRESS_DECODE.m38_LC_10_9_1  (
            .in0(N__11498),
            .in1(N__8976),
            .in2(N__7825),
            .in3(N__8942),
            .lcout(N_23),
            .ltout(N_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_9_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_9_2 .LUT_INIT=16'b0011000011000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(N__8223),
            .in2(N__7822),
            .in3(N__8567),
            .lcout(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__8674));
    defparam \U409_ADDRESS_DECODE.m33_3_LC_10_9_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.m33_3_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.m33_3_LC_10_9_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.m33_3_LC_10_9_3  (
            .in0(N__8221),
            .in1(N__8187),
            .in2(N__8595),
            .in3(N__8269),
            .lcout(\U409_ADDRESS_DECODE.m33Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.m27_3_LC_10_9_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.m27_3_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.m27_3_LC_10_9_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.m27_3_LC_10_9_4  (
            .in0(N__8188),
            .in1(N__8222),
            .in2(N__8275),
            .in3(N__8586),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.m27Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.m27_LC_10_9_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.m27_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.m27_LC_10_9_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_ADDRESS_DECODE.m27_LC_10_9_5  (
            .in0(N__8566),
            .in1(N__8308),
            .in2(N__8287),
            .in3(N__8243),
            .lcout(N_70_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_9_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_9_6 .LUT_INIT=16'b0111000010000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_9_6  (
            .in0(N__8284),
            .in1(N__8979),
            .in2(N__8623),
            .in3(N__8309),
            .lcout(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__8674));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_7 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_7  (
            .in0(N__8978),
            .in1(N__8283),
            .in2(_gnd_net_),
            .in3(N__8619),
            .lcout(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__8674));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_10_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_10_0  (
            .in0(N__8244),
            .in1(N__8254),
            .in2(N__8206),
            .in3(N__8190),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_10_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_10_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_10_1 .LUT_INIT=16'b0110101000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_10_1  (
            .in0(N__8274),
            .in1(N__8160),
            .in2(N__8596),
            .in3(N__8621),
            .lcout(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net ),
            .ce(),
            .sr(N__8656));
    defparam \U409_ADDRESS_DECODE.m33_1_LC_10_10_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.m33_1_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.m33_1_LC_10_10_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_ADDRESS_DECODE.m33_1_LC_10_10_2  (
            .in0(_gnd_net_),
            .in1(N__8590),
            .in2(_gnd_net_),
            .in3(N__8273),
            .lcout(U409_ADDRESS_DECODE_m33_1),
            .ltout(U409_ADDRESS_DECODE_m33_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_10_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_10_3 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_10_3 .LUT_INIT=16'b0110101000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_10_3  (
            .in0(N__8245),
            .in1(N__8161),
            .in2(N__8248),
            .in3(N__8622),
            .lcout(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net ),
            .ce(),
            .sr(N__8656));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI7S9R_1_LC_10_10_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI7S9R_1_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI7S9R_1_LC_10_10_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI7S9R_1_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(N__8568),
            .in2(_gnd_net_),
            .in3(N__8224),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c2 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_10_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_10_10_5 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(N__8189),
            .in2(N__8164),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_10_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_10_6 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_10_6  (
            .in0(N__8620),
            .in1(_gnd_net_),
            .in2(N__8599),
            .in3(N__8591),
            .lcout(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net ),
            .ce(),
            .sr(N__8656));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_7 .LUT_INIT=16'b0111011001010101;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_7  (
            .in0(N__8569),
            .in1(N__8980),
            .in2(N__11497),
            .in3(N__8944),
            .lcout(U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net ),
            .ce(),
            .sr(N__8656));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER16_LC_10_11_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER16_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER16_LC_10_11_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER16_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(N__10395),
            .in2(_gnd_net_),
            .in3(N__11202),
            .lcout(N_52_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_10_11_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_10_11_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_10_11_2  (
            .in0(N__10245),
            .in1(N__8548),
            .in2(N__8503),
            .in3(N__9724),
            .lcout(U409_ADDRESS_DECODE_un1_REGSPACEn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_1_0_LC_11_7_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_1_0_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_1_0_LC_11_7_4 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_1_0_LC_11_7_4  (
            .in0(N__10110),
            .in1(N__8454),
            .in2(N__10009),
            .in3(N__8439),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACE_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.LV_SPACE_LC_11_7_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.LV_SPACE_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.LV_SPACE_LC_11_7_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.LV_SPACE_LC_11_7_5  (
            .in0(N__8742),
            .in1(N__8688),
            .in2(N__8362),
            .in3(N__8422),
            .lcout(BUFENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_LC_11_7_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_LC_11_7_6 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(N__8358),
            .in2(_gnd_net_),
            .in3(N__8344),
            .lcout(U409_ADDRESS_DECODE_un1_ATA_ENn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_LC_11_8_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_LC_11_8_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_LC_11_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8310),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_EN_nerC_net ),
            .ce(N__8926),
            .sr(N__8666));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_11_9_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_11_9_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_11_9_0  (
            .in0(N__9018),
            .in1(N__9399),
            .in2(N__10219),
            .in3(N__9796),
            .lcout(U409_ADDRESS_DECODE_un1_RAMSPACEn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_1_LC_11_9_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_1_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.STATE_1_LC_11_9_1 .LUT_INIT=16'b0001000011000000;
    LogicCell40 \U409_AUTOCONFIG.STATE_1_LC_11_9_1  (
            .in0(N__8837),
            .in1(N__8895),
            .in2(N__11836),
            .in3(N__8770),
            .lcout(\U409_AUTOCONFIG.STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.STATE_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_0_LC_11_9_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_0_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.STATE_0_LC_11_9_2 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \U409_AUTOCONFIG.STATE_0_LC_11_9_2  (
            .in0(N__8769),
            .in1(N__11788),
            .in2(N__8903),
            .in3(N__8989),
            .lcout(\U409_AUTOCONFIG.STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.STATE_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_sbtinv_LC_11_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_sbtinv_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_sbtinv_LC_11_9_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_sbtinv_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__8977),
            .in2(N__8953),
            .in3(N__8943),
            .lcout(\U409_TRANSFER_ACK.N_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNIF4QU_0_LC_11_9_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNIF4QU_0_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNIF4QU_0_LC_11_9_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNIF4QU_0_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__8891),
            .in2(_gnd_net_),
            .in3(N__8768),
            .lcout(\U409_AUTOCONFIG.STATE_d_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_TACK_LC_11_10_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_TACK_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.AC_TACK_LC_11_10_0 .LUT_INIT=16'b1111111010001000;
    LogicCell40 \U409_AUTOCONFIG.AC_TACK_LC_11_10_0  (
            .in0(N__9522),
            .in1(N__8902),
            .in2(N__8869),
            .in3(N__8777),
            .lcout(AC_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.AC_TACKC_net ),
            .ce(),
            .sr(N__11383));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_11_11_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_11_11_4 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_11_11_4  (
            .in0(N__8726),
            .in1(N__8710),
            .in2(N__8692),
            .in3(N__11795),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_1_LC_11_12_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_1_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_1_LC_11_12_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_0_a3_1_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(N__9912),
            .in2(_gnd_net_),
            .in3(N__9723),
            .lcout(\U409_ADDRESS_DECODE.N_60_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_3.C_ON=1'b0;
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_3.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11206),
            .lcout(GB_BUFFER_CLK40_IN_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CS0_LC_12_3_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CS0_LC_12_3_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CS0_LC_12_3_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_ADDRESS_DECODE.CS0_LC_12_3_1  (
            .in0(N__9296),
            .in1(N__9237),
            .in2(N__9215),
            .in3(N__9150),
            .lcout(\U409_ADDRESS_DECODE.CSZ0Z0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CS1_LC_12_3_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CS1_LC_12_3_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CS1_LC_12_3_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_ADDRESS_DECODE.CS1_LC_12_3_5  (
            .in0(N__9297),
            .in1(N__9238),
            .in2(N__9216),
            .in3(N__9151),
            .lcout(\U409_ADDRESS_DECODE.CSZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_12_5_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_12_5_1 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_12_5_1  (
            .in0(N__9217),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9160),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS1n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNI692L_0_LC_12_5_5 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNI692L_0_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNI692L_0_LC_12_5_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_CIA.VMA_RNI692L_0_LC_12_5_5  (
            .in0(N__11731),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10924),
            .lcout(CIA_ENABLE),
            .ltout(CIA_ENABLE_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_12_5_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_12_5_6 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_12_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9154),
            .in3(N__9141),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS0n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.N_77_mux_i_LC_12_6_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.N_77_mux_i_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.N_77_mux_i_LC_12_6_0 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \U409_ADDRESS_DECODE.N_77_mux_i_LC_12_6_0  (
            .in0(N__9403),
            .in1(N__9096),
            .in2(N__10010),
            .in3(N__9759),
            .lcout(N_77_mux_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_12_7_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_12_7_3 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_12_7_3  (
            .in0(N__9397),
            .in1(N__9785),
            .in2(N__9025),
            .in3(N__10190),
            .lcout(U409_ADDRESS_DECODE_un1_RAMSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_12_8_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_12_8_2 .LUT_INIT=16'b0010000000110000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_12_8_2  (
            .in0(N__9450),
            .in1(N__9432),
            .in2(N__11775),
            .in3(N__9414),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_12_8_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_12_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_12_8_3 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_12_8_3  (
            .in0(N__9431),
            .in1(N__11738),
            .in2(_gnd_net_),
            .in3(N__9449),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_RNIKDE9_LC_12_8_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_RNIKDE9_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_RNIKDE9_LC_12_8_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_RNIKDE9_LC_12_8_4  (
            .in0(_gnd_net_),
            .in1(N__9529),
            .in2(_gnd_net_),
            .in3(N__10332),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIFT8M_LC_12_8_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIFT8M_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIFT8M_LC_12_8_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNIFT8M_LC_12_8_5  (
            .in0(N__9523),
            .in1(N__10939),
            .in2(N__9508),
            .in3(N__10314),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER6 ),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_12_8_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_12_8_6 .LUT_INIT=16'b0000000111011101;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_12_8_6  (
            .in0(N__9448),
            .in1(N__9430),
            .in2(N__9505),
            .in3(N__9469),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_12_8_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_12_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_12_8_7 .LUT_INIT=16'b0000111110101010;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_LC_12_8_7  (
            .in0(N__9470),
            .in1(_gnd_net_),
            .in2(N__9502),
            .in3(N__11739),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_9_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_9_0 .LUT_INIT=16'b0000000010011001;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_9_0  (
            .in0(N__10888),
            .in1(N__10806),
            .in2(_gnd_net_),
            .in3(N__11463),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__11382));
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_12_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_12_9_7 .LUT_INIT=16'b0111000001110001;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_LC_12_9_7  (
            .in0(N__9451),
            .in1(N__9433),
            .in2(N__9589),
            .in3(N__9415),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__11382));
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a2_LC_12_10_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a2_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a2_LC_12_10_0 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_0_a2_LC_12_10_0  (
            .in0(N__10024),
            .in1(N__9388),
            .in2(N__10234),
            .in3(N__9622),
            .lcout(ROMEN),
            .ltout(ROMEN_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIRHPR5_0_LC_12_10_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIRHPR5_0_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIRHPR5_0_LC_12_10_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIRHPR5_0_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9307),
            .in3(N__11434),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0 ),
            .ltout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_10_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_10_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_10_2  (
            .in0(N__10755),
            .in1(N__10805),
            .in2(N__9304),
            .in3(N__10858),
            .lcout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_0_LC_12_10_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_0_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_0_LC_12_10_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_0_a3_0_LC_12_10_3  (
            .in0(N__9740),
            .in1(N__10252),
            .in2(N__10218),
            .in3(N__10011),
            .lcout(\U409_ADDRESS_DECODE.N_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIV1RD_3_LC_12_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIV1RD_3_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIV1RD_3_LC_12_10_5 .LUT_INIT=16'b0100010010111011;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIV1RD_3_LC_12_10_5  (
            .in0(N__10647),
            .in1(N__10715),
            .in2(_gnd_net_),
            .in3(N__10754),
            .lcout(\U409_TRANSFER_ACK.N_42_i ),
            .ltout(\U409_TRANSFER_ACK.N_42_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_2_LC_12_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_2_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_2_LC_12_10_6 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_2_LC_12_10_6  (
            .in0(N__11435),
            .in1(N__10648),
            .in2(N__10222),
            .in3(N__10707),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER22_NE_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_1_0_LC_12_10_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_1_0_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_1_0_LC_12_10_7 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_0_a3_1_0_LC_12_10_7  (
            .in0(N__10213),
            .in1(N__10109),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_2_LC_12_11_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_2_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_2_LC_12_11_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_0_a3_2_LC_12_11_5  (
            .in0(N__10012),
            .in1(N__9916),
            .in2(N__9795),
            .in3(N__9728),
            .lcout(\U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_RNIPUKQ5_LC_12_13_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_RNIPUKQ5_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_EN_RNIPUKQ5_LC_12_13_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_RNIPUKQ5_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__9616),
            .in2(_gnd_net_),
            .in3(N__9590),
            .lcout(TCIn_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_2.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_2.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11796),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_13_8_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_13_8_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_13_8_1  (
            .in0(N__10425),
            .in1(N__11203),
            .in2(N__10407),
            .in3(N__10348),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .ce(),
            .sr(N__11386));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_13_8_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_13_8_5 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_13_8_5  (
            .in0(N__10426),
            .in1(_gnd_net_),
            .in2(N__10408),
            .in3(N__11842),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_13_8_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_13_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_13_8_6 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_13_8_6  (
            .in0(N__11204),
            .in1(N__10347),
            .in2(N__10336),
            .in3(N__10333),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .ce(),
            .sr(N__11386));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_13_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_13_9_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_13_9_4 .LUT_INIT=16'b1111111101001100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_LC_13_9_4  (
            .in0(N__10321),
            .in1(N__10315),
            .in2(N__10726),
            .in3(N__10258),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .ce(),
            .sr(N__11385));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_13_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_13_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_13_9_5 .LUT_INIT=16'b0011000100000010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_13_9_5  (
            .in0(N__10807),
            .in1(N__11459),
            .in2(N__10887),
            .in3(N__10759),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .ce(),
            .sr(N__11385));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_13_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_13_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_13_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_13_9_6  (
            .in0(N__11458),
            .in1(N__10859),
            .in2(_gnd_net_),
            .in3(N__11440),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .ce(),
            .sr(N__11385));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI87LI_2_LC_13_10_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI87LI_2_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI87LI_2_LC_13_10_1 .LUT_INIT=16'b1100010000000010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI87LI_2_LC_13_10_1  (
            .in0(N__10646),
            .in1(N__10795),
            .in2(N__10717),
            .in3(N__10848),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_NE_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIGEA51_3_LC_13_10_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIGEA51_3_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIGEA51_3_LC_13_10_2 .LUT_INIT=16'b1000000000010000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIGEA51_3_LC_13_10_2  (
            .in0(N__10602),
            .in1(N__11436),
            .in2(N__10303),
            .in3(N__10756),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ),
            .ltout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_LC_13_10_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_13_10_3 .SEQ_MODE=4'b1001;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_13_10_3 .LUT_INIT=16'b1111010011111100;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_LC_13_10_3  (
            .in0(N__11505),
            .in1(N__10275),
            .in2(N__10300),
            .in3(N__10297),
            .lcout(ROMENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROMENnC_net ),
            .ce(),
            .sr(N__11384));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_13_10_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_13_10_7 .LUT_INIT=16'b0100100000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_13_10_7  (
            .in0(N__10861),
            .in1(N__10867),
            .in2(N__10808),
            .in3(N__10264),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER21_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.m43_LC_13_14_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.m43_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.m43_LC_13_14_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.m43_LC_13_14_4  (
            .in0(N__10489),
            .in1(N__10510),
            .in2(_gnd_net_),
            .in3(N__10534),
            .lcout(PCIAT_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.m45_LC_13_15_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.m45_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.m45_LC_13_15_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_ADDRESS_DECODE.m45_LC_13_15_3  (
            .in0(N__10533),
            .in1(N__10509),
            .in2(_gnd_net_),
            .in3(N__10482),
            .lcout(PCIAT_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_6_0 .C_ON=1'b1;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_6_0  (
            .in0(_gnd_net_),
            .in1(N__11315),
            .in2(N__10963),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_6_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_2_LC_14_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_2_LC_14_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_2_LC_14_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_2_LC_14_6_1  (
            .in0(_gnd_net_),
            .in1(N__11334),
            .in2(_gnd_net_),
            .in3(N__10444),
            .lcout(\U409_TICK.COUNTER60Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .clk(N__12598),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_3_LC_14_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_3_LC_14_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_3_LC_14_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_3_LC_14_6_2  (
            .in0(_gnd_net_),
            .in1(N__11265),
            .in2(_gnd_net_),
            .in3(N__10441),
            .lcout(\U409_TICK.COUNTER60Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .clk(N__12598),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_14_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_14_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_4_LC_14_6_3  (
            .in0(_gnd_net_),
            .in1(N__11067),
            .in2(_gnd_net_),
            .in3(N__10438),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_5_LC_14_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_5_LC_14_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_5_LC_14_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_5_LC_14_6_4  (
            .in0(_gnd_net_),
            .in1(N__11085),
            .in2(_gnd_net_),
            .in3(N__10435),
            .lcout(\U409_TICK.COUNTER60Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .clk(N__12598),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_14_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_14_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_6_LC_14_6_5  (
            .in0(_gnd_net_),
            .in1(N__11016),
            .in2(_gnd_net_),
            .in3(N__10432),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_7_LC_14_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_7_LC_14_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_7_LC_14_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_7_LC_14_6_6  (
            .in0(_gnd_net_),
            .in1(N__10977),
            .in2(_gnd_net_),
            .in3(N__10429),
            .lcout(\U409_TICK.COUNTER60Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .clk(N__12598),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_14_6_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_14_6_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_14_6_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_8_LC_14_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11044),
            .in3(N__10582),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_14_7_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_14_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_9_LC_14_7_0  (
            .in0(_gnd_net_),
            .in1(N__11055),
            .in2(_gnd_net_),
            .in3(N__10579),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_14_7_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_10_LC_14_7_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_10_LC_14_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_10_LC_14_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_10_LC_14_7_1  (
            .in0(_gnd_net_),
            .in1(N__10992),
            .in2(_gnd_net_),
            .in3(N__10576),
            .lcout(\U409_TICK.COUNTER60Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .clk(N__12599),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_11_LC_14_7_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_11_LC_14_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_11_LC_14_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_11_LC_14_7_2  (
            .in0(_gnd_net_),
            .in1(N__11280),
            .in2(_gnd_net_),
            .in3(N__10573),
            .lcout(\U409_TICK.COUNTER60Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .clk(N__12599),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_12_LC_14_7_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_12_LC_14_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_12_LC_14_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_12_LC_14_7_3  (
            .in0(_gnd_net_),
            .in1(N__11346),
            .in2(_gnd_net_),
            .in3(N__10570),
            .lcout(\U409_TICK.COUNTER60Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .clk(N__12599),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_13_LC_14_7_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_13_LC_14_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_13_LC_14_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_13_LC_14_7_4  (
            .in0(_gnd_net_),
            .in1(N__11004),
            .in2(_gnd_net_),
            .in3(N__10567),
            .lcout(\U409_TICK.COUNTER60Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .clk(N__12599),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_14_7_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_14_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_14_LC_14_7_5  (
            .in0(_gnd_net_),
            .in1(N__11244),
            .in2(_gnd_net_),
            .in3(N__10564),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_14_7_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_14_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_14_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_15_LC_14_7_6  (
            .in0(_gnd_net_),
            .in1(N__11220),
            .in2(_gnd_net_),
            .in3(N__10561),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_16_LC_14_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_16_LC_14_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_16_LC_14_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER60_16_LC_14_7_7  (
            .in0(_gnd_net_),
            .in1(N__11299),
            .in2(_gnd_net_),
            .in3(N__10558),
            .lcout(\U409_TICK.COUNTER60Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12599),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_14_8_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_14_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_14_8_0 .LUT_INIT=16'b0100111001001100;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_LC_14_8_0  (
            .in0(N__11627),
            .in1(N__10938),
            .in2(N__11650),
            .in3(N__11116),
            .lcout(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__11390));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_14_8_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_14_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_14_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_14_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11911),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__11390));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_14_8_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_14_8_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_14_8_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_14_8_5  (
            .in0(N__11838),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10923),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__11390));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_14_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_14_9_1 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_14_9_1  (
            .in0(N__11430),
            .in1(N__10812),
            .in2(N__10860),
            .in3(N__10758),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_0_LC_14_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_0_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_0_LC_14_9_6 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_0_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(N__10851),
            .in2(_gnd_net_),
            .in3(N__11429),
            .lcout(\U409_TRANSFER_ACK.N_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_3_LC_14_10_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_3_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_3_LC_14_10_2 .LUT_INIT=16'b0100001010000100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_3_LC_14_10_2  (
            .in0(N__10637),
            .in1(N__10849),
            .in2(N__10716),
            .in3(N__11420),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER21_NE_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_1_LC_14_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_1_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_1_LC_14_10_5 .LUT_INIT=16'b0100000110000010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_1_LC_14_10_5  (
            .in0(N__10850),
            .in1(N__10813),
            .in2(N__10603),
            .in3(N__10757),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER22_NE_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER21_0_i_0_x3_0_0_LC_14_11_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER21_0_i_0_x3_0_0_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER21_0_i_0_x3_0_0_LC_14_11_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER21_0_i_0_x3_0_0_LC_14_11_1  (
            .in0(_gnd_net_),
            .in1(N__10708),
            .in2(_gnd_net_),
            .in3(N__10628),
            .lcout(\U409_TRANSFER_ACK.N_31_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_9_LC_15_6_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_9_LC_15_6_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_9_LC_15_6_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_9_LC_15_6_0  (
            .in0(N__12049),
            .in1(N__12122),
            .in2(N__12090),
            .in3(N__10588),
            .lcout(\U409_TICK.COUNTER60Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12600),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_8_LC_15_6_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_8_LC_15_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_8_LC_15_6_1 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_8_LC_15_6_1  (
            .in0(N__12121),
            .in1(N__12051),
            .in2(N__11095),
            .in3(N__12086),
            .lcout(\U409_TICK.COUNTER60Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12600),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_1_LC_15_6_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_1_LC_15_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_1_LC_15_6_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER60_1_LC_15_6_3  (
            .in0(N__10961),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11319),
            .lcout(\U409_TICK.COUNTER60Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12600),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_15_6_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_15_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_15_6_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U409_TICK.COUNTER60_RNIHJU51_4_LC_15_6_4  (
            .in0(N__11086),
            .in1(N__10960),
            .in2(_gnd_net_),
            .in3(N__11068),
            .lcout(\U409_TICK.TICK603_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_4_LC_15_6_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_4_LC_15_6_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_4_LC_15_6_5 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \U409_TICK.COUNTER60_4_LC_15_6_5  (
            .in0(N__11074),
            .in1(N__12082),
            .in2(N__12124),
            .in3(N__12052),
            .lcout(\U409_TICK.COUNTER60Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12600),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_15_6_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_15_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_15_6_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNICDC71_14_LC_15_6_6  (
            .in0(N__11056),
            .in1(N__11043),
            .in2(N__11020),
            .in3(N__11245),
            .lcout(\U409_TICK.TICK603_9 ),
            .ltout(\U409_TICK.TICK603_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_6_LC_15_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_6_LC_15_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_6_LC_15_6_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_6_LC_15_6_7  (
            .in0(N__12120),
            .in1(N__12050),
            .in2(N__11029),
            .in3(N__11026),
            .lcout(\U409_TICK.COUNTER60Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12600),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_15_7_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_15_7_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_TICK.COUNTER60_RNI2USG_10_LC_15_7_0  (
            .in0(N__11005),
            .in1(N__10993),
            .in2(N__10981),
            .in3(N__11221),
            .lcout(\U409_TICK.TICK603_10 ),
            .ltout(\U409_TICK.TICK603_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_0_LC_15_7_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_0_LC_15_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_0_LC_15_7_1 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \U409_TICK.COUNTER60_0_LC_15_7_1  (
            .in0(N__12079),
            .in1(N__12053),
            .in2(N__10966),
            .in3(N__10962),
            .lcout(\U409_TICK.COUNTER60Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12603),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_15_7_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_15_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_15_7_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER60_RNIDB4S_16_LC_15_7_2  (
            .in0(N__11347),
            .in1(N__11335),
            .in2(N__11323),
            .in3(N__11298),
            .lcout(),
            .ltout(\U409_TICK.TICK603_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_15_7_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_15_7_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_15_7_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER60_RNI335G2_11_LC_15_7_3  (
            .in0(N__11287),
            .in1(N__11281),
            .in2(N__11269),
            .in3(N__11266),
            .lcout(\U409_TICK.TICK603_14 ),
            .ltout(\U409_TICK.TICK603_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_14_LC_15_7_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_14_LC_15_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_14_LC_15_7_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_14_LC_15_7_4  (
            .in0(N__12115),
            .in1(N__12081),
            .in2(N__11254),
            .in3(N__11251),
            .lcout(\U409_TICK.COUNTER60Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12603),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_15_LC_15_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_15_LC_15_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_15_LC_15_7_7 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_15_LC_15_7_7  (
            .in0(N__12080),
            .in1(N__12116),
            .in2(N__11233),
            .in3(N__12054),
            .lcout(\U409_TICK.COUNTER60Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12603),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_15_8_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_15_8_0 .LUT_INIT=16'b0000011111110111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_15_8_0  (
            .in0(N__11921),
            .in1(N__11909),
            .in2(N__11628),
            .in3(N__11115),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_15_8_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_15_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_15_8_1 .LUT_INIT=16'b0000001010001010;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_0_LC_15_8_1  (
            .in0(N__11846),
            .in1(N__11649),
            .in2(N__11209),
            .in3(N__11101),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_15_8_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_15_8_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_15_8_3  (
            .in0(N__11541),
            .in1(N__11601),
            .in2(_gnd_net_),
            .in3(N__11205),
            .lcout(\U409_TRANSFER_ACK.N_17_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_15_8_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_15_8_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_15_8_4  (
            .in0(N__11602),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11540),
            .lcout(\U409_TRANSFER_ACK.N_3_0 ),
            .ltout(\U409_TRANSFER_ACK.N_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_15_8_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_15_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_15_8_5 .LUT_INIT=16'b0011000001110100;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_15_8_5  (
            .in0(N__11908),
            .in1(N__11625),
            .in2(N__11104),
            .in3(N__11923),
            .lcout(\U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_15_8_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_15_8_6 .LUT_INIT=16'b0001000000011111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_15_8_6  (
            .in0(N__11922),
            .in1(N__11910),
            .in2(N__11629),
            .in3(N__11893),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.N_55_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_15_8_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_15_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_15_8_7 .LUT_INIT=16'b0010101000001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_1_LC_15_8_7  (
            .in0(N__11847),
            .in1(N__11648),
            .in2(N__11632),
            .in3(N__11626),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_15_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_15_9_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_15_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_1_LC_15_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11542),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .ce(),
            .sr(N__11391));
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_15_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_15_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_15_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_0_LC_15_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11586),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .ce(),
            .sr(N__11391));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_15_10_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_15_10_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_15_10_7 .LUT_INIT=16'b0000000011101100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_15_10_7  (
            .in0(N__11527),
            .in1(N__11518),
            .in2(N__11512),
            .in3(N__11464),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__11387));
    defparam \U409_TICK.COUNTER50_15_LC_16_5_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_15_LC_16_5_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_15_LC_16_5_1 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_15_LC_16_5_1  (
            .in0(N__12733),
            .in1(N__12704),
            .in2(N__12775),
            .in3(N__12660),
            .lcout(\U409_TICK.COUNTER50Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12601),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_13_LC_16_5_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_13_LC_16_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_13_LC_16_5_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_13_LC_16_5_2  (
            .in0(N__12702),
            .in1(N__12734),
            .in2(N__12668),
            .in3(N__12286),
            .lcout(\U409_TICK.COUNTER50Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12601),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_9_LC_16_5_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_9_LC_16_5_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_9_LC_16_5_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_9_LC_16_5_4  (
            .in0(N__12705),
            .in1(N__12736),
            .in2(N__12669),
            .in3(N__12346),
            .lcout(\U409_TICK.COUNTER50Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12601),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_16_5_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_16_5_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_16_5_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNII24V_14_LC_16_5_5  (
            .in0(N__12388),
            .in1(N__12811),
            .in2(N__12166),
            .in3(N__12787),
            .lcout(\U409_TICK.TICK503_10 ),
            .ltout(\U409_TICK.TICK503_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_14_LC_16_5_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_14_LC_16_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_14_LC_16_5_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_14_LC_16_5_6  (
            .in0(N__12703),
            .in1(N__12735),
            .in2(N__12127),
            .in3(N__12796),
            .lcout(\U409_TICK.COUNTER50Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12601),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK60_LC_16_6_4 .C_ON=1'b0;
    defparam \U409_TICK.TICK60_LC_16_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK60_LC_16_6_4 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK60_LC_16_6_4  (
            .in0(N__12123),
            .in1(N__12012),
            .in2(N__12091),
            .in3(N__12055),
            .lcout(TICK60_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12604),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_1_LC_16_6_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_1_LC_16_6_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_1_LC_16_6_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER50_1_LC_16_6_5  (
            .in0(N__12226),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12246),
            .lcout(\U409_TICK.COUNTER50Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12604),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_17_3_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_17_3_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_17_3_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_17_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_17_4_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_17_4_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_17_4_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_TICK.COUNTER50_RNID6CP_3_LC_17_4_0  (
            .in0(N__12148),
            .in1(N__12181),
            .in2(_gnd_net_),
            .in3(N__12220),
            .lcout(\U409_TICK.TICK503_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_17_4_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_17_4_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_17_4_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER50_RNIUHF01_16_LC_17_4_1  (
            .in0(N__12373),
            .in1(N__12247),
            .in2(N__12199),
            .in3(N__12757),
            .lcout(),
            .ltout(\U409_TICK.TICK503_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_17_4_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_17_4_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_17_4_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER50_RNITU182_10_LC_17_4_2  (
            .in0(N__11935),
            .in1(N__12316),
            .in2(N__11929),
            .in3(N__12337),
            .lcout(\U409_TICK.TICK503_14 ),
            .ltout(\U409_TICK.TICK503_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_6_LC_17_4_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_6_LC_17_4_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_6_LC_17_4_3 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \U409_TICK.COUNTER50_6_LC_17_4_3  (
            .in0(N__12397),
            .in1(N__12697),
            .in2(N__11926),
            .in3(N__12663),
            .lcout(\U409_TICK.COUNTER50Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12602),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK50_LC_17_4_4 .C_ON=1'b0;
    defparam \U409_TICK.TICK50_LC_17_4_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK50_LC_17_4_4 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \U409_TICK.TICK50_LC_17_4_4  (
            .in0(N__12661),
            .in1(N__12738),
            .in2(N__12706),
            .in3(N__12261),
            .lcout(TICK50_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12602),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_0_LC_17_4_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_0_LC_17_4_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_0_LC_17_4_5 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \U409_TICK.COUNTER50_0_LC_17_4_5  (
            .in0(N__12221),
            .in1(N__12696),
            .in2(N__12742),
            .in3(N__12662),
            .lcout(\U409_TICK.COUNTER50Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12602),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_17_4_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_17_4_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_17_4_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNIH14V_11_LC_17_4_6  (
            .in0(N__12298),
            .in1(N__12358),
            .in2(N__12415),
            .in3(N__12619),
            .lcout(\U409_TICK.TICK503_9 ),
            .ltout(\U409_TICK.TICK503_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_5_LC_17_4_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_5_LC_17_4_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_5_LC_17_4_7 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \U409_TICK.COUNTER50_5_LC_17_4_7  (
            .in0(N__12737),
            .in1(N__12136),
            .in2(N__12250),
            .in3(N__12664),
            .lcout(\U409_TICK.COUNTER50Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12602),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_17_5_0 .C_ON=1'b1;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_17_5_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_17_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_17_5_0  (
            .in0(_gnd_net_),
            .in1(N__12242),
            .in2(N__12225),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_5_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_2_LC_17_5_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_2_LC_17_5_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_2_LC_17_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_2_LC_17_5_1  (
            .in0(_gnd_net_),
            .in1(N__12195),
            .in2(_gnd_net_),
            .in3(N__12184),
            .lcout(\U409_TICK.COUNTER50Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .clk(N__12605),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_3_LC_17_5_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_3_LC_17_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_3_LC_17_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_3_LC_17_5_2  (
            .in0(_gnd_net_),
            .in1(N__12180),
            .in2(_gnd_net_),
            .in3(N__12169),
            .lcout(\U409_TICK.COUNTER50Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .clk(N__12605),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_4_LC_17_5_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_4_LC_17_5_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_4_LC_17_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_4_LC_17_5_3  (
            .in0(_gnd_net_),
            .in1(N__12162),
            .in2(_gnd_net_),
            .in3(N__12151),
            .lcout(\U409_TICK.COUNTER50Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .clk(N__12605),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_17_5_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_17_5_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_17_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_5_LC_17_5_4  (
            .in0(_gnd_net_),
            .in1(N__12147),
            .in2(_gnd_net_),
            .in3(N__12130),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_17_5_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_17_5_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_17_5_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_6_LC_17_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12414),
            .in3(N__12391),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_7_LC_17_5_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_7_LC_17_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_7_LC_17_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_7_LC_17_5_6  (
            .in0(_gnd_net_),
            .in1(N__12387),
            .in2(_gnd_net_),
            .in3(N__12376),
            .lcout(\U409_TICK.COUNTER50Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .clk(N__12605),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_8_LC_17_5_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_8_LC_17_5_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_8_LC_17_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_8_LC_17_5_7  (
            .in0(_gnd_net_),
            .in1(N__12372),
            .in2(_gnd_net_),
            .in3(N__12361),
            .lcout(\U409_TICK.COUNTER50Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .clk(N__12605),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_17_6_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_17_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_17_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_9_LC_17_6_0  (
            .in0(_gnd_net_),
            .in1(N__12357),
            .in2(_gnd_net_),
            .in3(N__12340),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_17_6_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_10_LC_17_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_10_LC_17_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_10_LC_17_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_10_LC_17_6_1  (
            .in0(_gnd_net_),
            .in1(N__12333),
            .in2(_gnd_net_),
            .in3(N__12322),
            .lcout(\U409_TICK.COUNTER50Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .clk(N__12606),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_17_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_17_6_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_17_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_11_LC_17_6_2  (
            .in0(_gnd_net_),
            .in1(N__12618),
            .in2(_gnd_net_),
            .in3(N__12319),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_12_LC_17_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_12_LC_17_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_12_LC_17_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_12_LC_17_6_3  (
            .in0(_gnd_net_),
            .in1(N__12312),
            .in2(_gnd_net_),
            .in3(N__12301),
            .lcout(\U409_TICK.COUNTER50Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .clk(N__12606),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_17_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_17_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_17_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_13_LC_17_6_4  (
            .in0(_gnd_net_),
            .in1(N__12297),
            .in2(_gnd_net_),
            .in3(N__12280),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_17_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_17_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_17_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_14_LC_17_6_5  (
            .in0(_gnd_net_),
            .in1(N__12810),
            .in2(_gnd_net_),
            .in3(N__12790),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_17_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_17_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_17_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_15_LC_17_6_6  (
            .in0(_gnd_net_),
            .in1(N__12786),
            .in2(_gnd_net_),
            .in3(N__12763),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_16_LC_17_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_16_LC_17_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_16_LC_17_6_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER50_16_LC_17_6_7  (
            .in0(_gnd_net_),
            .in1(N__12756),
            .in2(_gnd_net_),
            .in3(N__12760),
            .lcout(\U409_TICK.COUNTER50Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12606),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_11_LC_18_5_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_11_LC_18_5_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_11_LC_18_5_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_11_LC_18_5_3  (
            .in0(N__12732),
            .in1(N__12701),
            .in2(N__12670),
            .in3(N__12625),
            .lcout(\U409_TICK.COUNTER50Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12607),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PCS0_LC_19_2_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PCS0_LC_19_2_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PCS0_LC_19_2_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U409_ADDRESS_DECODE.PCS0_LC_19_2_5  (
            .in0(N__12528),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12471),
            .lcout(PCS0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.SCS1_LC_19_3_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.SCS1_LC_19_3_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.SCS1_LC_19_3_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \U409_ADDRESS_DECODE.SCS1_LC_19_3_2  (
            .in0(N__12472),
            .in1(N__12486),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(SCS1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PCS1_LC_20_2_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PCS1_LC_20_2_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PCS1_LC_20_2_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_ADDRESS_DECODE.PCS1_LC_20_2_2  (
            .in0(_gnd_net_),
            .in1(N__12532),
            .in2(_gnd_net_),
            .in3(N__12469),
            .lcout(PCS1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.SCS0_LC_20_3_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.SCS0_LC_20_3_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.SCS0_LC_20_3_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U409_ADDRESS_DECODE.SCS0_LC_20_3_5  (
            .in0(_gnd_net_),
            .in1(N__12487),
            .in2(_gnd_net_),
            .in3(N__12470),
            .lcout(SCS0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam AGNUS_CLK_obuf_RNO_LC_24_14_7.C_ON=1'b0;
    defparam AGNUS_CLK_obuf_RNO_LC_24_14_7.SEQ_MODE=4'b0000;
    defparam AGNUS_CLK_obuf_RNO_LC_24_14_7.LUT_INIT=16'b1110111001000100;
    LogicCell40 AGNUS_CLK_obuf_RNO_LC_24_14_7 (
            .in0(N__12874),
            .in1(N__12862),
            .in2(_gnd_net_),
            .in3(N__12850),
            .lcout(AGNUS_CLK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U409_TOP

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     May 31 2025 14:05:17

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U409_TOP" view "INTERFACE"

module U409_TOP (
    TT,
    TM,
    A,
    D,
    TICK60,
    CIACS0n,
    CLK6,
    CLK_CIA,
    BUFENn,
    RnW,
    CIACS1n,
    TICK50,
    TCIn,
    TBIn,
    RAMSPACEn,
    CLK40_IN,
    CLK28_IN,
    REGSPACEn,
    TSn,
    RTC_ENn,
    RESETn,
    OVL,
    TACKn,
    ROMENn,
    PORTSIZE);

    input [1:0] TT;
    input [1:0] TM;
    input [31:1] A;
    output [7:0] D;
    output TICK60;
    output CIACS0n;
    input CLK6;
    output CLK_CIA;
    output BUFENn;
    input RnW;
    output CIACS1n;
    output TICK50;
    output TCIn;
    output TBIn;
    output RAMSPACEn;
    input CLK40_IN;
    input CLK28_IN;
    output REGSPACEn;
    input TSn;
    output RTC_ENn;
    input RESETn;
    input OVL;
    inout TACKn;
    output ROMENn;
    output PORTSIZE;

    wire N__7928;
    wire N__7927;
    wire N__7926;
    wire N__7918;
    wire N__7917;
    wire N__7916;
    wire N__7907;
    wire N__7906;
    wire N__7905;
    wire N__7898;
    wire N__7897;
    wire N__7896;
    wire N__7889;
    wire N__7888;
    wire N__7887;
    wire N__7880;
    wire N__7879;
    wire N__7878;
    wire N__7871;
    wire N__7870;
    wire N__7869;
    wire N__7862;
    wire N__7861;
    wire N__7860;
    wire N__7853;
    wire N__7852;
    wire N__7851;
    wire N__7844;
    wire N__7843;
    wire N__7842;
    wire N__7835;
    wire N__7834;
    wire N__7833;
    wire N__7826;
    wire N__7825;
    wire N__7824;
    wire N__7817;
    wire N__7816;
    wire N__7815;
    wire N__7808;
    wire N__7807;
    wire N__7806;
    wire N__7799;
    wire N__7798;
    wire N__7797;
    wire N__7790;
    wire N__7789;
    wire N__7788;
    wire N__7781;
    wire N__7780;
    wire N__7779;
    wire N__7772;
    wire N__7771;
    wire N__7770;
    wire N__7763;
    wire N__7762;
    wire N__7761;
    wire N__7754;
    wire N__7753;
    wire N__7752;
    wire N__7745;
    wire N__7744;
    wire N__7743;
    wire N__7736;
    wire N__7735;
    wire N__7734;
    wire N__7727;
    wire N__7726;
    wire N__7725;
    wire N__7718;
    wire N__7717;
    wire N__7716;
    wire N__7709;
    wire N__7708;
    wire N__7707;
    wire N__7700;
    wire N__7699;
    wire N__7698;
    wire N__7691;
    wire N__7690;
    wire N__7689;
    wire N__7682;
    wire N__7681;
    wire N__7680;
    wire N__7673;
    wire N__7672;
    wire N__7671;
    wire N__7664;
    wire N__7663;
    wire N__7662;
    wire N__7655;
    wire N__7654;
    wire N__7653;
    wire N__7646;
    wire N__7645;
    wire N__7644;
    wire N__7637;
    wire N__7636;
    wire N__7635;
    wire N__7628;
    wire N__7627;
    wire N__7626;
    wire N__7619;
    wire N__7618;
    wire N__7617;
    wire N__7610;
    wire N__7609;
    wire N__7608;
    wire N__7601;
    wire N__7600;
    wire N__7599;
    wire N__7592;
    wire N__7591;
    wire N__7590;
    wire N__7583;
    wire N__7582;
    wire N__7581;
    wire N__7574;
    wire N__7573;
    wire N__7572;
    wire N__7565;
    wire N__7564;
    wire N__7563;
    wire N__7556;
    wire N__7555;
    wire N__7554;
    wire N__7547;
    wire N__7546;
    wire N__7545;
    wire N__7538;
    wire N__7537;
    wire N__7536;
    wire N__7529;
    wire N__7528;
    wire N__7527;
    wire N__7520;
    wire N__7519;
    wire N__7518;
    wire N__7511;
    wire N__7510;
    wire N__7509;
    wire N__7502;
    wire N__7501;
    wire N__7500;
    wire N__7493;
    wire N__7492;
    wire N__7491;
    wire N__7484;
    wire N__7483;
    wire N__7482;
    wire N__7475;
    wire N__7474;
    wire N__7473;
    wire N__7456;
    wire N__7455;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7438;
    wire N__7435;
    wire N__7432;
    wire N__7431;
    wire N__7430;
    wire N__7427;
    wire N__7422;
    wire N__7417;
    wire N__7416;
    wire N__7415;
    wire N__7414;
    wire N__7413;
    wire N__7412;
    wire N__7409;
    wire N__7406;
    wire N__7403;
    wire N__7398;
    wire N__7393;
    wire N__7384;
    wire N__7383;
    wire N__7382;
    wire N__7375;
    wire N__7372;
    wire N__7369;
    wire N__7366;
    wire N__7363;
    wire N__7360;
    wire N__7359;
    wire N__7356;
    wire N__7353;
    wire N__7348;
    wire N__7347;
    wire N__7346;
    wire N__7341;
    wire N__7338;
    wire N__7333;
    wire N__7330;
    wire N__7327;
    wire N__7326;
    wire N__7325;
    wire N__7324;
    wire N__7323;
    wire N__7322;
    wire N__7319;
    wire N__7314;
    wire N__7309;
    wire N__7306;
    wire N__7297;
    wire N__7296;
    wire N__7295;
    wire N__7294;
    wire N__7291;
    wire N__7286;
    wire N__7283;
    wire N__7276;
    wire N__7273;
    wire N__7272;
    wire N__7271;
    wire N__7270;
    wire N__7267;
    wire N__7262;
    wire N__7259;
    wire N__7252;
    wire N__7249;
    wire N__7246;
    wire N__7243;
    wire N__7242;
    wire N__7241;
    wire N__7240;
    wire N__7235;
    wire N__7232;
    wire N__7229;
    wire N__7222;
    wire N__7219;
    wire N__7218;
    wire N__7215;
    wire N__7214;
    wire N__7213;
    wire N__7210;
    wire N__7207;
    wire N__7204;
    wire N__7199;
    wire N__7192;
    wire N__7189;
    wire N__7186;
    wire N__7183;
    wire N__7180;
    wire N__7177;
    wire N__7174;
    wire N__7171;
    wire N__7170;
    wire N__7167;
    wire N__7166;
    wire N__7165;
    wire N__7162;
    wire N__7159;
    wire N__7156;
    wire N__7151;
    wire N__7144;
    wire N__7141;
    wire N__7138;
    wire N__7135;
    wire N__7132;
    wire N__7129;
    wire N__7126;
    wire N__7123;
    wire N__7122;
    wire N__7119;
    wire N__7116;
    wire N__7111;
    wire N__7108;
    wire N__7105;
    wire N__7102;
    wire N__7099;
    wire N__7096;
    wire N__7093;
    wire N__7092;
    wire N__7089;
    wire N__7086;
    wire N__7083;
    wire N__7078;
    wire N__7075;
    wire N__7072;
    wire N__7071;
    wire N__7068;
    wire N__7065;
    wire N__7060;
    wire N__7059;
    wire N__7056;
    wire N__7053;
    wire N__7048;
    wire N__7045;
    wire N__7044;
    wire N__7041;
    wire N__7038;
    wire N__7033;
    wire N__7032;
    wire N__7031;
    wire N__7030;
    wire N__7027;
    wire N__7024;
    wire N__7023;
    wire N__7020;
    wire N__7019;
    wire N__7018;
    wire N__7015;
    wire N__7014;
    wire N__7011;
    wire N__7008;
    wire N__7003;
    wire N__6994;
    wire N__6991;
    wire N__6982;
    wire N__6981;
    wire N__6980;
    wire N__6979;
    wire N__6978;
    wire N__6977;
    wire N__6976;
    wire N__6975;
    wire N__6972;
    wire N__6967;
    wire N__6962;
    wire N__6955;
    wire N__6946;
    wire N__6945;
    wire N__6944;
    wire N__6943;
    wire N__6942;
    wire N__6941;
    wire N__6940;
    wire N__6939;
    wire N__6932;
    wire N__6927;
    wire N__6924;
    wire N__6919;
    wire N__6916;
    wire N__6907;
    wire N__6904;
    wire N__6901;
    wire N__6898;
    wire N__6897;
    wire N__6894;
    wire N__6891;
    wire N__6886;
    wire N__6885;
    wire N__6884;
    wire N__6883;
    wire N__6882;
    wire N__6881;
    wire N__6880;
    wire N__6879;
    wire N__6878;
    wire N__6877;
    wire N__6876;
    wire N__6853;
    wire N__6850;
    wire N__6847;
    wire N__6844;
    wire N__6841;
    wire N__6838;
    wire N__6835;
    wire N__6834;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6820;
    wire N__6817;
    wire N__6814;
    wire N__6811;
    wire N__6810;
    wire N__6807;
    wire N__6804;
    wire N__6803;
    wire N__6800;
    wire N__6797;
    wire N__6794;
    wire N__6791;
    wire N__6788;
    wire N__6785;
    wire N__6778;
    wire N__6775;
    wire N__6774;
    wire N__6771;
    wire N__6768;
    wire N__6765;
    wire N__6764;
    wire N__6761;
    wire N__6758;
    wire N__6755;
    wire N__6748;
    wire N__6747;
    wire N__6744;
    wire N__6741;
    wire N__6736;
    wire N__6733;
    wire N__6730;
    wire N__6727;
    wire N__6724;
    wire N__6723;
    wire N__6720;
    wire N__6717;
    wire N__6712;
    wire N__6709;
    wire N__6706;
    wire N__6703;
    wire N__6700;
    wire N__6697;
    wire N__6694;
    wire N__6693;
    wire N__6690;
    wire N__6687;
    wire N__6682;
    wire N__6679;
    wire N__6678;
    wire N__6675;
    wire N__6672;
    wire N__6669;
    wire N__6666;
    wire N__6661;
    wire N__6658;
    wire N__6655;
    wire N__6652;
    wire N__6649;
    wire N__6646;
    wire N__6645;
    wire N__6642;
    wire N__6639;
    wire N__6634;
    wire N__6631;
    wire N__6630;
    wire N__6627;
    wire N__6624;
    wire N__6619;
    wire N__6616;
    wire N__6613;
    wire N__6610;
    wire N__6607;
    wire N__6606;
    wire N__6603;
    wire N__6600;
    wire N__6595;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6579;
    wire N__6578;
    wire N__6577;
    wire N__6574;
    wire N__6569;
    wire N__6566;
    wire N__6559;
    wire N__6558;
    wire N__6557;
    wire N__6554;
    wire N__6551;
    wire N__6548;
    wire N__6545;
    wire N__6538;
    wire N__6537;
    wire N__6534;
    wire N__6531;
    wire N__6526;
    wire N__6523;
    wire N__6522;
    wire N__6519;
    wire N__6516;
    wire N__6511;
    wire N__6508;
    wire N__6505;
    wire N__6502;
    wire N__6501;
    wire N__6500;
    wire N__6499;
    wire N__6496;
    wire N__6491;
    wire N__6488;
    wire N__6485;
    wire N__6482;
    wire N__6475;
    wire N__6472;
    wire N__6471;
    wire N__6470;
    wire N__6467;
    wire N__6462;
    wire N__6459;
    wire N__6456;
    wire N__6451;
    wire N__6450;
    wire N__6447;
    wire N__6446;
    wire N__6443;
    wire N__6442;
    wire N__6441;
    wire N__6438;
    wire N__6435;
    wire N__6434;
    wire N__6431;
    wire N__6428;
    wire N__6425;
    wire N__6420;
    wire N__6417;
    wire N__6412;
    wire N__6409;
    wire N__6408;
    wire N__6403;
    wire N__6400;
    wire N__6397;
    wire N__6394;
    wire N__6391;
    wire N__6382;
    wire N__6379;
    wire N__6378;
    wire N__6375;
    wire N__6372;
    wire N__6367;
    wire N__6364;
    wire N__6361;
    wire N__6360;
    wire N__6357;
    wire N__6354;
    wire N__6353;
    wire N__6348;
    wire N__6345;
    wire N__6342;
    wire N__6339;
    wire N__6334;
    wire N__6333;
    wire N__6330;
    wire N__6327;
    wire N__6326;
    wire N__6323;
    wire N__6320;
    wire N__6317;
    wire N__6314;
    wire N__6311;
    wire N__6308;
    wire N__6305;
    wire N__6300;
    wire N__6295;
    wire N__6292;
    wire N__6289;
    wire N__6286;
    wire N__6283;
    wire N__6280;
    wire N__6277;
    wire N__6274;
    wire N__6271;
    wire N__6268;
    wire N__6265;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6253;
    wire N__6250;
    wire N__6247;
    wire N__6244;
    wire N__6243;
    wire N__6242;
    wire N__6239;
    wire N__6236;
    wire N__6233;
    wire N__6232;
    wire N__6227;
    wire N__6226;
    wire N__6225;
    wire N__6222;
    wire N__6219;
    wire N__6216;
    wire N__6213;
    wire N__6212;
    wire N__6209;
    wire N__6208;
    wire N__6207;
    wire N__6204;
    wire N__6201;
    wire N__6196;
    wire N__6189;
    wire N__6188;
    wire N__6187;
    wire N__6186;
    wire N__6185;
    wire N__6182;
    wire N__6179;
    wire N__6176;
    wire N__6171;
    wire N__6168;
    wire N__6165;
    wire N__6162;
    wire N__6159;
    wire N__6156;
    wire N__6151;
    wire N__6142;
    wire N__6139;
    wire N__6134;
    wire N__6131;
    wire N__6128;
    wire N__6121;
    wire N__6118;
    wire N__6115;
    wire N__6112;
    wire N__6109;
    wire N__6106;
    wire N__6103;
    wire N__6100;
    wire N__6097;
    wire N__6094;
    wire N__6091;
    wire N__6088;
    wire N__6085;
    wire N__6082;
    wire N__6079;
    wire N__6076;
    wire N__6073;
    wire N__6070;
    wire N__6067;
    wire N__6064;
    wire N__6063;
    wire N__6060;
    wire N__6057;
    wire N__6052;
    wire N__6051;
    wire N__6048;
    wire N__6045;
    wire N__6040;
    wire N__6039;
    wire N__6038;
    wire N__6035;
    wire N__6032;
    wire N__6029;
    wire N__6026;
    wire N__6023;
    wire N__6016;
    wire N__6015;
    wire N__6012;
    wire N__6009;
    wire N__6004;
    wire N__6003;
    wire N__6000;
    wire N__5997;
    wire N__5992;
    wire N__5989;
    wire N__5986;
    wire N__5983;
    wire N__5982;
    wire N__5979;
    wire N__5976;
    wire N__5971;
    wire N__5968;
    wire N__5965;
    wire N__5962;
    wire N__5961;
    wire N__5958;
    wire N__5955;
    wire N__5950;
    wire N__5949;
    wire N__5946;
    wire N__5943;
    wire N__5938;
    wire N__5935;
    wire N__5934;
    wire N__5931;
    wire N__5928;
    wire N__5923;
    wire N__5920;
    wire N__5917;
    wire N__5914;
    wire N__5913;
    wire N__5910;
    wire N__5907;
    wire N__5902;
    wire N__5901;
    wire N__5898;
    wire N__5895;
    wire N__5890;
    wire N__5889;
    wire N__5886;
    wire N__5883;
    wire N__5878;
    wire N__5875;
    wire N__5874;
    wire N__5871;
    wire N__5868;
    wire N__5863;
    wire N__5860;
    wire N__5857;
    wire N__5854;
    wire N__5853;
    wire N__5850;
    wire N__5847;
    wire N__5842;
    wire N__5841;
    wire N__5840;
    wire N__5839;
    wire N__5838;
    wire N__5837;
    wire N__5836;
    wire N__5833;
    wire N__5828;
    wire N__5823;
    wire N__5818;
    wire N__5809;
    wire N__5808;
    wire N__5805;
    wire N__5802;
    wire N__5801;
    wire N__5800;
    wire N__5799;
    wire N__5798;
    wire N__5797;
    wire N__5794;
    wire N__5789;
    wire N__5784;
    wire N__5779;
    wire N__5770;
    wire N__5769;
    wire N__5768;
    wire N__5767;
    wire N__5766;
    wire N__5765;
    wire N__5762;
    wire N__5759;
    wire N__5758;
    wire N__5755;
    wire N__5750;
    wire N__5747;
    wire N__5744;
    wire N__5739;
    wire N__5736;
    wire N__5733;
    wire N__5730;
    wire N__5719;
    wire N__5716;
    wire N__5713;
    wire N__5712;
    wire N__5709;
    wire N__5706;
    wire N__5701;
    wire N__5698;
    wire N__5697;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5689;
    wire N__5688;
    wire N__5685;
    wire N__5680;
    wire N__5673;
    wire N__5670;
    wire N__5665;
    wire N__5662;
    wire N__5659;
    wire N__5656;
    wire N__5653;
    wire N__5650;
    wire N__5647;
    wire N__5646;
    wire N__5643;
    wire N__5640;
    wire N__5635;
    wire N__5632;
    wire N__5629;
    wire N__5626;
    wire N__5625;
    wire N__5622;
    wire N__5621;
    wire N__5618;
    wire N__5617;
    wire N__5614;
    wire N__5609;
    wire N__5606;
    wire N__5599;
    wire N__5598;
    wire N__5597;
    wire N__5592;
    wire N__5589;
    wire N__5584;
    wire N__5581;
    wire N__5578;
    wire N__5577;
    wire N__5576;
    wire N__5575;
    wire N__5572;
    wire N__5569;
    wire N__5564;
    wire N__5561;
    wire N__5554;
    wire N__5551;
    wire N__5548;
    wire N__5547;
    wire N__5546;
    wire N__5543;
    wire N__5542;
    wire N__5541;
    wire N__5538;
    wire N__5535;
    wire N__5534;
    wire N__5531;
    wire N__5528;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5518;
    wire N__5515;
    wire N__5512;
    wire N__5507;
    wire N__5500;
    wire N__5497;
    wire N__5496;
    wire N__5493;
    wire N__5490;
    wire N__5487;
    wire N__5484;
    wire N__5481;
    wire N__5478;
    wire N__5475;
    wire N__5470;
    wire N__5467;
    wire N__5458;
    wire N__5455;
    wire N__5452;
    wire N__5449;
    wire N__5446;
    wire N__5443;
    wire N__5440;
    wire N__5437;
    wire N__5434;
    wire N__5431;
    wire N__5428;
    wire N__5427;
    wire N__5424;
    wire N__5421;
    wire N__5416;
    wire N__5413;
    wire N__5410;
    wire N__5409;
    wire N__5406;
    wire N__5403;
    wire N__5402;
    wire N__5397;
    wire N__5394;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5361;
    wire N__5358;
    wire N__5355;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5332;
    wire N__5329;
    wire N__5326;
    wire N__5323;
    wire N__5320;
    wire N__5319;
    wire N__5318;
    wire N__5317;
    wire N__5314;
    wire N__5309;
    wire N__5306;
    wire N__5305;
    wire N__5304;
    wire N__5303;
    wire N__5296;
    wire N__5293;
    wire N__5290;
    wire N__5287;
    wire N__5282;
    wire N__5275;
    wire N__5274;
    wire N__5273;
    wire N__5270;
    wire N__5269;
    wire N__5268;
    wire N__5265;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5252;
    wire N__5251;
    wire N__5246;
    wire N__5241;
    wire N__5236;
    wire N__5233;
    wire N__5224;
    wire N__5223;
    wire N__5220;
    wire N__5219;
    wire N__5216;
    wire N__5215;
    wire N__5214;
    wire N__5213;
    wire N__5206;
    wire N__5203;
    wire N__5202;
    wire N__5201;
    wire N__5198;
    wire N__5195;
    wire N__5190;
    wire N__5185;
    wire N__5182;
    wire N__5179;
    wire N__5176;
    wire N__5167;
    wire N__5164;
    wire N__5163;
    wire N__5162;
    wire N__5161;
    wire N__5160;
    wire N__5157;
    wire N__5154;
    wire N__5151;
    wire N__5150;
    wire N__5145;
    wire N__5142;
    wire N__5137;
    wire N__5134;
    wire N__5125;
    wire N__5122;
    wire N__5119;
    wire N__5116;
    wire N__5113;
    wire N__5112;
    wire N__5111;
    wire N__5110;
    wire N__5103;
    wire N__5100;
    wire N__5095;
    wire N__5092;
    wire N__5089;
    wire N__5088;
    wire N__5087;
    wire N__5086;
    wire N__5083;
    wire N__5080;
    wire N__5077;
    wire N__5074;
    wire N__5073;
    wire N__5062;
    wire N__5059;
    wire N__5058;
    wire N__5057;
    wire N__5056;
    wire N__5053;
    wire N__5050;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5029;
    wire N__5028;
    wire N__5027;
    wire N__5026;
    wire N__5023;
    wire N__5020;
    wire N__5015;
    wire N__5008;
    wire N__5007;
    wire N__5002;
    wire N__4999;
    wire N__4998;
    wire N__4997;
    wire N__4996;
    wire N__4995;
    wire N__4994;
    wire N__4993;
    wire N__4988;
    wire N__4985;
    wire N__4982;
    wire N__4979;
    wire N__4974;
    wire N__4963;
    wire N__4962;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4945;
    wire N__4944;
    wire N__4943;
    wire N__4942;
    wire N__4937;
    wire N__4934;
    wire N__4931;
    wire N__4924;
    wire N__4923;
    wire N__4922;
    wire N__4919;
    wire N__4916;
    wire N__4913;
    wire N__4910;
    wire N__4907;
    wire N__4900;
    wire N__4899;
    wire N__4898;
    wire N__4897;
    wire N__4892;
    wire N__4891;
    wire N__4890;
    wire N__4887;
    wire N__4884;
    wire N__4881;
    wire N__4876;
    wire N__4867;
    wire N__4864;
    wire N__4863;
    wire N__4862;
    wire N__4861;
    wire N__4860;
    wire N__4857;
    wire N__4852;
    wire N__4847;
    wire N__4840;
    wire N__4837;
    wire N__4834;
    wire N__4831;
    wire N__4830;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4815;
    wire N__4812;
    wire N__4811;
    wire N__4806;
    wire N__4803;
    wire N__4798;
    wire N__4795;
    wire N__4792;
    wire N__4789;
    wire N__4788;
    wire N__4785;
    wire N__4782;
    wire N__4779;
    wire N__4776;
    wire N__4771;
    wire N__4768;
    wire N__4765;
    wire N__4762;
    wire N__4759;
    wire N__4756;
    wire N__4753;
    wire N__4750;
    wire N__4747;
    wire N__4746;
    wire N__4743;
    wire N__4740;
    wire N__4739;
    wire N__4736;
    wire N__4733;
    wire N__4730;
    wire N__4727;
    wire N__4722;
    wire N__4721;
    wire N__4716;
    wire N__4713;
    wire N__4708;
    wire N__4705;
    wire N__4702;
    wire N__4699;
    wire N__4696;
    wire N__4693;
    wire N__4690;
    wire N__4687;
    wire N__4684;
    wire N__4681;
    wire N__4678;
    wire N__4675;
    wire N__4672;
    wire N__4669;
    wire N__4668;
    wire N__4665;
    wire N__4662;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4648;
    wire N__4645;
    wire N__4642;
    wire N__4639;
    wire N__4636;
    wire N__4635;
    wire N__4630;
    wire N__4627;
    wire N__4624;
    wire N__4623;
    wire N__4620;
    wire N__4617;
    wire N__4612;
    wire N__4609;
    wire N__4608;
    wire N__4605;
    wire N__4604;
    wire N__4603;
    wire N__4600;
    wire N__4597;
    wire N__4592;
    wire N__4585;
    wire N__4582;
    wire N__4579;
    wire N__4576;
    wire N__4573;
    wire N__4570;
    wire N__4569;
    wire N__4564;
    wire N__4561;
    wire N__4558;
    wire N__4555;
    wire N__4554;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4543;
    wire N__4538;
    wire N__4533;
    wire N__4532;
    wire N__4527;
    wire N__4524;
    wire N__4521;
    wire N__4518;
    wire N__4515;
    wire N__4512;
    wire N__4509;
    wire N__4506;
    wire N__4503;
    wire N__4498;
    wire N__4497;
    wire N__4496;
    wire N__4493;
    wire N__4488;
    wire N__4483;
    wire N__4480;
    wire N__4477;
    wire N__4474;
    wire N__4471;
    wire N__4468;
    wire N__4465;
    wire N__4462;
    wire N__4459;
    wire N__4456;
    wire N__4453;
    wire N__4450;
    wire N__4447;
    wire N__4446;
    wire N__4443;
    wire N__4440;
    wire N__4439;
    wire N__4438;
    wire N__4437;
    wire N__4432;
    wire N__4429;
    wire N__4426;
    wire N__4425;
    wire N__4424;
    wire N__4423;
    wire N__4420;
    wire N__4417;
    wire N__4412;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4395;
    wire N__4390;
    wire N__4389;
    wire N__4386;
    wire N__4383;
    wire N__4378;
    wire N__4375;
    wire N__4366;
    wire N__4363;
    wire N__4362;
    wire N__4359;
    wire N__4356;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4343;
    wire N__4338;
    wire N__4333;
    wire N__4330;
    wire N__4327;
    wire N__4324;
    wire N__4321;
    wire N__4320;
    wire N__4317;
    wire N__4314;
    wire N__4309;
    wire N__4308;
    wire N__4305;
    wire N__4302;
    wire N__4297;
    wire N__4294;
    wire N__4291;
    wire N__4290;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4276;
    wire N__4273;
    wire N__4270;
    wire N__4267;
    wire N__4264;
    wire N__4261;
    wire N__4258;
    wire N__4255;
    wire N__4252;
    wire N__4249;
    wire N__4246;
    wire N__4243;
    wire N__4240;
    wire N__4239;
    wire N__4238;
    wire N__4235;
    wire N__4232;
    wire N__4229;
    wire N__4226;
    wire N__4221;
    wire N__4218;
    wire N__4215;
    wire N__4212;
    wire N__4209;
    wire N__4206;
    wire N__4205;
    wire N__4204;
    wire N__4201;
    wire N__4198;
    wire N__4195;
    wire N__4192;
    wire N__4183;
    wire N__4182;
    wire N__4181;
    wire N__4180;
    wire N__4177;
    wire N__4170;
    wire N__4165;
    wire N__4162;
    wire N__4161;
    wire N__4160;
    wire N__4159;
    wire N__4156;
    wire N__4153;
    wire N__4148;
    wire N__4141;
    wire N__4140;
    wire N__4137;
    wire N__4134;
    wire N__4129;
    wire N__4126;
    wire N__4123;
    wire N__4120;
    wire N__4117;
    wire N__4114;
    wire N__4111;
    wire N__4108;
    wire N__4107;
    wire N__4104;
    wire N__4101;
    wire N__4096;
    wire N__4095;
    wire N__4092;
    wire N__4089;
    wire N__4084;
    wire N__4083;
    wire N__4082;
    wire N__4081;
    wire N__4078;
    wire N__4073;
    wire N__4070;
    wire N__4063;
    wire N__4060;
    wire N__4057;
    wire N__4054;
    wire N__4051;
    wire N__4048;
    wire N__4047;
    wire N__4046;
    wire N__4045;
    wire N__4042;
    wire N__4037;
    wire N__4034;
    wire N__4027;
    wire N__4024;
    wire N__4021;
    wire N__4018;
    wire N__4015;
    wire N__4014;
    wire N__4013;
    wire N__4012;
    wire N__4007;
    wire N__4004;
    wire N__4001;
    wire N__3998;
    wire N__3995;
    wire N__3994;
    wire N__3993;
    wire N__3990;
    wire N__3989;
    wire N__3984;
    wire N__3981;
    wire N__3978;
    wire N__3975;
    wire N__3972;
    wire N__3965;
    wire N__3960;
    wire N__3955;
    wire N__3954;
    wire N__3953;
    wire N__3950;
    wire N__3947;
    wire N__3944;
    wire N__3943;
    wire N__3942;
    wire N__3941;
    wire N__3940;
    wire N__3935;
    wire N__3932;
    wire N__3929;
    wire N__3926;
    wire N__3921;
    wire N__3920;
    wire N__3913;
    wire N__3908;
    wire N__3905;
    wire N__3902;
    wire N__3897;
    wire N__3894;
    wire N__3891;
    wire N__3888;
    wire N__3883;
    wire N__3880;
    wire N__3877;
    wire N__3874;
    wire N__3871;
    wire N__3868;
    wire N__3865;
    wire N__3862;
    wire N__3859;
    wire N__3856;
    wire N__3855;
    wire N__3854;
    wire N__3853;
    wire N__3852;
    wire N__3847;
    wire N__3844;
    wire N__3839;
    wire N__3836;
    wire N__3833;
    wire N__3830;
    wire N__3827;
    wire N__3822;
    wire N__3819;
    wire N__3816;
    wire N__3811;
    wire N__3808;
    wire N__3807;
    wire N__3802;
    wire N__3799;
    wire N__3796;
    wire N__3793;
    wire N__3792;
    wire N__3789;
    wire N__3784;
    wire N__3781;
    wire N__3778;
    wire N__3777;
    wire N__3772;
    wire N__3769;
    wire N__3766;
    wire N__3765;
    wire N__3762;
    wire N__3759;
    wire N__3754;
    wire N__3751;
    wire N__3748;
    wire N__3745;
    wire N__3742;
    wire N__3739;
    wire N__3736;
    wire N__3733;
    wire N__3730;
    wire N__3727;
    wire N__3724;
    wire N__3721;
    wire N__3718;
    wire N__3715;
    wire N__3712;
    wire N__3709;
    wire N__3706;
    wire N__3703;
    wire N__3700;
    wire N__3697;
    wire N__3694;
    wire N__3691;
    wire N__3688;
    wire N__3685;
    wire N__3682;
    wire N__3679;
    wire N__3676;
    wire N__3673;
    wire N__3670;
    wire N__3667;
    wire N__3666;
    wire N__3663;
    wire N__3660;
    wire N__3655;
    wire N__3654;
    wire N__3651;
    wire N__3648;
    wire N__3647;
    wire N__3646;
    wire N__3645;
    wire N__3642;
    wire N__3639;
    wire N__3634;
    wire N__3631;
    wire N__3628;
    wire N__3625;
    wire N__3620;
    wire N__3617;
    wire N__3612;
    wire N__3607;
    wire N__3604;
    wire N__3601;
    wire N__3598;
    wire N__3597;
    wire N__3596;
    wire N__3595;
    wire N__3590;
    wire N__3585;
    wire N__3584;
    wire N__3583;
    wire N__3580;
    wire N__3579;
    wire N__3576;
    wire N__3573;
    wire N__3570;
    wire N__3569;
    wire N__3566;
    wire N__3563;
    wire N__3560;
    wire N__3557;
    wire N__3554;
    wire N__3551;
    wire N__3546;
    wire N__3539;
    wire N__3536;
    wire N__3529;
    wire N__3526;
    wire N__3525;
    wire N__3522;
    wire N__3521;
    wire N__3518;
    wire N__3515;
    wire N__3512;
    wire N__3511;
    wire N__3510;
    wire N__3503;
    wire N__3500;
    wire N__3499;
    wire N__3498;
    wire N__3495;
    wire N__3492;
    wire N__3489;
    wire N__3484;
    wire N__3481;
    wire N__3478;
    wire N__3471;
    wire N__3468;
    wire N__3465;
    wire N__3462;
    wire N__3459;
    wire N__3454;
    wire N__3451;
    wire N__3448;
    wire N__3447;
    wire N__3442;
    wire N__3441;
    wire N__3438;
    wire N__3435;
    wire N__3432;
    wire N__3429;
    wire N__3428;
    wire N__3423;
    wire N__3420;
    wire N__3417;
    wire N__3414;
    wire N__3409;
    wire N__3406;
    wire N__3403;
    wire N__3400;
    wire N__3397;
    wire N__3396;
    wire N__3393;
    wire N__3390;
    wire N__3385;
    wire N__3382;
    wire N__3381;
    wire N__3378;
    wire N__3373;
    wire N__3370;
    wire N__3367;
    wire N__3364;
    wire N__3363;
    wire N__3358;
    wire N__3355;
    wire N__3352;
    wire N__3349;
    wire N__3346;
    wire N__3343;
    wire N__3340;
    wire N__3337;
    wire N__3334;
    wire N__3331;
    wire N__3328;
    wire N__3325;
    wire N__3324;
    wire N__3323;
    wire N__3322;
    wire N__3319;
    wire N__3316;
    wire N__3313;
    wire N__3310;
    wire N__3309;
    wire N__3308;
    wire N__3307;
    wire N__3300;
    wire N__3297;
    wire N__3294;
    wire N__3291;
    wire N__3288;
    wire N__3281;
    wire N__3276;
    wire N__3275;
    wire N__3270;
    wire N__3267;
    wire N__3262;
    wire N__3259;
    wire N__3256;
    wire N__3253;
    wire N__3250;
    wire N__3247;
    wire N__3244;
    wire N__3241;
    wire N__3238;
    wire N__3235;
    wire N__3232;
    wire N__3229;
    wire N__3226;
    wire N__3223;
    wire N__3220;
    wire N__3217;
    wire N__3214;
    wire N__3211;
    wire N__3208;
    wire N__3205;
    wire N__3202;
    wire N__3199;
    wire N__3196;
    wire N__3193;
    wire N__3190;
    wire N__3187;
    wire N__3184;
    wire N__3181;
    wire N__3178;
    wire N__3175;
    wire N__3172;
    wire N__3169;
    wire N__3166;
    wire N__3163;
    wire N__3160;
    wire N__3159;
    wire N__3154;
    wire N__3151;
    wire N__3148;
    wire N__3145;
    wire N__3142;
    wire N__3141;
    wire N__3136;
    wire N__3133;
    wire N__3130;
    wire N__3127;
    wire N__3124;
    wire N__3123;
    wire N__3120;
    wire N__3115;
    wire N__3112;
    wire N__3109;
    wire N__3106;
    wire N__3103;
    wire N__3100;
    wire N__3099;
    wire N__3094;
    wire N__3091;
    wire N__3088;
    wire N__3085;
    wire N__3082;
    wire N__3079;
    wire N__3076;
    wire N__3075;
    wire N__3072;
    wire N__3069;
    wire N__3064;
    wire N__3061;
    wire N__3058;
    wire N__3055;
    wire N__3052;
    wire N__3049;
    wire N__3046;
    wire N__3043;
    wire N__3042;
    wire N__3037;
    wire N__3034;
    wire N__3031;
    wire N__3028;
    wire N__3025;
    wire N__3024;
    wire N__3021;
    wire N__3016;
    wire N__3013;
    wire N__3010;
    wire N__3007;
    wire N__3004;
    wire N__3001;
    wire N__3000;
    wire N__2995;
    wire N__2992;
    wire N__2989;
    wire N__2986;
    wire N__2983;
    wire N__2980;
    wire N__2979;
    wire N__2976;
    wire N__2973;
    wire N__2968;
    wire N__2965;
    wire N__2962;
    wire N__2959;
    wire N__2958;
    wire N__2957;
    wire N__2956;
    wire N__2955;
    wire N__2954;
    wire N__2953;
    wire N__2952;
    wire N__2951;
    wire N__2950;
    wire N__2949;
    wire N__2948;
    wire N__2947;
    wire N__2920;
    wire CLK80_OUT;
    wire GNDG0;
    wire VCCG0;
    wire A_c_27;
    wire A_c_26;
    wire A_c_25;
    wire A_c_24;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5 ;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_ ;
    wire A_c_31;
    wire A_c_30;
    wire A_c_28;
    wire A_c_29;
    wire \U409_ADDRESS_DECODE.CIA_SPACE_0Z0Z_1_cascade_ ;
    wire A_c_16;
    wire \U409_ADDRESS_DECODE.RAN_SPACEZ0Z_0_cascade_ ;
    wire \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_4 ;
    wire \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_5 ;
    wire \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_0_cascade_ ;
    wire RnW_c;
    wire D_1_i;
    wire U409_ADDRESS_DECODE_un1_RTC_ENn_i;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3 ;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3_cascade_ ;
    wire \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_0 ;
    wire \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_5 ;
    wire U409_ADDRESS_DECODE_LOWROM_3_cascade_;
    wire \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_3 ;
    wire U409_ADDRESS_DECODE_AUTOVECTOR_3;
    wire TT_c_1;
    wire TT_c_0;
    wire U409_ADDRESS_DECODE_AUTOVECTOR_2;
    wire U409_ADDRESS_DECODE_LOWROM_2_cascade_;
    wire \U409_TRANSFER_ACK.N_45 ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2Z0Z_1_cascade_ ;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2 ;
    wire A_c_18;
    wire A_c_20;
    wire A_c_19;
    wire A_c_17;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_0 ;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4_cascade_ ;
    wire TM_c_1;
    wire TM_c_0;
    wire A_c_23;
    wire A_c_22;
    wire U409_ADDRESS_DECODE_un1_REGSPACEn_i;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0 ;
    wire \U409_ADDRESS_DECODE.un2_REGSPACEn_0_0 ;
    wire \U409_ADDRESS_DECODE.REG_SPACE_3_0 ;
    wire \U409_ADDRESS_DECODE.REG_SPACEZ0Z_2 ;
    wire U409_ADDRESS_DECODE_un1_RTC_ENn;
    wire PORTSIZE_0_i;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0_0_cascade_ ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_EN_nerC_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ;
    wire \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ;
    wire TACK_OUTn;
    wire \INVU409_TRANSFER_ACK.TACK_OUTnC_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER6 ;
    wire \U409_TRANSFER_ACK.N_35 ;
    wire ROMENn_c;
    wire \U409_TRANSFER_ACK.CIA_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.ROM_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.IRQ_TACK_EN_nesrC_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ;
    wire \U409_TRANSFER_ACK.N_47 ;
    wire \U409_TRANSFER_ACK.N_142 ;
    wire \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_0 ;
    wire TSn_c;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_cascade_ ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1_0 ;
    wire U409_ADDRESS_DECODE_un1_RAMSPACEn_i;
    wire A_c_21;
    wire OVL_c;
    wire U409_ADDRESS_DECODE_LOWROM_3;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_3_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_2_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5 ;
    wire U409_ADDRESS_DECODE_ROMEN_1;
    wire \U409_TRANSFER_ACK.N_23 ;
    wire TACKn_in;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ;
    wire CONSTANT_ONE_NET;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_1_0 ;
    wire \U409_TRANSFER_ACK.N_35_1 ;
    wire \U409_TRANSFER_ACK.N_29 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.N_36 ;
    wire \U409_TICK.COUNTER60Z0Z_0 ;
    wire bfn_12_9_0_;
    wire \U409_TICK.un3_COUNTER60_1_cry_1 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_2 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_3 ;
    wire \U409_TICK.COUNTER60Z0Z_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_4 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_6 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_8 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_8 ;
    wire bfn_12_10_0_;
    wire \U409_TICK.un3_COUNTER60_1_cry_9 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_10 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_13 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_15 ;
    wire U409_ADDRESS_DECODE_un1_RAMSPACEn;
    wire U409_ADDRESS_DECODE_un1_REGSPACEn;
    wire BUFENn_c;
    wire \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ;
    wire \U409_TRANSFER_ACK.i6_mux_0_cascade_ ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ;
    wire \U409_TRANSFER_ACK.N_9_cascade_ ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_1C_net ;
    wire TICK60_c;
    wire \U409_TRANSFER_ACK.N_4 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ;
    wire \U409_TRANSFER_ACK.N_4_cascade_ ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ;
    wire \U409_TRANSFER_ACK.N_5 ;
    wire CLK40_IN_c;
    wire \U409_TRANSFER_ACK.m8_ns_1 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_6 ;
    wire \U409_TICK.COUNTER60Z0Z_12 ;
    wire \U409_TICK.COUNTER60Z0Z_2 ;
    wire \U409_TICK.COUNTER60Z0Z_1 ;
    wire \U409_TICK.COUNTER60Z0Z_16 ;
    wire \U409_TICK.COUNTER60Z0Z_11 ;
    wire \U409_TICK.TICK603_8 ;
    wire \U409_TICK.TICK603_11_cascade_ ;
    wire \U409_TICK.COUNTER60Z0Z_3 ;
    wire \U409_TICK.TICK603_14_cascade_ ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_4 ;
    wire \U409_TICK.COUNTER60Z0Z_4 ;
    wire \U409_TICK.COUNTER60Z0Z_8 ;
    wire \U409_TICK.COUNTER60Z0Z_6 ;
    wire \U409_TICK.TICK603_9_cascade_ ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_14 ;
    wire \U409_TICK.COUNTER60Z0Z_14 ;
    wire \U409_TICK.COUNTER60Z0Z_13 ;
    wire \U409_TICK.COUNTER60Z0Z_10 ;
    wire \U409_TICK.COUNTER60Z0Z_7 ;
    wire \U409_TICK.TICK603_10_cascade_ ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER60Z0Z_15 ;
    wire \U409_TICK.TICK603_9 ;
    wire \U409_TICK.TICK603_14 ;
    wire \U409_TICK.TICK603_10 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_9 ;
    wire \U409_TICK.COUNTER60Z0Z_9 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_0 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.LASTCLK_0C_net ;
    wire RESETn_c_i;
    wire TACK_EN;
    wire AUTOCONFIG_SPACE;
    wire TCIn_1_i;
    wire A_c_13;
    wire U409_ADDRESS_DECODE_un1_CIACS1n_i;
    wire RESETn_c;
    wire CIA_ENABLE;
    wire A_c_12;
    wire CIA_ENABLE_cascade_;
    wire U409_ADDRESS_DECODE_un1_CIACS0n_i;
    wire \U409_TICK.TICK503_11_cascade_ ;
    wire \U409_TICK.TICK503_14_cascade_ ;
    wire \U409_TICK.TICK503_8 ;
    wire \U409_TICK.TICK503_9_cascade_ ;
    wire \U409_TICK.COUNTER50Z0Z_0 ;
    wire \U409_TICK.COUNTER50Z0Z_1 ;
    wire bfn_14_9_0_;
    wire \U409_TICK.COUNTER50Z0Z_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_1 ;
    wire \U409_TICK.COUNTER50Z0Z_3 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_3 ;
    wire \U409_TICK.COUNTER50Z0Z_5 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_4 ;
    wire \U409_TICK.COUNTER50Z0Z_6 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_6 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_6 ;
    wire \U409_TICK.COUNTER50Z0Z_8 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_8 ;
    wire \U409_TICK.COUNTER50Z0Z_9 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_9 ;
    wire bfn_14_10_0_;
    wire \U409_TICK.COUNTER50Z0Z_10 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_9 ;
    wire \U409_TICK.COUNTER50Z0Z_11 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_11 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_10 ;
    wire \U409_TICK.COUNTER50Z0Z_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_11 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_13 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_15 ;
    wire \U409_TICK.COUNTER50Z0Z_16 ;
    wire \U409_CIA.CLK_CIA6_3_cascade_ ;
    wire \U409_CIA.un1_CIA_CLK_COUNT_3_2_cascade_ ;
    wire CIA_SPACE;
    wire \U409_CIA.VMA_RNOZ0Z_0_cascade_ ;
    wire \U409_CIA.VMAZ0 ;
    wire CLK_CIA_c;
    wire \U409_CIA.CLK_CIA_r_1_0 ;
    wire TICK50_c;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_13 ;
    wire \U409_TICK.COUNTER50Z0Z_13 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_14 ;
    wire \U409_TICK.COUNTER50Z0Z_14 ;
    wire \U409_TICK.COUNTER50Z0Z_4 ;
    wire \U409_TICK.COUNTER50Z0Z_7 ;
    wire \U409_TICK.TICK503_10 ;
    wire \U409_TICK.TICK503_9 ;
    wire \U409_TICK.TICK503_14 ;
    wire \U409_TICK.TICK503_10_cascade_ ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER50Z0Z_15 ;
    wire CLK6_c_g;
    wire \U409_CIA.CIA_CLK_COUNT11_2 ;
    wire \U409_CIA.CIA_CLK_COUNT11_2_0 ;
    wire \U409_CIA.CLK_CIA6_4 ;
    wire \U409_CIA.CIA_CLK_COUNT11_2_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_1 ;
    wire bfn_15_11_0_;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_1 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_3 ;
    wire \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_4 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_3 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_5 ;
    wire \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_6 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_5 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_6 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_7 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_0 ;
    wire CLK28_IN_c_g;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="SIMPLE";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0001111;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE pll (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__5548),
            .RESETB(N__4699),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(CLK80_OUT));
    PRE_IO_GBUF CLK28_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__7926),
            .GLOBALBUFFEROUTPUT(CLK28_IN_c_g));
    IO_PAD CLK28_IN_ibuf_gb_io_iopad (
            .OE(N__7928),
            .DIN(N__7927),
            .DOUT(N__7926),
            .PACKAGEPIN(CLK28_IN));
    defparam CLK28_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK28_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK28_IN_ibuf_gb_io_preio (
            .PADOEN(N__7928),
            .PADOUT(N__7927),
            .PADIN(N__7926),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK6_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__7916),
            .GLOBALBUFFEROUTPUT(CLK6_c_g));
    IO_PAD CLK6_ibuf_gb_io_iopad (
            .OE(N__7918),
            .DIN(N__7917),
            .DOUT(N__7916),
            .PACKAGEPIN(CLK6));
    defparam CLK6_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK6_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK6_ibuf_gb_io_preio (
            .PADOEN(N__7918),
            .PADOUT(N__7917),
            .PADIN(N__7916),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_0_iopad (
            .OE(N__7907),
            .DIN(N__7906),
            .DOUT(N__7905),
            .PACKAGEPIN(TT[0]));
    defparam TT_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_0_preio (
            .PADOEN(N__7907),
            .PADOUT(N__7906),
            .PADIN(N__7905),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_6_iopad (
            .OE(N__7898),
            .DIN(N__7897),
            .DOUT(N__7896),
            .PACKAGEPIN(D[6]));
    defparam D_obuft_6_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_6_preio (
            .PADOEN(N__7898),
            .PADOUT(N__7897),
            .PADIN(N__7896),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3324),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RTC_ENn_obuf_iopad (
            .OE(N__7889),
            .DIN(N__7888),
            .DOUT(N__7887),
            .PACKAGEPIN(RTC_ENn));
    defparam RTC_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RTC_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RTC_ENn_obuf_preio (
            .PADOEN(N__7889),
            .PADOUT(N__7888),
            .PADIN(N__7887),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3253),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_24_iopad (
            .OE(N__7880),
            .DIN(N__7879),
            .DOUT(N__7878),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__7880),
            .PADOUT(N__7879),
            .PADIN(N__7878),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_5_iopad (
            .OE(N__7871),
            .DIN(N__7870),
            .DOUT(N__7869),
            .PACKAGEPIN(D[5]));
    defparam D_obuft_5_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_5_preio (
            .PADOEN(N__7871),
            .PADOUT(N__7870),
            .PADIN(N__7869),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3323),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TM_ibuf_1_iopad (
            .OE(N__7862),
            .DIN(N__7861),
            .DOUT(N__7860),
            .PACKAGEPIN(TM[1]));
    defparam TM_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TM_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TM_ibuf_1_preio (
            .PADOEN(N__7862),
            .PADOUT(N__7861),
            .PADIN(N__7860),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TM_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__7853),
            .DIN(N__7852),
            .DOUT(N__7851),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__7853),
            .PADOUT(N__7852),
            .PADIN(N__7851),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_CIA_obuf_iopad (
            .OE(N__7844),
            .DIN(N__7843),
            .DOUT(N__7842),
            .PACKAGEPIN(CLK_CIA));
    defparam CLK_CIA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_CIA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_CIA_obuf_preio (
            .PADOEN(N__7844),
            .PADOUT(N__7843),
            .PADIN(N__7842),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7183),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_21_iopad (
            .OE(N__7835),
            .DIN(N__7834),
            .DOUT(N__7833),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__7835),
            .PADOUT(N__7834),
            .PADIN(N__7833),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_obuf_iopad (
            .OE(N__7826),
            .DIN(N__7825),
            .DOUT(N__7824),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMSPACEn_obuf_preio (
            .PADOEN(N__7826),
            .PADOUT(N__7825),
            .PADIN(N__7824),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4468),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__7817),
            .DIN(N__7816),
            .DOUT(N__7815),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__7817),
            .PADOUT(N__7816),
            .PADIN(N__7815),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6378),
            .DIN0(TACKn_in),
            .DOUT0(N__4243),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__7808),
            .DIN(N__7807),
            .DOUT(N__7806),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__7808),
            .PADOUT(N__7807),
            .PADIN(N__7806),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ROMENn_obuf_iopad (
            .OE(N__7799),
            .DIN(N__7798),
            .DOUT(N__7797),
            .PACKAGEPIN(ROMENn));
    defparam ROMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ROMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ROMENn_obuf_preio (
            .PADOEN(N__7799),
            .PADOUT(N__7798),
            .PADIN(N__7797),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4123),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuft_iopad (
            .OE(N__7790),
            .DIN(N__7789),
            .DOUT(N__7788),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TBIn_obuft_preio (
            .PADOEN(N__7790),
            .PADOUT(N__7789),
            .PADIN(N__7788),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6382),
            .DIN0(),
            .DOUT0(N__4238),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_0_iopad (
            .OE(N__7781),
            .DIN(N__7780),
            .DOUT(N__7779),
            .PACKAGEPIN(D[0]));
    defparam D_obuft_0_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_0_preio (
            .PADOEN(N__7781),
            .PADOUT(N__7780),
            .PADIN(N__7779),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3308),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_1_iopad (
            .OE(N__7772),
            .DIN(N__7771),
            .DOUT(N__7770),
            .PACKAGEPIN(TT[1]));
    defparam TT_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_1_preio (
            .PADOEN(N__7772),
            .PADOUT(N__7771),
            .PADIN(N__7770),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__7763),
            .DIN(N__7762),
            .DOUT(N__7761),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__7763),
            .PADOUT(N__7762),
            .PADIN(N__7761),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__7754),
            .DIN(N__7753),
            .DOUT(N__7752),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__7754),
            .PADOUT(N__7753),
            .PADIN(N__7752),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5389),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORTSIZE_obuf_iopad (
            .OE(N__7745),
            .DIN(N__7744),
            .DOUT(N__7743),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PORTSIZE_obuf_preio (
            .PADOEN(N__7745),
            .PADOUT(N__7744),
            .PADIN(N__7743),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3751),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_7_iopad (
            .OE(N__7736),
            .DIN(N__7735),
            .DOUT(N__7734),
            .PACKAGEPIN(D[7]));
    defparam D_obuft_7_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_7_preio (
            .PADOEN(N__7736),
            .PADOUT(N__7735),
            .PADIN(N__7734),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3328),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__7727),
            .DIN(N__7726),
            .DOUT(N__7725),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__7727),
            .PADOUT(N__7726),
            .PADIN(N__7725),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_29_iopad (
            .OE(N__7718),
            .DIN(N__7717),
            .DOUT(N__7716),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__7718),
            .PADOUT(N__7717),
            .PADIN(N__7716),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_22_iopad (
            .OE(N__7709),
            .DIN(N__7708),
            .DOUT(N__7707),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__7709),
            .PADOUT(N__7708),
            .PADIN(N__7707),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_27_iopad (
            .OE(N__7700),
            .DIN(N__7699),
            .DOUT(N__7698),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__7700),
            .PADOUT(N__7699),
            .PADIN(N__7698),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__7691),
            .DIN(N__7690),
            .DOUT(N__7689),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__7691),
            .PADOUT(N__7690),
            .PADIN(N__7689),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_2_iopad (
            .OE(N__7682),
            .DIN(N__7681),
            .DOUT(N__7680),
            .PACKAGEPIN(D[2]));
    defparam D_obuft_2_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_2_preio (
            .PADOEN(N__7682),
            .PADOUT(N__7681),
            .PADIN(N__7680),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3275),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__7673),
            .DIN(N__7672),
            .DOUT(N__7671),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__7673),
            .PADOUT(N__7672),
            .PADIN(N__7671),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TM_ibuf_0_iopad (
            .OE(N__7664),
            .DIN(N__7663),
            .DOUT(N__7662),
            .PACKAGEPIN(TM[0]));
    defparam TM_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TM_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TM_ibuf_0_preio (
            .PADOEN(N__7664),
            .PADOUT(N__7663),
            .PADIN(N__7662),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TM_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__7655),
            .DIN(N__7654),
            .DOUT(N__7653),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__7655),
            .PADOUT(N__7654),
            .PADIN(N__7653),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__7646),
            .DIN(N__7645),
            .DOUT(N__7644),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__7646),
            .PADOUT(N__7645),
            .PADIN(N__7644),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_25_iopad (
            .OE(N__7637),
            .DIN(N__7636),
            .DOUT(N__7635),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__7637),
            .PADOUT(N__7636),
            .PADIN(N__7635),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_1_iopad (
            .OE(N__7628),
            .DIN(N__7627),
            .DOUT(N__7626),
            .PACKAGEPIN(D[1]));
    defparam D_obuft_1_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_1_preio (
            .PADOEN(N__7628),
            .PADOUT(N__7627),
            .PADIN(N__7626),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3307),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS0n_obuf_iopad (
            .OE(N__7619),
            .DIN(N__7618),
            .DOUT(N__7617),
            .PACKAGEPIN(CIACS0n));
    defparam CIACS0n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS0n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS0n_obuf_preio (
            .PADOEN(N__7619),
            .PADOUT(N__7618),
            .PADIN(N__7617),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6088),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_4_iopad (
            .OE(N__7610),
            .DIN(N__7609),
            .DOUT(N__7608),
            .PACKAGEPIN(D[4]));
    defparam D_obuft_4_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_4_preio (
            .PADOEN(N__7610),
            .PADOUT(N__7609),
            .PADIN(N__7608),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3322),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK50_obuf_iopad (
            .OE(N__7601),
            .DIN(N__7600),
            .DOUT(N__7599),
            .PACKAGEPIN(TICK50));
    defparam TICK50_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK50_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK50_obuf_preio (
            .PADOEN(N__7601),
            .PADOUT(N__7600),
            .PADIN(N__7599),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7138),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__7592),
            .DIN(N__7591),
            .DOUT(N__7590),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__7592),
            .PADOUT(N__7591),
            .PADIN(N__7590),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_28_iopad (
            .OE(N__7583),
            .DIN(N__7582),
            .DOUT(N__7581),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__7583),
            .PADOUT(N__7582),
            .PADIN(N__7581),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_30_iopad (
            .OE(N__7574),
            .DIN(N__7573),
            .DOUT(N__7572),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__7574),
            .PADOUT(N__7573),
            .PADIN(N__7572),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD OVL_ibuf_iopad (
            .OE(N__7565),
            .DIN(N__7564),
            .DOUT(N__7563),
            .PACKAGEPIN(OVL));
    defparam OVL_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam OVL_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO OVL_ibuf_preio (
            .PADOEN(N__7565),
            .PADOUT(N__7564),
            .PADIN(N__7563),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(OVL_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuft_iopad (
            .OE(N__7556),
            .DIN(N__7555),
            .DOUT(N__7554),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TCIn_obuft_preio (
            .PADOEN(N__7556),
            .PADOUT(N__7555),
            .PADIN(N__7554),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6295),
            .DIN0(),
            .DOUT0(N__4239),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__7547),
            .DIN(N__7546),
            .DOUT(N__7545),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__7547),
            .PADOUT(N__7546),
            .PADIN(N__7545),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__7538),
            .DIN(N__7537),
            .DOUT(N__7536),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__7538),
            .PADOUT(N__7537),
            .PADIN(N__7536),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK60_obuf_iopad (
            .OE(N__7529),
            .DIN(N__7528),
            .DOUT(N__7527),
            .PACKAGEPIN(TICK60));
    defparam TICK60_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK60_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK60_obuf_preio (
            .PADOEN(N__7529),
            .PADOUT(N__7528),
            .PADIN(N__7527),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5662),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_26_iopad (
            .OE(N__7520),
            .DIN(N__7519),
            .DOUT(N__7518),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__7520),
            .PADOUT(N__7519),
            .PADIN(N__7518),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_3_iopad (
            .OE(N__7511),
            .DIN(N__7510),
            .DOUT(N__7509),
            .PACKAGEPIN(D[3]));
    defparam D_obuft_3_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_3_preio (
            .PADOEN(N__7511),
            .PADOUT(N__7510),
            .PADIN(N__7509),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3309),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_23_iopad (
            .OE(N__7502),
            .DIN(N__7501),
            .DOUT(N__7500),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__7502),
            .PADOUT(N__7501),
            .PADIN(N__7500),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_31_iopad (
            .OE(N__7493),
            .DIN(N__7492),
            .DOUT(N__7491),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__7493),
            .PADOUT(N__7492),
            .PADIN(N__7491),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS1n_obuf_iopad (
            .OE(N__7484),
            .DIN(N__7483),
            .DOUT(N__7482),
            .PACKAGEPIN(CIACS1n));
    defparam CIACS1n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS1n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS1n_obuf_preio (
            .PADOEN(N__7484),
            .PADOUT(N__7483),
            .PADIN(N__7482),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6265),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_obuf_iopad (
            .OE(N__7475),
            .DIN(N__7474),
            .DOUT(N__7473),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGSPACEn_obuf_preio (
            .PADOEN(N__7475),
            .PADOUT(N__7474),
            .PADIN(N__7473),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3883),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1767 (
            .O(N__7456),
            .I(N__7451));
    InMux I__1766 (
            .O(N__7455),
            .I(N__7448));
    InMux I__1765 (
            .O(N__7454),
            .I(N__7445));
    LocalMux I__1764 (
            .O(N__7451),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__1763 (
            .O(N__7448),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__1762 (
            .O(N__7445),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    InMux I__1761 (
            .O(N__7438),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ));
    InMux I__1760 (
            .O(N__7435),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ));
    InMux I__1759 (
            .O(N__7432),
            .I(N__7427));
    InMux I__1758 (
            .O(N__7431),
            .I(N__7422));
    InMux I__1757 (
            .O(N__7430),
            .I(N__7422));
    LocalMux I__1756 (
            .O(N__7427),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    LocalMux I__1755 (
            .O(N__7422),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    CascadeMux I__1754 (
            .O(N__7417),
            .I(N__7409));
    InMux I__1753 (
            .O(N__7416),
            .I(N__7406));
    InMux I__1752 (
            .O(N__7415),
            .I(N__7403));
    InMux I__1751 (
            .O(N__7414),
            .I(N__7398));
    InMux I__1750 (
            .O(N__7413),
            .I(N__7398));
    InMux I__1749 (
            .O(N__7412),
            .I(N__7393));
    InMux I__1748 (
            .O(N__7409),
            .I(N__7393));
    LocalMux I__1747 (
            .O(N__7406),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1746 (
            .O(N__7403),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1745 (
            .O(N__7398),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1744 (
            .O(N__7393),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    ClkMux I__1743 (
            .O(N__7384),
            .I(N__7375));
    ClkMux I__1742 (
            .O(N__7383),
            .I(N__7375));
    ClkMux I__1741 (
            .O(N__7382),
            .I(N__7375));
    GlobalMux I__1740 (
            .O(N__7375),
            .I(N__7372));
    gio2CtrlBuf I__1739 (
            .O(N__7372),
            .I(CLK28_IN_c_g));
    InMux I__1738 (
            .O(N__7369),
            .I(N__7366));
    LocalMux I__1737 (
            .O(N__7366),
            .I(\U409_CIA.CIA_CLK_COUNT11_2 ));
    CascadeMux I__1736 (
            .O(N__7363),
            .I(N__7360));
    InMux I__1735 (
            .O(N__7360),
            .I(N__7356));
    InMux I__1734 (
            .O(N__7359),
            .I(N__7353));
    LocalMux I__1733 (
            .O(N__7356),
            .I(\U409_CIA.CIA_CLK_COUNT11_2_0 ));
    LocalMux I__1732 (
            .O(N__7353),
            .I(\U409_CIA.CIA_CLK_COUNT11_2_0 ));
    InMux I__1731 (
            .O(N__7348),
            .I(N__7341));
    InMux I__1730 (
            .O(N__7347),
            .I(N__7341));
    InMux I__1729 (
            .O(N__7346),
            .I(N__7338));
    LocalMux I__1728 (
            .O(N__7341),
            .I(\U409_CIA.CLK_CIA6_4 ));
    LocalMux I__1727 (
            .O(N__7338),
            .I(\U409_CIA.CLK_CIA6_4 ));
    CascadeMux I__1726 (
            .O(N__7333),
            .I(\U409_CIA.CIA_CLK_COUNT11_2_cascade_ ));
    CascadeMux I__1725 (
            .O(N__7330),
            .I(N__7327));
    InMux I__1724 (
            .O(N__7327),
            .I(N__7319));
    InMux I__1723 (
            .O(N__7326),
            .I(N__7314));
    InMux I__1722 (
            .O(N__7325),
            .I(N__7314));
    InMux I__1721 (
            .O(N__7324),
            .I(N__7309));
    InMux I__1720 (
            .O(N__7323),
            .I(N__7309));
    InMux I__1719 (
            .O(N__7322),
            .I(N__7306));
    LocalMux I__1718 (
            .O(N__7319),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1717 (
            .O(N__7314),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1716 (
            .O(N__7309),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1715 (
            .O(N__7306),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    InMux I__1714 (
            .O(N__7297),
            .I(N__7291));
    InMux I__1713 (
            .O(N__7296),
            .I(N__7286));
    InMux I__1712 (
            .O(N__7295),
            .I(N__7286));
    InMux I__1711 (
            .O(N__7294),
            .I(N__7283));
    LocalMux I__1710 (
            .O(N__7291),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1709 (
            .O(N__7286),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1708 (
            .O(N__7283),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    InMux I__1707 (
            .O(N__7276),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ));
    InMux I__1706 (
            .O(N__7273),
            .I(N__7267));
    InMux I__1705 (
            .O(N__7272),
            .I(N__7262));
    InMux I__1704 (
            .O(N__7271),
            .I(N__7262));
    InMux I__1703 (
            .O(N__7270),
            .I(N__7259));
    LocalMux I__1702 (
            .O(N__7267),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__1701 (
            .O(N__7262),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__1700 (
            .O(N__7259),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    InMux I__1699 (
            .O(N__7252),
            .I(N__7249));
    LocalMux I__1698 (
            .O(N__7249),
            .I(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_3 ));
    InMux I__1697 (
            .O(N__7246),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ));
    InMux I__1696 (
            .O(N__7243),
            .I(N__7235));
    InMux I__1695 (
            .O(N__7242),
            .I(N__7235));
    InMux I__1694 (
            .O(N__7241),
            .I(N__7232));
    InMux I__1693 (
            .O(N__7240),
            .I(N__7229));
    LocalMux I__1692 (
            .O(N__7235),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1691 (
            .O(N__7232),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1690 (
            .O(N__7229),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    InMux I__1689 (
            .O(N__7222),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ));
    CascadeMux I__1688 (
            .O(N__7219),
            .I(N__7215));
    CascadeMux I__1687 (
            .O(N__7218),
            .I(N__7210));
    InMux I__1686 (
            .O(N__7215),
            .I(N__7207));
    InMux I__1685 (
            .O(N__7214),
            .I(N__7204));
    InMux I__1684 (
            .O(N__7213),
            .I(N__7199));
    InMux I__1683 (
            .O(N__7210),
            .I(N__7199));
    LocalMux I__1682 (
            .O(N__7207),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1681 (
            .O(N__7204),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1680 (
            .O(N__7199),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    InMux I__1679 (
            .O(N__7192),
            .I(N__7189));
    LocalMux I__1678 (
            .O(N__7189),
            .I(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5 ));
    InMux I__1677 (
            .O(N__7186),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ));
    IoInMux I__1676 (
            .O(N__7183),
            .I(N__7180));
    LocalMux I__1675 (
            .O(N__7180),
            .I(N__7177));
    Span4Mux_s3_v I__1674 (
            .O(N__7177),
            .I(N__7174));
    Span4Mux_v I__1673 (
            .O(N__7174),
            .I(N__7171));
    Span4Mux_v I__1672 (
            .O(N__7171),
            .I(N__7167));
    CascadeMux I__1671 (
            .O(N__7170),
            .I(N__7162));
    Span4Mux_v I__1670 (
            .O(N__7167),
            .I(N__7159));
    InMux I__1669 (
            .O(N__7166),
            .I(N__7156));
    InMux I__1668 (
            .O(N__7165),
            .I(N__7151));
    InMux I__1667 (
            .O(N__7162),
            .I(N__7151));
    Odrv4 I__1666 (
            .O(N__7159),
            .I(CLK_CIA_c));
    LocalMux I__1665 (
            .O(N__7156),
            .I(CLK_CIA_c));
    LocalMux I__1664 (
            .O(N__7151),
            .I(CLK_CIA_c));
    InMux I__1663 (
            .O(N__7144),
            .I(N__7141));
    LocalMux I__1662 (
            .O(N__7141),
            .I(\U409_CIA.CLK_CIA_r_1_0 ));
    IoInMux I__1661 (
            .O(N__7138),
            .I(N__7135));
    LocalMux I__1660 (
            .O(N__7135),
            .I(N__7132));
    Span4Mux_s3_v I__1659 (
            .O(N__7132),
            .I(N__7129));
    Span4Mux_v I__1658 (
            .O(N__7129),
            .I(N__7126));
    Span4Mux_v I__1657 (
            .O(N__7126),
            .I(N__7123));
    Span4Mux_h I__1656 (
            .O(N__7123),
            .I(N__7119));
    InMux I__1655 (
            .O(N__7122),
            .I(N__7116));
    Odrv4 I__1654 (
            .O(N__7119),
            .I(TICK50_c));
    LocalMux I__1653 (
            .O(N__7116),
            .I(TICK50_c));
    CascadeMux I__1652 (
            .O(N__7111),
            .I(N__7108));
    InMux I__1651 (
            .O(N__7108),
            .I(N__7105));
    LocalMux I__1650 (
            .O(N__7105),
            .I(N__7102));
    Span4Mux_h I__1649 (
            .O(N__7102),
            .I(N__7099));
    Odrv4 I__1648 (
            .O(N__7099),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ));
    CascadeMux I__1647 (
            .O(N__7096),
            .I(N__7093));
    InMux I__1646 (
            .O(N__7093),
            .I(N__7089));
    InMux I__1645 (
            .O(N__7092),
            .I(N__7086));
    LocalMux I__1644 (
            .O(N__7089),
            .I(N__7083));
    LocalMux I__1643 (
            .O(N__7086),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    Odrv4 I__1642 (
            .O(N__7083),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    InMux I__1641 (
            .O(N__7078),
            .I(N__7075));
    LocalMux I__1640 (
            .O(N__7075),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ));
    InMux I__1639 (
            .O(N__7072),
            .I(N__7068));
    InMux I__1638 (
            .O(N__7071),
            .I(N__7065));
    LocalMux I__1637 (
            .O(N__7068),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    LocalMux I__1636 (
            .O(N__7065),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    InMux I__1635 (
            .O(N__7060),
            .I(N__7056));
    InMux I__1634 (
            .O(N__7059),
            .I(N__7053));
    LocalMux I__1633 (
            .O(N__7056),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    LocalMux I__1632 (
            .O(N__7053),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    CascadeMux I__1631 (
            .O(N__7048),
            .I(N__7045));
    InMux I__1630 (
            .O(N__7045),
            .I(N__7041));
    InMux I__1629 (
            .O(N__7044),
            .I(N__7038));
    LocalMux I__1628 (
            .O(N__7041),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    LocalMux I__1627 (
            .O(N__7038),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    CascadeMux I__1626 (
            .O(N__7033),
            .I(N__7027));
    CascadeMux I__1625 (
            .O(N__7032),
            .I(N__7024));
    CascadeMux I__1624 (
            .O(N__7031),
            .I(N__7020));
    CascadeMux I__1623 (
            .O(N__7030),
            .I(N__7015));
    InMux I__1622 (
            .O(N__7027),
            .I(N__7011));
    InMux I__1621 (
            .O(N__7024),
            .I(N__7008));
    InMux I__1620 (
            .O(N__7023),
            .I(N__7003));
    InMux I__1619 (
            .O(N__7020),
            .I(N__7003));
    InMux I__1618 (
            .O(N__7019),
            .I(N__6994));
    InMux I__1617 (
            .O(N__7018),
            .I(N__6994));
    InMux I__1616 (
            .O(N__7015),
            .I(N__6994));
    InMux I__1615 (
            .O(N__7014),
            .I(N__6994));
    LocalMux I__1614 (
            .O(N__7011),
            .I(N__6991));
    LocalMux I__1613 (
            .O(N__7008),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__1612 (
            .O(N__7003),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__1611 (
            .O(N__6994),
            .I(\U409_TICK.TICK503_10 ));
    Odrv4 I__1610 (
            .O(N__6991),
            .I(\U409_TICK.TICK503_10 ));
    InMux I__1609 (
            .O(N__6982),
            .I(N__6972));
    InMux I__1608 (
            .O(N__6981),
            .I(N__6967));
    InMux I__1607 (
            .O(N__6980),
            .I(N__6967));
    InMux I__1606 (
            .O(N__6979),
            .I(N__6962));
    InMux I__1605 (
            .O(N__6978),
            .I(N__6962));
    InMux I__1604 (
            .O(N__6977),
            .I(N__6955));
    InMux I__1603 (
            .O(N__6976),
            .I(N__6955));
    InMux I__1602 (
            .O(N__6975),
            .I(N__6955));
    LocalMux I__1601 (
            .O(N__6972),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__1600 (
            .O(N__6967),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__1599 (
            .O(N__6962),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__1598 (
            .O(N__6955),
            .I(\U409_TICK.TICK503_9 ));
    InMux I__1597 (
            .O(N__6946),
            .I(N__6932));
    InMux I__1596 (
            .O(N__6945),
            .I(N__6932));
    InMux I__1595 (
            .O(N__6944),
            .I(N__6932));
    InMux I__1594 (
            .O(N__6943),
            .I(N__6927));
    InMux I__1593 (
            .O(N__6942),
            .I(N__6927));
    InMux I__1592 (
            .O(N__6941),
            .I(N__6924));
    InMux I__1591 (
            .O(N__6940),
            .I(N__6919));
    InMux I__1590 (
            .O(N__6939),
            .I(N__6919));
    LocalMux I__1589 (
            .O(N__6932),
            .I(N__6916));
    LocalMux I__1588 (
            .O(N__6927),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__1587 (
            .O(N__6924),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__1586 (
            .O(N__6919),
            .I(\U409_TICK.TICK503_14 ));
    Odrv4 I__1585 (
            .O(N__6916),
            .I(\U409_TICK.TICK503_14 ));
    CascadeMux I__1584 (
            .O(N__6907),
            .I(\U409_TICK.TICK503_10_cascade_ ));
    InMux I__1583 (
            .O(N__6904),
            .I(N__6901));
    LocalMux I__1582 (
            .O(N__6901),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ));
    InMux I__1581 (
            .O(N__6898),
            .I(N__6894));
    InMux I__1580 (
            .O(N__6897),
            .I(N__6891));
    LocalMux I__1579 (
            .O(N__6894),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    LocalMux I__1578 (
            .O(N__6891),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    ClkMux I__1577 (
            .O(N__6886),
            .I(N__6853));
    ClkMux I__1576 (
            .O(N__6885),
            .I(N__6853));
    ClkMux I__1575 (
            .O(N__6884),
            .I(N__6853));
    ClkMux I__1574 (
            .O(N__6883),
            .I(N__6853));
    ClkMux I__1573 (
            .O(N__6882),
            .I(N__6853));
    ClkMux I__1572 (
            .O(N__6881),
            .I(N__6853));
    ClkMux I__1571 (
            .O(N__6880),
            .I(N__6853));
    ClkMux I__1570 (
            .O(N__6879),
            .I(N__6853));
    ClkMux I__1569 (
            .O(N__6878),
            .I(N__6853));
    ClkMux I__1568 (
            .O(N__6877),
            .I(N__6853));
    ClkMux I__1567 (
            .O(N__6876),
            .I(N__6853));
    GlobalMux I__1566 (
            .O(N__6853),
            .I(N__6850));
    gio2CtrlBuf I__1565 (
            .O(N__6850),
            .I(CLK6_c_g));
    InMux I__1564 (
            .O(N__6847),
            .I(\U409_TICK.un2_COUNTER50_1_cry_12 ));
    InMux I__1563 (
            .O(N__6844),
            .I(\U409_TICK.un2_COUNTER50_1_cry_13 ));
    InMux I__1562 (
            .O(N__6841),
            .I(\U409_TICK.un2_COUNTER50_1_cry_14 ));
    InMux I__1561 (
            .O(N__6838),
            .I(\U409_TICK.un2_COUNTER50_1_cry_15 ));
    InMux I__1560 (
            .O(N__6835),
            .I(N__6831));
    InMux I__1559 (
            .O(N__6834),
            .I(N__6828));
    LocalMux I__1558 (
            .O(N__6831),
            .I(N__6825));
    LocalMux I__1557 (
            .O(N__6828),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    Odrv4 I__1556 (
            .O(N__6825),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    CascadeMux I__1555 (
            .O(N__6820),
            .I(\U409_CIA.CLK_CIA6_3_cascade_ ));
    CascadeMux I__1554 (
            .O(N__6817),
            .I(\U409_CIA.un1_CIA_CLK_COUNT_3_2_cascade_ ));
    InMux I__1553 (
            .O(N__6814),
            .I(N__6811));
    LocalMux I__1552 (
            .O(N__6811),
            .I(N__6807));
    InMux I__1551 (
            .O(N__6810),
            .I(N__6804));
    Span4Mux_v I__1550 (
            .O(N__6807),
            .I(N__6800));
    LocalMux I__1549 (
            .O(N__6804),
            .I(N__6797));
    InMux I__1548 (
            .O(N__6803),
            .I(N__6794));
    Span4Mux_h I__1547 (
            .O(N__6800),
            .I(N__6791));
    Span12Mux_h I__1546 (
            .O(N__6797),
            .I(N__6788));
    LocalMux I__1545 (
            .O(N__6794),
            .I(N__6785));
    Odrv4 I__1544 (
            .O(N__6791),
            .I(CIA_SPACE));
    Odrv12 I__1543 (
            .O(N__6788),
            .I(CIA_SPACE));
    Odrv4 I__1542 (
            .O(N__6785),
            .I(CIA_SPACE));
    CascadeMux I__1541 (
            .O(N__6778),
            .I(\U409_CIA.VMA_RNOZ0Z_0_cascade_ ));
    InMux I__1540 (
            .O(N__6775),
            .I(N__6771));
    InMux I__1539 (
            .O(N__6774),
            .I(N__6768));
    LocalMux I__1538 (
            .O(N__6771),
            .I(N__6765));
    LocalMux I__1537 (
            .O(N__6768),
            .I(N__6761));
    Span4Mux_v I__1536 (
            .O(N__6765),
            .I(N__6758));
    InMux I__1535 (
            .O(N__6764),
            .I(N__6755));
    Odrv12 I__1534 (
            .O(N__6761),
            .I(\U409_CIA.VMAZ0 ));
    Odrv4 I__1533 (
            .O(N__6758),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__1532 (
            .O(N__6755),
            .I(\U409_CIA.VMAZ0 ));
    InMux I__1531 (
            .O(N__6748),
            .I(N__6744));
    InMux I__1530 (
            .O(N__6747),
            .I(N__6741));
    LocalMux I__1529 (
            .O(N__6744),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    LocalMux I__1528 (
            .O(N__6741),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    InMux I__1527 (
            .O(N__6736),
            .I(N__6733));
    LocalMux I__1526 (
            .O(N__6733),
            .I(N__6730));
    Odrv4 I__1525 (
            .O(N__6730),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ));
    InMux I__1524 (
            .O(N__6727),
            .I(\U409_TICK.un2_COUNTER50_1_cry_4 ));
    InMux I__1523 (
            .O(N__6724),
            .I(N__6720));
    InMux I__1522 (
            .O(N__6723),
            .I(N__6717));
    LocalMux I__1521 (
            .O(N__6720),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    LocalMux I__1520 (
            .O(N__6717),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    CascadeMux I__1519 (
            .O(N__6712),
            .I(N__6709));
    InMux I__1518 (
            .O(N__6709),
            .I(N__6706));
    LocalMux I__1517 (
            .O(N__6706),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ));
    InMux I__1516 (
            .O(N__6703),
            .I(\U409_TICK.un2_COUNTER50_1_cry_5 ));
    InMux I__1515 (
            .O(N__6700),
            .I(\U409_TICK.un2_COUNTER50_1_cry_6 ));
    CascadeMux I__1514 (
            .O(N__6697),
            .I(N__6694));
    InMux I__1513 (
            .O(N__6694),
            .I(N__6690));
    InMux I__1512 (
            .O(N__6693),
            .I(N__6687));
    LocalMux I__1511 (
            .O(N__6690),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    LocalMux I__1510 (
            .O(N__6687),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    InMux I__1509 (
            .O(N__6682),
            .I(\U409_TICK.un2_COUNTER50_1_cry_7 ));
    CascadeMux I__1508 (
            .O(N__6679),
            .I(N__6675));
    InMux I__1507 (
            .O(N__6678),
            .I(N__6672));
    InMux I__1506 (
            .O(N__6675),
            .I(N__6669));
    LocalMux I__1505 (
            .O(N__6672),
            .I(N__6666));
    LocalMux I__1504 (
            .O(N__6669),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    Odrv4 I__1503 (
            .O(N__6666),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    InMux I__1502 (
            .O(N__6661),
            .I(N__6658));
    LocalMux I__1501 (
            .O(N__6658),
            .I(N__6655));
    Odrv4 I__1500 (
            .O(N__6655),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ));
    InMux I__1499 (
            .O(N__6652),
            .I(bfn_14_10_0_));
    InMux I__1498 (
            .O(N__6649),
            .I(N__6646));
    LocalMux I__1497 (
            .O(N__6646),
            .I(N__6642));
    InMux I__1496 (
            .O(N__6645),
            .I(N__6639));
    Odrv4 I__1495 (
            .O(N__6642),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    LocalMux I__1494 (
            .O(N__6639),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    InMux I__1493 (
            .O(N__6634),
            .I(\U409_TICK.un2_COUNTER50_1_cry_9 ));
    InMux I__1492 (
            .O(N__6631),
            .I(N__6627));
    InMux I__1491 (
            .O(N__6630),
            .I(N__6624));
    LocalMux I__1490 (
            .O(N__6627),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    LocalMux I__1489 (
            .O(N__6624),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    InMux I__1488 (
            .O(N__6619),
            .I(N__6616));
    LocalMux I__1487 (
            .O(N__6616),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ));
    InMux I__1486 (
            .O(N__6613),
            .I(\U409_TICK.un2_COUNTER50_1_cry_10 ));
    InMux I__1485 (
            .O(N__6610),
            .I(N__6607));
    LocalMux I__1484 (
            .O(N__6607),
            .I(N__6603));
    InMux I__1483 (
            .O(N__6606),
            .I(N__6600));
    Odrv4 I__1482 (
            .O(N__6603),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    LocalMux I__1481 (
            .O(N__6600),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    InMux I__1480 (
            .O(N__6595),
            .I(\U409_TICK.un2_COUNTER50_1_cry_11 ));
    CascadeMux I__1479 (
            .O(N__6592),
            .I(\U409_TICK.TICK503_14_cascade_ ));
    InMux I__1478 (
            .O(N__6589),
            .I(N__6586));
    LocalMux I__1477 (
            .O(N__6586),
            .I(\U409_TICK.TICK503_8 ));
    CascadeMux I__1476 (
            .O(N__6583),
            .I(\U409_TICK.TICK503_9_cascade_ ));
    InMux I__1475 (
            .O(N__6580),
            .I(N__6574));
    InMux I__1474 (
            .O(N__6579),
            .I(N__6569));
    InMux I__1473 (
            .O(N__6578),
            .I(N__6569));
    InMux I__1472 (
            .O(N__6577),
            .I(N__6566));
    LocalMux I__1471 (
            .O(N__6574),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__1470 (
            .O(N__6569),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__1469 (
            .O(N__6566),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    CascadeMux I__1468 (
            .O(N__6559),
            .I(N__6554));
    InMux I__1467 (
            .O(N__6558),
            .I(N__6551));
    InMux I__1466 (
            .O(N__6557),
            .I(N__6548));
    InMux I__1465 (
            .O(N__6554),
            .I(N__6545));
    LocalMux I__1464 (
            .O(N__6551),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__1463 (
            .O(N__6548),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__1462 (
            .O(N__6545),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    InMux I__1461 (
            .O(N__6538),
            .I(N__6534));
    InMux I__1460 (
            .O(N__6537),
            .I(N__6531));
    LocalMux I__1459 (
            .O(N__6534),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    LocalMux I__1458 (
            .O(N__6531),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    InMux I__1457 (
            .O(N__6526),
            .I(\U409_TICK.un2_COUNTER50_1_cry_1 ));
    InMux I__1456 (
            .O(N__6523),
            .I(N__6519));
    InMux I__1455 (
            .O(N__6522),
            .I(N__6516));
    LocalMux I__1454 (
            .O(N__6519),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    LocalMux I__1453 (
            .O(N__6516),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    InMux I__1452 (
            .O(N__6511),
            .I(\U409_TICK.un2_COUNTER50_1_cry_2 ));
    InMux I__1451 (
            .O(N__6508),
            .I(\U409_TICK.un2_COUNTER50_1_cry_3 ));
    InMux I__1450 (
            .O(N__6505),
            .I(N__6502));
    LocalMux I__1449 (
            .O(N__6502),
            .I(N__6496));
    InMux I__1448 (
            .O(N__6501),
            .I(N__6491));
    InMux I__1447 (
            .O(N__6500),
            .I(N__6491));
    InMux I__1446 (
            .O(N__6499),
            .I(N__6488));
    Span4Mux_h I__1445 (
            .O(N__6496),
            .I(N__6485));
    LocalMux I__1444 (
            .O(N__6491),
            .I(N__6482));
    LocalMux I__1443 (
            .O(N__6488),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    Odrv4 I__1442 (
            .O(N__6485),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    Odrv4 I__1441 (
            .O(N__6482),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    InMux I__1440 (
            .O(N__6475),
            .I(N__6472));
    LocalMux I__1439 (
            .O(N__6472),
            .I(N__6467));
    InMux I__1438 (
            .O(N__6471),
            .I(N__6462));
    InMux I__1437 (
            .O(N__6470),
            .I(N__6462));
    Span4Mux_h I__1436 (
            .O(N__6467),
            .I(N__6459));
    LocalMux I__1435 (
            .O(N__6462),
            .I(N__6456));
    Odrv4 I__1434 (
            .O(N__6459),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    Odrv12 I__1433 (
            .O(N__6456),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    SRMux I__1432 (
            .O(N__6451),
            .I(N__6447));
    SRMux I__1431 (
            .O(N__6450),
            .I(N__6443));
    LocalMux I__1430 (
            .O(N__6447),
            .I(N__6438));
    SRMux I__1429 (
            .O(N__6446),
            .I(N__6435));
    LocalMux I__1428 (
            .O(N__6443),
            .I(N__6431));
    SRMux I__1427 (
            .O(N__6442),
            .I(N__6428));
    SRMux I__1426 (
            .O(N__6441),
            .I(N__6425));
    Span4Mux_v I__1425 (
            .O(N__6438),
            .I(N__6420));
    LocalMux I__1424 (
            .O(N__6435),
            .I(N__6420));
    SRMux I__1423 (
            .O(N__6434),
            .I(N__6417));
    Span4Mux_h I__1422 (
            .O(N__6431),
            .I(N__6412));
    LocalMux I__1421 (
            .O(N__6428),
            .I(N__6412));
    LocalMux I__1420 (
            .O(N__6425),
            .I(N__6409));
    Span4Mux_v I__1419 (
            .O(N__6420),
            .I(N__6403));
    LocalMux I__1418 (
            .O(N__6417),
            .I(N__6403));
    Span4Mux_v I__1417 (
            .O(N__6412),
            .I(N__6400));
    Span4Mux_h I__1416 (
            .O(N__6409),
            .I(N__6397));
    InMux I__1415 (
            .O(N__6408),
            .I(N__6394));
    Span4Mux_v I__1414 (
            .O(N__6403),
            .I(N__6391));
    Odrv4 I__1413 (
            .O(N__6400),
            .I(RESETn_c_i));
    Odrv4 I__1412 (
            .O(N__6397),
            .I(RESETn_c_i));
    LocalMux I__1411 (
            .O(N__6394),
            .I(RESETn_c_i));
    Odrv4 I__1410 (
            .O(N__6391),
            .I(RESETn_c_i));
    IoInMux I__1409 (
            .O(N__6382),
            .I(N__6379));
    LocalMux I__1408 (
            .O(N__6379),
            .I(N__6375));
    IoInMux I__1407 (
            .O(N__6378),
            .I(N__6372));
    IoSpan4Mux I__1406 (
            .O(N__6375),
            .I(N__6367));
    LocalMux I__1405 (
            .O(N__6372),
            .I(N__6367));
    IoSpan4Mux I__1404 (
            .O(N__6367),
            .I(N__6364));
    Span4Mux_s2_v I__1403 (
            .O(N__6364),
            .I(N__6361));
    Sp12to4 I__1402 (
            .O(N__6361),
            .I(N__6357));
    InMux I__1401 (
            .O(N__6360),
            .I(N__6354));
    Span12Mux_s10_v I__1400 (
            .O(N__6357),
            .I(N__6348));
    LocalMux I__1399 (
            .O(N__6354),
            .I(N__6348));
    CascadeMux I__1398 (
            .O(N__6353),
            .I(N__6345));
    Span12Mux_h I__1397 (
            .O(N__6348),
            .I(N__6342));
    InMux I__1396 (
            .O(N__6345),
            .I(N__6339));
    Odrv12 I__1395 (
            .O(N__6342),
            .I(TACK_EN));
    LocalMux I__1394 (
            .O(N__6339),
            .I(TACK_EN));
    InMux I__1393 (
            .O(N__6334),
            .I(N__6330));
    InMux I__1392 (
            .O(N__6333),
            .I(N__6327));
    LocalMux I__1391 (
            .O(N__6330),
            .I(N__6323));
    LocalMux I__1390 (
            .O(N__6327),
            .I(N__6320));
    InMux I__1389 (
            .O(N__6326),
            .I(N__6317));
    Span4Mux_v I__1388 (
            .O(N__6323),
            .I(N__6314));
    Span4Mux_v I__1387 (
            .O(N__6320),
            .I(N__6311));
    LocalMux I__1386 (
            .O(N__6317),
            .I(N__6308));
    Sp12to4 I__1385 (
            .O(N__6314),
            .I(N__6305));
    Span4Mux_h I__1384 (
            .O(N__6311),
            .I(N__6300));
    Span4Mux_v I__1383 (
            .O(N__6308),
            .I(N__6300));
    Odrv12 I__1382 (
            .O(N__6305),
            .I(AUTOCONFIG_SPACE));
    Odrv4 I__1381 (
            .O(N__6300),
            .I(AUTOCONFIG_SPACE));
    IoInMux I__1380 (
            .O(N__6295),
            .I(N__6292));
    LocalMux I__1379 (
            .O(N__6292),
            .I(N__6289));
    Span12Mux_s1_v I__1378 (
            .O(N__6289),
            .I(N__6286));
    Span12Mux_h I__1377 (
            .O(N__6286),
            .I(N__6283));
    Odrv12 I__1376 (
            .O(N__6283),
            .I(TCIn_1_i));
    InMux I__1375 (
            .O(N__6280),
            .I(N__6277));
    LocalMux I__1374 (
            .O(N__6277),
            .I(N__6274));
    Span12Mux_v I__1373 (
            .O(N__6274),
            .I(N__6271));
    Span12Mux_h I__1372 (
            .O(N__6271),
            .I(N__6268));
    Odrv12 I__1371 (
            .O(N__6268),
            .I(A_c_13));
    IoInMux I__1370 (
            .O(N__6265),
            .I(N__6262));
    LocalMux I__1369 (
            .O(N__6262),
            .I(N__6259));
    Span4Mux_s2_h I__1368 (
            .O(N__6259),
            .I(N__6256));
    Span4Mux_h I__1367 (
            .O(N__6256),
            .I(N__6253));
    Sp12to4 I__1366 (
            .O(N__6253),
            .I(N__6250));
    Span12Mux_s9_v I__1365 (
            .O(N__6250),
            .I(N__6247));
    Odrv12 I__1364 (
            .O(N__6247),
            .I(U409_ADDRESS_DECODE_un1_CIACS1n_i));
    InMux I__1363 (
            .O(N__6244),
            .I(N__6239));
    InMux I__1362 (
            .O(N__6243),
            .I(N__6236));
    InMux I__1361 (
            .O(N__6242),
            .I(N__6233));
    LocalMux I__1360 (
            .O(N__6239),
            .I(N__6227));
    LocalMux I__1359 (
            .O(N__6236),
            .I(N__6227));
    LocalMux I__1358 (
            .O(N__6233),
            .I(N__6222));
    CascadeMux I__1357 (
            .O(N__6232),
            .I(N__6219));
    Span4Mux_v I__1356 (
            .O(N__6227),
            .I(N__6216));
    InMux I__1355 (
            .O(N__6226),
            .I(N__6213));
    CascadeMux I__1354 (
            .O(N__6225),
            .I(N__6209));
    Span4Mux_v I__1353 (
            .O(N__6222),
            .I(N__6204));
    InMux I__1352 (
            .O(N__6219),
            .I(N__6201));
    Span4Mux_h I__1351 (
            .O(N__6216),
            .I(N__6196));
    LocalMux I__1350 (
            .O(N__6213),
            .I(N__6196));
    InMux I__1349 (
            .O(N__6212),
            .I(N__6189));
    InMux I__1348 (
            .O(N__6209),
            .I(N__6189));
    InMux I__1347 (
            .O(N__6208),
            .I(N__6189));
    InMux I__1346 (
            .O(N__6207),
            .I(N__6182));
    Span4Mux_h I__1345 (
            .O(N__6204),
            .I(N__6179));
    LocalMux I__1344 (
            .O(N__6201),
            .I(N__6176));
    Span4Mux_v I__1343 (
            .O(N__6196),
            .I(N__6171));
    LocalMux I__1342 (
            .O(N__6189),
            .I(N__6171));
    InMux I__1341 (
            .O(N__6188),
            .I(N__6168));
    InMux I__1340 (
            .O(N__6187),
            .I(N__6165));
    InMux I__1339 (
            .O(N__6186),
            .I(N__6162));
    InMux I__1338 (
            .O(N__6185),
            .I(N__6159));
    LocalMux I__1337 (
            .O(N__6182),
            .I(N__6156));
    Span4Mux_h I__1336 (
            .O(N__6179),
            .I(N__6151));
    Span4Mux_v I__1335 (
            .O(N__6176),
            .I(N__6151));
    Span4Mux_h I__1334 (
            .O(N__6171),
            .I(N__6142));
    LocalMux I__1333 (
            .O(N__6168),
            .I(N__6142));
    LocalMux I__1332 (
            .O(N__6165),
            .I(N__6142));
    LocalMux I__1331 (
            .O(N__6162),
            .I(N__6142));
    LocalMux I__1330 (
            .O(N__6159),
            .I(N__6139));
    Span12Mux_h I__1329 (
            .O(N__6156),
            .I(N__6134));
    Sp12to4 I__1328 (
            .O(N__6151),
            .I(N__6134));
    Span4Mux_v I__1327 (
            .O(N__6142),
            .I(N__6131));
    Span4Mux_v I__1326 (
            .O(N__6139),
            .I(N__6128));
    Span12Mux_v I__1325 (
            .O(N__6134),
            .I(N__6121));
    Sp12to4 I__1324 (
            .O(N__6131),
            .I(N__6121));
    Sp12to4 I__1323 (
            .O(N__6128),
            .I(N__6121));
    Span12Mux_h I__1322 (
            .O(N__6121),
            .I(N__6118));
    Odrv12 I__1321 (
            .O(N__6118),
            .I(RESETn_c));
    InMux I__1320 (
            .O(N__6115),
            .I(N__6112));
    LocalMux I__1319 (
            .O(N__6112),
            .I(CIA_ENABLE));
    InMux I__1318 (
            .O(N__6109),
            .I(N__6106));
    LocalMux I__1317 (
            .O(N__6106),
            .I(N__6103));
    Span4Mux_v I__1316 (
            .O(N__6103),
            .I(N__6100));
    Sp12to4 I__1315 (
            .O(N__6100),
            .I(N__6097));
    Span12Mux_h I__1314 (
            .O(N__6097),
            .I(N__6094));
    Odrv12 I__1313 (
            .O(N__6094),
            .I(A_c_12));
    CascadeMux I__1312 (
            .O(N__6091),
            .I(CIA_ENABLE_cascade_));
    IoInMux I__1311 (
            .O(N__6088),
            .I(N__6085));
    LocalMux I__1310 (
            .O(N__6085),
            .I(N__6082));
    IoSpan4Mux I__1309 (
            .O(N__6082),
            .I(N__6079));
    Sp12to4 I__1308 (
            .O(N__6079),
            .I(N__6076));
    Span12Mux_s7_v I__1307 (
            .O(N__6076),
            .I(N__6073));
    Span12Mux_h I__1306 (
            .O(N__6073),
            .I(N__6070));
    Odrv12 I__1305 (
            .O(N__6070),
            .I(U409_ADDRESS_DECODE_un1_CIACS0n_i));
    CascadeMux I__1304 (
            .O(N__6067),
            .I(\U409_TICK.TICK503_11_cascade_ ));
    InMux I__1303 (
            .O(N__6064),
            .I(N__6060));
    InMux I__1302 (
            .O(N__6063),
            .I(N__6057));
    LocalMux I__1301 (
            .O(N__6060),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    LocalMux I__1300 (
            .O(N__6057),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    InMux I__1299 (
            .O(N__6052),
            .I(N__6048));
    InMux I__1298 (
            .O(N__6051),
            .I(N__6045));
    LocalMux I__1297 (
            .O(N__6048),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    LocalMux I__1296 (
            .O(N__6045),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    CascadeMux I__1295 (
            .O(N__6040),
            .I(N__6035));
    CascadeMux I__1294 (
            .O(N__6039),
            .I(N__6032));
    InMux I__1293 (
            .O(N__6038),
            .I(N__6029));
    InMux I__1292 (
            .O(N__6035),
            .I(N__6026));
    InMux I__1291 (
            .O(N__6032),
            .I(N__6023));
    LocalMux I__1290 (
            .O(N__6029),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__1289 (
            .O(N__6026),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__1288 (
            .O(N__6023),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    InMux I__1287 (
            .O(N__6016),
            .I(N__6012));
    InMux I__1286 (
            .O(N__6015),
            .I(N__6009));
    LocalMux I__1285 (
            .O(N__6012),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    LocalMux I__1284 (
            .O(N__6009),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    InMux I__1283 (
            .O(N__6004),
            .I(N__6000));
    InMux I__1282 (
            .O(N__6003),
            .I(N__5997));
    LocalMux I__1281 (
            .O(N__6000),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    LocalMux I__1280 (
            .O(N__5997),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    InMux I__1279 (
            .O(N__5992),
            .I(N__5989));
    LocalMux I__1278 (
            .O(N__5989),
            .I(\U409_TICK.TICK603_8 ));
    CascadeMux I__1277 (
            .O(N__5986),
            .I(\U409_TICK.TICK603_11_cascade_ ));
    InMux I__1276 (
            .O(N__5983),
            .I(N__5979));
    InMux I__1275 (
            .O(N__5982),
            .I(N__5976));
    LocalMux I__1274 (
            .O(N__5979),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    LocalMux I__1273 (
            .O(N__5976),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    CascadeMux I__1272 (
            .O(N__5971),
            .I(\U409_TICK.TICK603_14_cascade_ ));
    InMux I__1271 (
            .O(N__5968),
            .I(N__5965));
    LocalMux I__1270 (
            .O(N__5965),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ));
    InMux I__1269 (
            .O(N__5962),
            .I(N__5958));
    InMux I__1268 (
            .O(N__5961),
            .I(N__5955));
    LocalMux I__1267 (
            .O(N__5958),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    LocalMux I__1266 (
            .O(N__5955),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    InMux I__1265 (
            .O(N__5950),
            .I(N__5946));
    InMux I__1264 (
            .O(N__5949),
            .I(N__5943));
    LocalMux I__1263 (
            .O(N__5946),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    LocalMux I__1262 (
            .O(N__5943),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    CascadeMux I__1261 (
            .O(N__5938),
            .I(N__5935));
    InMux I__1260 (
            .O(N__5935),
            .I(N__5931));
    InMux I__1259 (
            .O(N__5934),
            .I(N__5928));
    LocalMux I__1258 (
            .O(N__5931),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    LocalMux I__1257 (
            .O(N__5928),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    CascadeMux I__1256 (
            .O(N__5923),
            .I(\U409_TICK.TICK603_9_cascade_ ));
    InMux I__1255 (
            .O(N__5920),
            .I(N__5917));
    LocalMux I__1254 (
            .O(N__5917),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ));
    InMux I__1253 (
            .O(N__5914),
            .I(N__5910));
    InMux I__1252 (
            .O(N__5913),
            .I(N__5907));
    LocalMux I__1251 (
            .O(N__5910),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    LocalMux I__1250 (
            .O(N__5907),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    InMux I__1249 (
            .O(N__5902),
            .I(N__5898));
    InMux I__1248 (
            .O(N__5901),
            .I(N__5895));
    LocalMux I__1247 (
            .O(N__5898),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    LocalMux I__1246 (
            .O(N__5895),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    InMux I__1245 (
            .O(N__5890),
            .I(N__5886));
    InMux I__1244 (
            .O(N__5889),
            .I(N__5883));
    LocalMux I__1243 (
            .O(N__5886),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    LocalMux I__1242 (
            .O(N__5883),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    CascadeMux I__1241 (
            .O(N__5878),
            .I(N__5875));
    InMux I__1240 (
            .O(N__5875),
            .I(N__5871));
    InMux I__1239 (
            .O(N__5874),
            .I(N__5868));
    LocalMux I__1238 (
            .O(N__5871),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    LocalMux I__1237 (
            .O(N__5868),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    CascadeMux I__1236 (
            .O(N__5863),
            .I(\U409_TICK.TICK603_10_cascade_ ));
    InMux I__1235 (
            .O(N__5860),
            .I(N__5857));
    LocalMux I__1234 (
            .O(N__5857),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ));
    InMux I__1233 (
            .O(N__5854),
            .I(N__5850));
    InMux I__1232 (
            .O(N__5853),
            .I(N__5847));
    LocalMux I__1231 (
            .O(N__5850),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    LocalMux I__1230 (
            .O(N__5847),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    InMux I__1229 (
            .O(N__5842),
            .I(N__5833));
    InMux I__1228 (
            .O(N__5841),
            .I(N__5828));
    InMux I__1227 (
            .O(N__5840),
            .I(N__5828));
    InMux I__1226 (
            .O(N__5839),
            .I(N__5823));
    InMux I__1225 (
            .O(N__5838),
            .I(N__5823));
    InMux I__1224 (
            .O(N__5837),
            .I(N__5818));
    InMux I__1223 (
            .O(N__5836),
            .I(N__5818));
    LocalMux I__1222 (
            .O(N__5833),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__1221 (
            .O(N__5828),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__1220 (
            .O(N__5823),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__1219 (
            .O(N__5818),
            .I(\U409_TICK.TICK603_9 ));
    CascadeMux I__1218 (
            .O(N__5809),
            .I(N__5805));
    CascadeMux I__1217 (
            .O(N__5808),
            .I(N__5802));
    InMux I__1216 (
            .O(N__5805),
            .I(N__5794));
    InMux I__1215 (
            .O(N__5802),
            .I(N__5789));
    InMux I__1214 (
            .O(N__5801),
            .I(N__5789));
    InMux I__1213 (
            .O(N__5800),
            .I(N__5784));
    InMux I__1212 (
            .O(N__5799),
            .I(N__5784));
    InMux I__1211 (
            .O(N__5798),
            .I(N__5779));
    InMux I__1210 (
            .O(N__5797),
            .I(N__5779));
    LocalMux I__1209 (
            .O(N__5794),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__1208 (
            .O(N__5789),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__1207 (
            .O(N__5784),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__1206 (
            .O(N__5779),
            .I(\U409_TICK.TICK603_14 ));
    InMux I__1205 (
            .O(N__5770),
            .I(N__5762));
    CascadeMux I__1204 (
            .O(N__5769),
            .I(N__5759));
    CascadeMux I__1203 (
            .O(N__5768),
            .I(N__5755));
    InMux I__1202 (
            .O(N__5767),
            .I(N__5750));
    InMux I__1201 (
            .O(N__5766),
            .I(N__5750));
    InMux I__1200 (
            .O(N__5765),
            .I(N__5747));
    LocalMux I__1199 (
            .O(N__5762),
            .I(N__5744));
    InMux I__1198 (
            .O(N__5759),
            .I(N__5739));
    InMux I__1197 (
            .O(N__5758),
            .I(N__5739));
    InMux I__1196 (
            .O(N__5755),
            .I(N__5736));
    LocalMux I__1195 (
            .O(N__5750),
            .I(N__5733));
    LocalMux I__1194 (
            .O(N__5747),
            .I(N__5730));
    Odrv12 I__1193 (
            .O(N__5744),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__1192 (
            .O(N__5739),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__1191 (
            .O(N__5736),
            .I(\U409_TICK.TICK603_10 ));
    Odrv4 I__1190 (
            .O(N__5733),
            .I(\U409_TICK.TICK603_10 ));
    Odrv4 I__1189 (
            .O(N__5730),
            .I(\U409_TICK.TICK603_10 ));
    InMux I__1188 (
            .O(N__5719),
            .I(N__5716));
    LocalMux I__1187 (
            .O(N__5716),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ));
    InMux I__1186 (
            .O(N__5713),
            .I(N__5709));
    InMux I__1185 (
            .O(N__5712),
            .I(N__5706));
    LocalMux I__1184 (
            .O(N__5709),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    LocalMux I__1183 (
            .O(N__5706),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    CascadeMux I__1182 (
            .O(N__5701),
            .I(N__5698));
    InMux I__1181 (
            .O(N__5698),
            .I(N__5693));
    InMux I__1180 (
            .O(N__5697),
            .I(N__5690));
    CascadeMux I__1179 (
            .O(N__5696),
            .I(N__5685));
    LocalMux I__1178 (
            .O(N__5693),
            .I(N__5680));
    LocalMux I__1177 (
            .O(N__5690),
            .I(N__5680));
    InMux I__1176 (
            .O(N__5689),
            .I(N__5673));
    InMux I__1175 (
            .O(N__5688),
            .I(N__5673));
    InMux I__1174 (
            .O(N__5685),
            .I(N__5673));
    Span4Mux_h I__1173 (
            .O(N__5680),
            .I(N__5670));
    LocalMux I__1172 (
            .O(N__5673),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    Odrv4 I__1171 (
            .O(N__5670),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    CascadeMux I__1170 (
            .O(N__5665),
            .I(\U409_TRANSFER_ACK.N_9_cascade_ ));
    IoInMux I__1169 (
            .O(N__5662),
            .I(N__5659));
    LocalMux I__1168 (
            .O(N__5659),
            .I(N__5656));
    Span4Mux_s3_v I__1167 (
            .O(N__5656),
            .I(N__5653));
    Span4Mux_v I__1166 (
            .O(N__5653),
            .I(N__5650));
    Span4Mux_v I__1165 (
            .O(N__5650),
            .I(N__5647));
    Span4Mux_h I__1164 (
            .O(N__5647),
            .I(N__5643));
    InMux I__1163 (
            .O(N__5646),
            .I(N__5640));
    Odrv4 I__1162 (
            .O(N__5643),
            .I(TICK60_c));
    LocalMux I__1161 (
            .O(N__5640),
            .I(TICK60_c));
    InMux I__1160 (
            .O(N__5635),
            .I(N__5632));
    LocalMux I__1159 (
            .O(N__5632),
            .I(\U409_TRANSFER_ACK.N_4 ));
    InMux I__1158 (
            .O(N__5629),
            .I(N__5626));
    LocalMux I__1157 (
            .O(N__5626),
            .I(N__5622));
    CascadeMux I__1156 (
            .O(N__5625),
            .I(N__5618));
    Span4Mux_h I__1155 (
            .O(N__5622),
            .I(N__5614));
    InMux I__1154 (
            .O(N__5621),
            .I(N__5609));
    InMux I__1153 (
            .O(N__5618),
            .I(N__5609));
    InMux I__1152 (
            .O(N__5617),
            .I(N__5606));
    Odrv4 I__1151 (
            .O(N__5614),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__1150 (
            .O(N__5609),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__1149 (
            .O(N__5606),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    InMux I__1148 (
            .O(N__5599),
            .I(N__5592));
    InMux I__1147 (
            .O(N__5598),
            .I(N__5592));
    InMux I__1146 (
            .O(N__5597),
            .I(N__5589));
    LocalMux I__1145 (
            .O(N__5592),
            .I(N__5584));
    LocalMux I__1144 (
            .O(N__5589),
            .I(N__5584));
    Odrv4 I__1143 (
            .O(N__5584),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    CascadeMux I__1142 (
            .O(N__5581),
            .I(\U409_TRANSFER_ACK.N_4_cascade_ ));
    InMux I__1141 (
            .O(N__5578),
            .I(N__5572));
    InMux I__1140 (
            .O(N__5577),
            .I(N__5569));
    InMux I__1139 (
            .O(N__5576),
            .I(N__5564));
    InMux I__1138 (
            .O(N__5575),
            .I(N__5564));
    LocalMux I__1137 (
            .O(N__5572),
            .I(N__5561));
    LocalMux I__1136 (
            .O(N__5569),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__1135 (
            .O(N__5564),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    Odrv4 I__1134 (
            .O(N__5561),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    InMux I__1133 (
            .O(N__5554),
            .I(N__5551));
    LocalMux I__1132 (
            .O(N__5551),
            .I(\U409_TRANSFER_ACK.N_5 ));
    IoInMux I__1131 (
            .O(N__5548),
            .I(N__5543));
    CascadeMux I__1130 (
            .O(N__5547),
            .I(N__5538));
    CascadeMux I__1129 (
            .O(N__5546),
            .I(N__5535));
    LocalMux I__1128 (
            .O(N__5543),
            .I(N__5531));
    CascadeMux I__1127 (
            .O(N__5542),
            .I(N__5528));
    InMux I__1126 (
            .O(N__5541),
            .I(N__5524));
    InMux I__1125 (
            .O(N__5538),
            .I(N__5521));
    InMux I__1124 (
            .O(N__5535),
            .I(N__5518));
    InMux I__1123 (
            .O(N__5534),
            .I(N__5515));
    IoSpan4Mux I__1122 (
            .O(N__5531),
            .I(N__5512));
    InMux I__1121 (
            .O(N__5528),
            .I(N__5507));
    InMux I__1120 (
            .O(N__5527),
            .I(N__5507));
    LocalMux I__1119 (
            .O(N__5524),
            .I(N__5500));
    LocalMux I__1118 (
            .O(N__5521),
            .I(N__5500));
    LocalMux I__1117 (
            .O(N__5518),
            .I(N__5500));
    LocalMux I__1116 (
            .O(N__5515),
            .I(N__5497));
    Span4Mux_s0_v I__1115 (
            .O(N__5512),
            .I(N__5493));
    LocalMux I__1114 (
            .O(N__5507),
            .I(N__5490));
    Span4Mux_v I__1113 (
            .O(N__5500),
            .I(N__5487));
    Span4Mux_v I__1112 (
            .O(N__5497),
            .I(N__5484));
    InMux I__1111 (
            .O(N__5496),
            .I(N__5481));
    Sp12to4 I__1110 (
            .O(N__5493),
            .I(N__5478));
    Span4Mux_h I__1109 (
            .O(N__5490),
            .I(N__5475));
    Sp12to4 I__1108 (
            .O(N__5487),
            .I(N__5470));
    Sp12to4 I__1107 (
            .O(N__5484),
            .I(N__5470));
    LocalMux I__1106 (
            .O(N__5481),
            .I(N__5467));
    Span12Mux_v I__1105 (
            .O(N__5478),
            .I(N__5458));
    Sp12to4 I__1104 (
            .O(N__5475),
            .I(N__5458));
    Span12Mux_h I__1103 (
            .O(N__5470),
            .I(N__5458));
    Span12Mux_h I__1102 (
            .O(N__5467),
            .I(N__5458));
    Span12Mux_v I__1101 (
            .O(N__5458),
            .I(N__5455));
    Odrv12 I__1100 (
            .O(N__5455),
            .I(CLK40_IN_c));
    InMux I__1099 (
            .O(N__5452),
            .I(N__5449));
    LocalMux I__1098 (
            .O(N__5449),
            .I(\U409_TRANSFER_ACK.m8_ns_1 ));
    InMux I__1097 (
            .O(N__5446),
            .I(N__5443));
    LocalMux I__1096 (
            .O(N__5443),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ));
    InMux I__1095 (
            .O(N__5440),
            .I(\U409_TICK.un3_COUNTER60_1_cry_12 ));
    InMux I__1094 (
            .O(N__5437),
            .I(\U409_TICK.un3_COUNTER60_1_cry_13 ));
    InMux I__1093 (
            .O(N__5434),
            .I(\U409_TICK.un3_COUNTER60_1_cry_14 ));
    InMux I__1092 (
            .O(N__5431),
            .I(\U409_TICK.un3_COUNTER60_1_cry_15 ));
    InMux I__1091 (
            .O(N__5428),
            .I(N__5424));
    InMux I__1090 (
            .O(N__5427),
            .I(N__5421));
    LocalMux I__1089 (
            .O(N__5424),
            .I(N__5416));
    LocalMux I__1088 (
            .O(N__5421),
            .I(N__5416));
    Span4Mux_v I__1087 (
            .O(N__5416),
            .I(N__5413));
    Odrv4 I__1086 (
            .O(N__5413),
            .I(U409_ADDRESS_DECODE_un1_RAMSPACEn));
    InMux I__1085 (
            .O(N__5410),
            .I(N__5406));
    InMux I__1084 (
            .O(N__5409),
            .I(N__5403));
    LocalMux I__1083 (
            .O(N__5406),
            .I(N__5397));
    LocalMux I__1082 (
            .O(N__5403),
            .I(N__5397));
    InMux I__1081 (
            .O(N__5402),
            .I(N__5394));
    Odrv12 I__1080 (
            .O(N__5397),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn));
    LocalMux I__1079 (
            .O(N__5394),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn));
    IoInMux I__1078 (
            .O(N__5389),
            .I(N__5386));
    LocalMux I__1077 (
            .O(N__5386),
            .I(N__5383));
    IoSpan4Mux I__1076 (
            .O(N__5383),
            .I(N__5380));
    Span4Mux_s2_v I__1075 (
            .O(N__5380),
            .I(N__5377));
    Sp12to4 I__1074 (
            .O(N__5377),
            .I(N__5374));
    Span12Mux_s10_v I__1073 (
            .O(N__5374),
            .I(N__5371));
    Odrv12 I__1072 (
            .O(N__5371),
            .I(BUFENn_c));
    CascadeMux I__1071 (
            .O(N__5368),
            .I(\U409_TRANSFER_ACK.i6_mux_0_cascade_ ));
    InMux I__1070 (
            .O(N__5365),
            .I(\U409_TICK.un3_COUNTER60_1_cry_3 ));
    InMux I__1069 (
            .O(N__5362),
            .I(N__5358));
    InMux I__1068 (
            .O(N__5361),
            .I(N__5355));
    LocalMux I__1067 (
            .O(N__5358),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    LocalMux I__1066 (
            .O(N__5355),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    InMux I__1065 (
            .O(N__5350),
            .I(\U409_TICK.un3_COUNTER60_1_cry_4 ));
    InMux I__1064 (
            .O(N__5347),
            .I(\U409_TICK.un3_COUNTER60_1_cry_5 ));
    InMux I__1063 (
            .O(N__5344),
            .I(\U409_TICK.un3_COUNTER60_1_cry_6 ));
    InMux I__1062 (
            .O(N__5341),
            .I(N__5338));
    LocalMux I__1061 (
            .O(N__5338),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ));
    InMux I__1060 (
            .O(N__5335),
            .I(\U409_TICK.un3_COUNTER60_1_cry_7 ));
    InMux I__1059 (
            .O(N__5332),
            .I(bfn_12_10_0_));
    InMux I__1058 (
            .O(N__5329),
            .I(\U409_TICK.un3_COUNTER60_1_cry_9 ));
    InMux I__1057 (
            .O(N__5326),
            .I(\U409_TICK.un3_COUNTER60_1_cry_10 ));
    InMux I__1056 (
            .O(N__5323),
            .I(\U409_TICK.un3_COUNTER60_1_cry_11 ));
    InMux I__1055 (
            .O(N__5320),
            .I(N__5314));
    InMux I__1054 (
            .O(N__5319),
            .I(N__5309));
    InMux I__1053 (
            .O(N__5318),
            .I(N__5309));
    InMux I__1052 (
            .O(N__5317),
            .I(N__5306));
    LocalMux I__1051 (
            .O(N__5314),
            .I(N__5296));
    LocalMux I__1050 (
            .O(N__5309),
            .I(N__5296));
    LocalMux I__1049 (
            .O(N__5306),
            .I(N__5296));
    InMux I__1048 (
            .O(N__5305),
            .I(N__5293));
    InMux I__1047 (
            .O(N__5304),
            .I(N__5290));
    InMux I__1046 (
            .O(N__5303),
            .I(N__5287));
    Span4Mux_v I__1045 (
            .O(N__5296),
            .I(N__5282));
    LocalMux I__1044 (
            .O(N__5293),
            .I(N__5282));
    LocalMux I__1043 (
            .O(N__5290),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1042 (
            .O(N__5287),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    Odrv4 I__1041 (
            .O(N__5282),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    InMux I__1040 (
            .O(N__5275),
            .I(N__5270));
    CascadeMux I__1039 (
            .O(N__5274),
            .I(N__5265));
    InMux I__1038 (
            .O(N__5273),
            .I(N__5261));
    LocalMux I__1037 (
            .O(N__5270),
            .I(N__5258));
    InMux I__1036 (
            .O(N__5269),
            .I(N__5255));
    InMux I__1035 (
            .O(N__5268),
            .I(N__5252));
    InMux I__1034 (
            .O(N__5265),
            .I(N__5246));
    InMux I__1033 (
            .O(N__5264),
            .I(N__5246));
    LocalMux I__1032 (
            .O(N__5261),
            .I(N__5241));
    Span4Mux_v I__1031 (
            .O(N__5258),
            .I(N__5241));
    LocalMux I__1030 (
            .O(N__5255),
            .I(N__5236));
    LocalMux I__1029 (
            .O(N__5252),
            .I(N__5236));
    InMux I__1028 (
            .O(N__5251),
            .I(N__5233));
    LocalMux I__1027 (
            .O(N__5246),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    Odrv4 I__1026 (
            .O(N__5241),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    Odrv4 I__1025 (
            .O(N__5236),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1024 (
            .O(N__5233),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    CascadeMux I__1023 (
            .O(N__5224),
            .I(N__5220));
    CascadeMux I__1022 (
            .O(N__5223),
            .I(N__5216));
    InMux I__1021 (
            .O(N__5220),
            .I(N__5206));
    InMux I__1020 (
            .O(N__5219),
            .I(N__5206));
    InMux I__1019 (
            .O(N__5216),
            .I(N__5206));
    InMux I__1018 (
            .O(N__5215),
            .I(N__5203));
    InMux I__1017 (
            .O(N__5214),
            .I(N__5198));
    CascadeMux I__1016 (
            .O(N__5213),
            .I(N__5195));
    LocalMux I__1015 (
            .O(N__5206),
            .I(N__5190));
    LocalMux I__1014 (
            .O(N__5203),
            .I(N__5190));
    InMux I__1013 (
            .O(N__5202),
            .I(N__5185));
    InMux I__1012 (
            .O(N__5201),
            .I(N__5185));
    LocalMux I__1011 (
            .O(N__5198),
            .I(N__5182));
    InMux I__1010 (
            .O(N__5195),
            .I(N__5179));
    Span4Mux_v I__1009 (
            .O(N__5190),
            .I(N__5176));
    LocalMux I__1008 (
            .O(N__5185),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    Odrv4 I__1007 (
            .O(N__5182),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1006 (
            .O(N__5179),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    Odrv4 I__1005 (
            .O(N__5176),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    InMux I__1004 (
            .O(N__5167),
            .I(N__5164));
    LocalMux I__1003 (
            .O(N__5164),
            .I(N__5157));
    InMux I__1002 (
            .O(N__5163),
            .I(N__5154));
    InMux I__1001 (
            .O(N__5162),
            .I(N__5151));
    InMux I__1000 (
            .O(N__5161),
            .I(N__5145));
    InMux I__999 (
            .O(N__5160),
            .I(N__5145));
    Span4Mux_h I__998 (
            .O(N__5157),
            .I(N__5142));
    LocalMux I__997 (
            .O(N__5154),
            .I(N__5137));
    LocalMux I__996 (
            .O(N__5151),
            .I(N__5137));
    InMux I__995 (
            .O(N__5150),
            .I(N__5134));
    LocalMux I__994 (
            .O(N__5145),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    Odrv4 I__993 (
            .O(N__5142),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    Odrv4 I__992 (
            .O(N__5137),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__991 (
            .O(N__5134),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    InMux I__990 (
            .O(N__5125),
            .I(N__5122));
    LocalMux I__989 (
            .O(N__5122),
            .I(N__5119));
    Odrv4 I__988 (
            .O(N__5119),
            .I(\U409_TRANSFER_ACK.N_36 ));
    CascadeMux I__987 (
            .O(N__5116),
            .I(N__5113));
    InMux I__986 (
            .O(N__5113),
            .I(N__5103));
    InMux I__985 (
            .O(N__5112),
            .I(N__5103));
    InMux I__984 (
            .O(N__5111),
            .I(N__5103));
    InMux I__983 (
            .O(N__5110),
            .I(N__5100));
    LocalMux I__982 (
            .O(N__5103),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__981 (
            .O(N__5100),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    InMux I__980 (
            .O(N__5095),
            .I(\U409_TICK.un3_COUNTER60_1_cry_1 ));
    InMux I__979 (
            .O(N__5092),
            .I(\U409_TICK.un3_COUNTER60_1_cry_2 ));
    CascadeMux I__978 (
            .O(N__5089),
            .I(N__5083));
    CascadeMux I__977 (
            .O(N__5088),
            .I(N__5080));
    CascadeMux I__976 (
            .O(N__5087),
            .I(N__5077));
    CascadeMux I__975 (
            .O(N__5086),
            .I(N__5074));
    InMux I__974 (
            .O(N__5083),
            .I(N__5062));
    InMux I__973 (
            .O(N__5080),
            .I(N__5062));
    InMux I__972 (
            .O(N__5077),
            .I(N__5062));
    InMux I__971 (
            .O(N__5074),
            .I(N__5062));
    InMux I__970 (
            .O(N__5073),
            .I(N__5062));
    LocalMux I__969 (
            .O(N__5062),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    CascadeMux I__968 (
            .O(N__5059),
            .I(N__5053));
    CascadeMux I__967 (
            .O(N__5058),
            .I(N__5050));
    InMux I__966 (
            .O(N__5057),
            .I(N__5047));
    InMux I__965 (
            .O(N__5056),
            .I(N__5044));
    InMux I__964 (
            .O(N__5053),
            .I(N__5041));
    InMux I__963 (
            .O(N__5050),
            .I(N__5038));
    LocalMux I__962 (
            .O(N__5047),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__961 (
            .O(N__5044),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__960 (
            .O(N__5041),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__959 (
            .O(N__5038),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    InMux I__958 (
            .O(N__5029),
            .I(N__5023));
    InMux I__957 (
            .O(N__5028),
            .I(N__5020));
    InMux I__956 (
            .O(N__5027),
            .I(N__5015));
    InMux I__955 (
            .O(N__5026),
            .I(N__5015));
    LocalMux I__954 (
            .O(N__5023),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__953 (
            .O(N__5020),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__952 (
            .O(N__5015),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    InMux I__951 (
            .O(N__5008),
            .I(N__5002));
    InMux I__950 (
            .O(N__5007),
            .I(N__5002));
    LocalMux I__949 (
            .O(N__5002),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ));
    InMux I__948 (
            .O(N__4999),
            .I(N__4988));
    InMux I__947 (
            .O(N__4998),
            .I(N__4988));
    InMux I__946 (
            .O(N__4997),
            .I(N__4985));
    InMux I__945 (
            .O(N__4996),
            .I(N__4982));
    InMux I__944 (
            .O(N__4995),
            .I(N__4979));
    InMux I__943 (
            .O(N__4994),
            .I(N__4974));
    InMux I__942 (
            .O(N__4993),
            .I(N__4974));
    LocalMux I__941 (
            .O(N__4988),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__940 (
            .O(N__4985),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__939 (
            .O(N__4982),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__938 (
            .O(N__4979),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__937 (
            .O(N__4974),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    InMux I__936 (
            .O(N__4963),
            .I(N__4958));
    InMux I__935 (
            .O(N__4962),
            .I(N__4955));
    InMux I__934 (
            .O(N__4961),
            .I(N__4952));
    LocalMux I__933 (
            .O(N__4958),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__932 (
            .O(N__4955),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__931 (
            .O(N__4952),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    InMux I__930 (
            .O(N__4945),
            .I(N__4937));
    InMux I__929 (
            .O(N__4944),
            .I(N__4937));
    InMux I__928 (
            .O(N__4943),
            .I(N__4934));
    InMux I__927 (
            .O(N__4942),
            .I(N__4931));
    LocalMux I__926 (
            .O(N__4937),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__925 (
            .O(N__4934),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__924 (
            .O(N__4931),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    InMux I__923 (
            .O(N__4924),
            .I(N__4919));
    CascadeMux I__922 (
            .O(N__4923),
            .I(N__4916));
    InMux I__921 (
            .O(N__4922),
            .I(N__4913));
    LocalMux I__920 (
            .O(N__4919),
            .I(N__4910));
    InMux I__919 (
            .O(N__4916),
            .I(N__4907));
    LocalMux I__918 (
            .O(N__4913),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ));
    Odrv4 I__917 (
            .O(N__4910),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ));
    LocalMux I__916 (
            .O(N__4907),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ));
    InMux I__915 (
            .O(N__4900),
            .I(N__4892));
    InMux I__914 (
            .O(N__4899),
            .I(N__4892));
    InMux I__913 (
            .O(N__4898),
            .I(N__4887));
    InMux I__912 (
            .O(N__4897),
            .I(N__4884));
    LocalMux I__911 (
            .O(N__4892),
            .I(N__4881));
    InMux I__910 (
            .O(N__4891),
            .I(N__4876));
    InMux I__909 (
            .O(N__4890),
            .I(N__4876));
    LocalMux I__908 (
            .O(N__4887),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__907 (
            .O(N__4884),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    Odrv4 I__906 (
            .O(N__4881),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__905 (
            .O(N__4876),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    CascadeMux I__904 (
            .O(N__4867),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ));
    InMux I__903 (
            .O(N__4864),
            .I(N__4857));
    InMux I__902 (
            .O(N__4863),
            .I(N__4852));
    InMux I__901 (
            .O(N__4862),
            .I(N__4852));
    InMux I__900 (
            .O(N__4861),
            .I(N__4847));
    InMux I__899 (
            .O(N__4860),
            .I(N__4847));
    LocalMux I__898 (
            .O(N__4857),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__897 (
            .O(N__4852),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__896 (
            .O(N__4847),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    InMux I__895 (
            .O(N__4840),
            .I(N__4837));
    LocalMux I__894 (
            .O(N__4837),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5 ));
    InMux I__893 (
            .O(N__4834),
            .I(N__4831));
    LocalMux I__892 (
            .O(N__4831),
            .I(N__4826));
    InMux I__891 (
            .O(N__4830),
            .I(N__4823));
    CascadeMux I__890 (
            .O(N__4829),
            .I(N__4820));
    Span4Mux_h I__889 (
            .O(N__4826),
            .I(N__4815));
    LocalMux I__888 (
            .O(N__4823),
            .I(N__4815));
    InMux I__887 (
            .O(N__4820),
            .I(N__4812));
    Span4Mux_h I__886 (
            .O(N__4815),
            .I(N__4806));
    LocalMux I__885 (
            .O(N__4812),
            .I(N__4806));
    InMux I__884 (
            .O(N__4811),
            .I(N__4803));
    Span4Mux_v I__883 (
            .O(N__4806),
            .I(N__4798));
    LocalMux I__882 (
            .O(N__4803),
            .I(N__4798));
    Span4Mux_h I__881 (
            .O(N__4798),
            .I(N__4795));
    Odrv4 I__880 (
            .O(N__4795),
            .I(U409_ADDRESS_DECODE_ROMEN_1));
    CascadeMux I__879 (
            .O(N__4792),
            .I(N__4789));
    InMux I__878 (
            .O(N__4789),
            .I(N__4785));
    CascadeMux I__877 (
            .O(N__4788),
            .I(N__4782));
    LocalMux I__876 (
            .O(N__4785),
            .I(N__4779));
    InMux I__875 (
            .O(N__4782),
            .I(N__4776));
    Span4Mux_h I__874 (
            .O(N__4779),
            .I(N__4771));
    LocalMux I__873 (
            .O(N__4776),
            .I(N__4771));
    Span4Mux_h I__872 (
            .O(N__4771),
            .I(N__4768));
    Odrv4 I__871 (
            .O(N__4768),
            .I(\U409_TRANSFER_ACK.N_23 ));
    InMux I__870 (
            .O(N__4765),
            .I(N__4762));
    LocalMux I__869 (
            .O(N__4762),
            .I(N__4759));
    Sp12to4 I__868 (
            .O(N__4759),
            .I(N__4756));
    Span12Mux_s9_v I__867 (
            .O(N__4756),
            .I(N__4753));
    Span12Mux_h I__866 (
            .O(N__4753),
            .I(N__4750));
    Odrv12 I__865 (
            .O(N__4750),
            .I(TACKn_in));
    SRMux I__864 (
            .O(N__4747),
            .I(N__4743));
    SRMux I__863 (
            .O(N__4746),
            .I(N__4740));
    LocalMux I__862 (
            .O(N__4743),
            .I(N__4736));
    LocalMux I__861 (
            .O(N__4740),
            .I(N__4733));
    SRMux I__860 (
            .O(N__4739),
            .I(N__4730));
    Span4Mux_h I__859 (
            .O(N__4736),
            .I(N__4727));
    Span4Mux_h I__858 (
            .O(N__4733),
            .I(N__4722));
    LocalMux I__857 (
            .O(N__4730),
            .I(N__4722));
    Span4Mux_v I__856 (
            .O(N__4727),
            .I(N__4716));
    Span4Mux_v I__855 (
            .O(N__4722),
            .I(N__4716));
    SRMux I__854 (
            .O(N__4721),
            .I(N__4713));
    Span4Mux_v I__853 (
            .O(N__4716),
            .I(N__4708));
    LocalMux I__852 (
            .O(N__4713),
            .I(N__4708));
    Span4Mux_v I__851 (
            .O(N__4708),
            .I(N__4705));
    Span4Mux_v I__850 (
            .O(N__4705),
            .I(N__4702));
    Odrv4 I__849 (
            .O(N__4702),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    IoInMux I__848 (
            .O(N__4699),
            .I(N__4696));
    LocalMux I__847 (
            .O(N__4696),
            .I(N__4693));
    Span4Mux_s2_v I__846 (
            .O(N__4693),
            .I(N__4690));
    Span4Mux_v I__845 (
            .O(N__4690),
            .I(N__4687));
    Odrv4 I__844 (
            .O(N__4687),
            .I(CONSTANT_ONE_NET));
    InMux I__843 (
            .O(N__4684),
            .I(N__4681));
    LocalMux I__842 (
            .O(N__4681),
            .I(N__4678));
    Odrv4 I__841 (
            .O(N__4678),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_1_0 ));
    CascadeMux I__840 (
            .O(N__4675),
            .I(N__4672));
    InMux I__839 (
            .O(N__4672),
            .I(N__4669));
    LocalMux I__838 (
            .O(N__4669),
            .I(N__4665));
    InMux I__837 (
            .O(N__4668),
            .I(N__4662));
    Span4Mux_v I__836 (
            .O(N__4665),
            .I(N__4657));
    LocalMux I__835 (
            .O(N__4662),
            .I(N__4657));
    Odrv4 I__834 (
            .O(N__4657),
            .I(\U409_TRANSFER_ACK.N_35_1 ));
    InMux I__833 (
            .O(N__4654),
            .I(N__4651));
    LocalMux I__832 (
            .O(N__4651),
            .I(N__4648));
    Odrv12 I__831 (
            .O(N__4648),
            .I(\U409_TRANSFER_ACK.N_29 ));
    CascadeMux I__830 (
            .O(N__4645),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_3_cascade_ ));
    InMux I__829 (
            .O(N__4642),
            .I(N__4639));
    LocalMux I__828 (
            .O(N__4639),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ));
    InMux I__827 (
            .O(N__4636),
            .I(N__4630));
    InMux I__826 (
            .O(N__4635),
            .I(N__4630));
    LocalMux I__825 (
            .O(N__4630),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ));
    CascadeMux I__824 (
            .O(N__4627),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_2_cascade_ ));
    InMux I__823 (
            .O(N__4624),
            .I(N__4620));
    InMux I__822 (
            .O(N__4623),
            .I(N__4617));
    LocalMux I__821 (
            .O(N__4620),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    LocalMux I__820 (
            .O(N__4617),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    InMux I__819 (
            .O(N__4612),
            .I(N__4609));
    LocalMux I__818 (
            .O(N__4609),
            .I(N__4605));
    InMux I__817 (
            .O(N__4608),
            .I(N__4600));
    Span4Mux_v I__816 (
            .O(N__4605),
            .I(N__4597));
    InMux I__815 (
            .O(N__4604),
            .I(N__4592));
    InMux I__814 (
            .O(N__4603),
            .I(N__4592));
    LocalMux I__813 (
            .O(N__4600),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    Odrv4 I__812 (
            .O(N__4597),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    LocalMux I__811 (
            .O(N__4592),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    InMux I__810 (
            .O(N__4585),
            .I(N__4582));
    LocalMux I__809 (
            .O(N__4582),
            .I(N__4579));
    Odrv4 I__808 (
            .O(N__4579),
            .I(\U409_TRANSFER_ACK.N_47 ));
    InMux I__807 (
            .O(N__4576),
            .I(N__4573));
    LocalMux I__806 (
            .O(N__4573),
            .I(\U409_TRANSFER_ACK.N_142 ));
    InMux I__805 (
            .O(N__4570),
            .I(N__4564));
    InMux I__804 (
            .O(N__4569),
            .I(N__4564));
    LocalMux I__803 (
            .O(N__4564),
            .I(N__4561));
    Span12Mux_v I__802 (
            .O(N__4561),
            .I(N__4558));
    Odrv12 I__801 (
            .O(N__4558),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_0 ));
    InMux I__800 (
            .O(N__4555),
            .I(N__4550));
    InMux I__799 (
            .O(N__4554),
            .I(N__4547));
    CascadeMux I__798 (
            .O(N__4553),
            .I(N__4544));
    LocalMux I__797 (
            .O(N__4550),
            .I(N__4538));
    LocalMux I__796 (
            .O(N__4547),
            .I(N__4538));
    InMux I__795 (
            .O(N__4544),
            .I(N__4533));
    InMux I__794 (
            .O(N__4543),
            .I(N__4533));
    Span4Mux_v I__793 (
            .O(N__4538),
            .I(N__4527));
    LocalMux I__792 (
            .O(N__4533),
            .I(N__4527));
    InMux I__791 (
            .O(N__4532),
            .I(N__4524));
    Span4Mux_v I__790 (
            .O(N__4527),
            .I(N__4521));
    LocalMux I__789 (
            .O(N__4524),
            .I(N__4518));
    Sp12to4 I__788 (
            .O(N__4521),
            .I(N__4515));
    Span12Mux_h I__787 (
            .O(N__4518),
            .I(N__4512));
    Span12Mux_h I__786 (
            .O(N__4515),
            .I(N__4509));
    Span12Mux_v I__785 (
            .O(N__4512),
            .I(N__4506));
    Span12Mux_v I__784 (
            .O(N__4509),
            .I(N__4503));
    Odrv12 I__783 (
            .O(N__4506),
            .I(TSn_c));
    Odrv12 I__782 (
            .O(N__4503),
            .I(TSn_c));
    InMux I__781 (
            .O(N__4498),
            .I(N__4493));
    InMux I__780 (
            .O(N__4497),
            .I(N__4488));
    InMux I__779 (
            .O(N__4496),
            .I(N__4488));
    LocalMux I__778 (
            .O(N__4493),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    LocalMux I__777 (
            .O(N__4488),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    CascadeMux I__776 (
            .O(N__4483),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_cascade_ ));
    CEMux I__775 (
            .O(N__4480),
            .I(N__4477));
    LocalMux I__774 (
            .O(N__4477),
            .I(N__4474));
    Span4Mux_h I__773 (
            .O(N__4474),
            .I(N__4471));
    Odrv4 I__772 (
            .O(N__4471),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1_0 ));
    IoInMux I__771 (
            .O(N__4468),
            .I(N__4465));
    LocalMux I__770 (
            .O(N__4465),
            .I(N__4462));
    IoSpan4Mux I__769 (
            .O(N__4462),
            .I(N__4459));
    Span4Mux_s1_v I__768 (
            .O(N__4459),
            .I(N__4456));
    Sp12to4 I__767 (
            .O(N__4456),
            .I(N__4453));
    Span12Mux_v I__766 (
            .O(N__4453),
            .I(N__4450));
    Odrv12 I__765 (
            .O(N__4450),
            .I(U409_ADDRESS_DECODE_un1_RAMSPACEn_i));
    InMux I__764 (
            .O(N__4447),
            .I(N__4443));
    InMux I__763 (
            .O(N__4446),
            .I(N__4440));
    LocalMux I__762 (
            .O(N__4443),
            .I(N__4432));
    LocalMux I__761 (
            .O(N__4440),
            .I(N__4432));
    InMux I__760 (
            .O(N__4439),
            .I(N__4429));
    InMux I__759 (
            .O(N__4438),
            .I(N__4426));
    InMux I__758 (
            .O(N__4437),
            .I(N__4420));
    Span4Mux_v I__757 (
            .O(N__4432),
            .I(N__4417));
    LocalMux I__756 (
            .O(N__4429),
            .I(N__4412));
    LocalMux I__755 (
            .O(N__4426),
            .I(N__4412));
    InMux I__754 (
            .O(N__4425),
            .I(N__4409));
    InMux I__753 (
            .O(N__4424),
            .I(N__4406));
    InMux I__752 (
            .O(N__4423),
            .I(N__4403));
    LocalMux I__751 (
            .O(N__4420),
            .I(N__4400));
    Span4Mux_h I__750 (
            .O(N__4417),
            .I(N__4395));
    Span4Mux_v I__749 (
            .O(N__4412),
            .I(N__4395));
    LocalMux I__748 (
            .O(N__4409),
            .I(N__4390));
    LocalMux I__747 (
            .O(N__4406),
            .I(N__4390));
    LocalMux I__746 (
            .O(N__4403),
            .I(N__4386));
    Span4Mux_v I__745 (
            .O(N__4400),
            .I(N__4383));
    Span4Mux_h I__744 (
            .O(N__4395),
            .I(N__4378));
    Span4Mux_v I__743 (
            .O(N__4390),
            .I(N__4378));
    InMux I__742 (
            .O(N__4389),
            .I(N__4375));
    Span12Mux_v I__741 (
            .O(N__4386),
            .I(N__4366));
    Sp12to4 I__740 (
            .O(N__4383),
            .I(N__4366));
    Sp12to4 I__739 (
            .O(N__4378),
            .I(N__4366));
    LocalMux I__738 (
            .O(N__4375),
            .I(N__4366));
    Odrv12 I__737 (
            .O(N__4366),
            .I(A_c_21));
    InMux I__736 (
            .O(N__4363),
            .I(N__4359));
    CascadeMux I__735 (
            .O(N__4362),
            .I(N__4356));
    LocalMux I__734 (
            .O(N__4359),
            .I(N__4352));
    InMux I__733 (
            .O(N__4356),
            .I(N__4349));
    InMux I__732 (
            .O(N__4355),
            .I(N__4346));
    Span4Mux_v I__731 (
            .O(N__4352),
            .I(N__4343));
    LocalMux I__730 (
            .O(N__4349),
            .I(N__4338));
    LocalMux I__729 (
            .O(N__4346),
            .I(N__4338));
    Span4Mux_h I__728 (
            .O(N__4343),
            .I(N__4333));
    Span4Mux_v I__727 (
            .O(N__4338),
            .I(N__4333));
    Sp12to4 I__726 (
            .O(N__4333),
            .I(N__4330));
    Span12Mux_h I__725 (
            .O(N__4330),
            .I(N__4327));
    Span12Mux_v I__724 (
            .O(N__4327),
            .I(N__4324));
    Odrv12 I__723 (
            .O(N__4324),
            .I(OVL_c));
    InMux I__722 (
            .O(N__4321),
            .I(N__4317));
    InMux I__721 (
            .O(N__4320),
            .I(N__4314));
    LocalMux I__720 (
            .O(N__4317),
            .I(N__4309));
    LocalMux I__719 (
            .O(N__4314),
            .I(N__4309));
    Span4Mux_v I__718 (
            .O(N__4309),
            .I(N__4305));
    InMux I__717 (
            .O(N__4308),
            .I(N__4302));
    Span4Mux_h I__716 (
            .O(N__4305),
            .I(N__4297));
    LocalMux I__715 (
            .O(N__4302),
            .I(N__4297));
    Odrv4 I__714 (
            .O(N__4297),
            .I(U409_ADDRESS_DECODE_LOWROM_3));
    CascadeMux I__713 (
            .O(N__4294),
            .I(N__4291));
    InMux I__712 (
            .O(N__4291),
            .I(N__4287));
    InMux I__711 (
            .O(N__4290),
            .I(N__4284));
    LocalMux I__710 (
            .O(N__4287),
            .I(N__4281));
    LocalMux I__709 (
            .O(N__4284),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    Odrv4 I__708 (
            .O(N__4281),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    InMux I__707 (
            .O(N__4276),
            .I(N__4273));
    LocalMux I__706 (
            .O(N__4273),
            .I(N__4270));
    Odrv12 I__705 (
            .O(N__4270),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    InMux I__704 (
            .O(N__4267),
            .I(N__4264));
    LocalMux I__703 (
            .O(N__4264),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23 ));
    CascadeMux I__702 (
            .O(N__4261),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_cascade_ ));
    CascadeMux I__701 (
            .O(N__4258),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ));
    InMux I__700 (
            .O(N__4255),
            .I(N__4252));
    LocalMux I__699 (
            .O(N__4252),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    CascadeMux I__698 (
            .O(N__4249),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ));
    CascadeMux I__697 (
            .O(N__4246),
            .I(\U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ));
    IoInMux I__696 (
            .O(N__4243),
            .I(N__4240));
    LocalMux I__695 (
            .O(N__4240),
            .I(N__4235));
    IoInMux I__694 (
            .O(N__4239),
            .I(N__4232));
    IoInMux I__693 (
            .O(N__4238),
            .I(N__4229));
    Span4Mux_s3_v I__692 (
            .O(N__4235),
            .I(N__4226));
    LocalMux I__691 (
            .O(N__4232),
            .I(N__4221));
    LocalMux I__690 (
            .O(N__4229),
            .I(N__4221));
    Span4Mux_v I__689 (
            .O(N__4226),
            .I(N__4218));
    Span12Mux_s7_v I__688 (
            .O(N__4221),
            .I(N__4215));
    Sp12to4 I__687 (
            .O(N__4218),
            .I(N__4212));
    Span12Mux_v I__686 (
            .O(N__4215),
            .I(N__4209));
    Span12Mux_s7_h I__685 (
            .O(N__4212),
            .I(N__4206));
    Span12Mux_h I__684 (
            .O(N__4209),
            .I(N__4201));
    Span12Mux_v I__683 (
            .O(N__4206),
            .I(N__4198));
    InMux I__682 (
            .O(N__4205),
            .I(N__4195));
    InMux I__681 (
            .O(N__4204),
            .I(N__4192));
    Odrv12 I__680 (
            .O(N__4201),
            .I(TACK_OUTn));
    Odrv12 I__679 (
            .O(N__4198),
            .I(TACK_OUTn));
    LocalMux I__678 (
            .O(N__4195),
            .I(TACK_OUTn));
    LocalMux I__677 (
            .O(N__4192),
            .I(TACK_OUTn));
    InMux I__676 (
            .O(N__4183),
            .I(N__4177));
    InMux I__675 (
            .O(N__4182),
            .I(N__4170));
    InMux I__674 (
            .O(N__4181),
            .I(N__4170));
    InMux I__673 (
            .O(N__4180),
            .I(N__4170));
    LocalMux I__672 (
            .O(N__4177),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    LocalMux I__671 (
            .O(N__4170),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    CascadeMux I__670 (
            .O(N__4165),
            .I(N__4162));
    InMux I__669 (
            .O(N__4162),
            .I(N__4156));
    InMux I__668 (
            .O(N__4161),
            .I(N__4153));
    InMux I__667 (
            .O(N__4160),
            .I(N__4148));
    InMux I__666 (
            .O(N__4159),
            .I(N__4148));
    LocalMux I__665 (
            .O(N__4156),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    LocalMux I__664 (
            .O(N__4153),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    LocalMux I__663 (
            .O(N__4148),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    InMux I__662 (
            .O(N__4141),
            .I(N__4137));
    InMux I__661 (
            .O(N__4140),
            .I(N__4134));
    LocalMux I__660 (
            .O(N__4137),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    LocalMux I__659 (
            .O(N__4134),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    InMux I__658 (
            .O(N__4129),
            .I(N__4126));
    LocalMux I__657 (
            .O(N__4126),
            .I(\U409_TRANSFER_ACK.N_35 ));
    IoInMux I__656 (
            .O(N__4123),
            .I(N__4120));
    LocalMux I__655 (
            .O(N__4120),
            .I(N__4117));
    IoSpan4Mux I__654 (
            .O(N__4117),
            .I(N__4114));
    Sp12to4 I__653 (
            .O(N__4114),
            .I(N__4111));
    Span12Mux_s6_v I__652 (
            .O(N__4111),
            .I(N__4108));
    Span12Mux_v I__651 (
            .O(N__4108),
            .I(N__4104));
    InMux I__650 (
            .O(N__4107),
            .I(N__4101));
    Odrv12 I__649 (
            .O(N__4104),
            .I(ROMENn_c));
    LocalMux I__648 (
            .O(N__4101),
            .I(ROMENn_c));
    InMux I__647 (
            .O(N__4096),
            .I(N__4092));
    InMux I__646 (
            .O(N__4095),
            .I(N__4089));
    LocalMux I__645 (
            .O(N__4092),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    LocalMux I__644 (
            .O(N__4089),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    InMux I__643 (
            .O(N__4084),
            .I(N__4078));
    InMux I__642 (
            .O(N__4083),
            .I(N__4073));
    InMux I__641 (
            .O(N__4082),
            .I(N__4073));
    InMux I__640 (
            .O(N__4081),
            .I(N__4070));
    LocalMux I__639 (
            .O(N__4078),
            .I(N__4063));
    LocalMux I__638 (
            .O(N__4073),
            .I(N__4063));
    LocalMux I__637 (
            .O(N__4070),
            .I(N__4063));
    Span4Mux_v I__636 (
            .O(N__4063),
            .I(N__4060));
    Sp12to4 I__635 (
            .O(N__4060),
            .I(N__4057));
    Span12Mux_h I__634 (
            .O(N__4057),
            .I(N__4054));
    Odrv12 I__633 (
            .O(N__4054),
            .I(TM_c_1));
    InMux I__632 (
            .O(N__4051),
            .I(N__4048));
    LocalMux I__631 (
            .O(N__4048),
            .I(N__4042));
    InMux I__630 (
            .O(N__4047),
            .I(N__4037));
    InMux I__629 (
            .O(N__4046),
            .I(N__4037));
    InMux I__628 (
            .O(N__4045),
            .I(N__4034));
    Span4Mux_h I__627 (
            .O(N__4042),
            .I(N__4027));
    LocalMux I__626 (
            .O(N__4037),
            .I(N__4027));
    LocalMux I__625 (
            .O(N__4034),
            .I(N__4027));
    Span4Mux_v I__624 (
            .O(N__4027),
            .I(N__4024));
    Sp12to4 I__623 (
            .O(N__4024),
            .I(N__4021));
    Span12Mux_h I__622 (
            .O(N__4021),
            .I(N__4018));
    Odrv12 I__621 (
            .O(N__4018),
            .I(TM_c_0));
    InMux I__620 (
            .O(N__4015),
            .I(N__4007));
    InMux I__619 (
            .O(N__4014),
            .I(N__4007));
    InMux I__618 (
            .O(N__4013),
            .I(N__4004));
    InMux I__617 (
            .O(N__4012),
            .I(N__4001));
    LocalMux I__616 (
            .O(N__4007),
            .I(N__3998));
    LocalMux I__615 (
            .O(N__4004),
            .I(N__3995));
    LocalMux I__614 (
            .O(N__4001),
            .I(N__3990));
    Span4Mux_v I__613 (
            .O(N__3998),
            .I(N__3984));
    Span4Mux_v I__612 (
            .O(N__3995),
            .I(N__3984));
    InMux I__611 (
            .O(N__3994),
            .I(N__3981));
    InMux I__610 (
            .O(N__3993),
            .I(N__3978));
    Span4Mux_v I__609 (
            .O(N__3990),
            .I(N__3975));
    InMux I__608 (
            .O(N__3989),
            .I(N__3972));
    Sp12to4 I__607 (
            .O(N__3984),
            .I(N__3965));
    LocalMux I__606 (
            .O(N__3981),
            .I(N__3965));
    LocalMux I__605 (
            .O(N__3978),
            .I(N__3965));
    Sp12to4 I__604 (
            .O(N__3975),
            .I(N__3960));
    LocalMux I__603 (
            .O(N__3972),
            .I(N__3960));
    Odrv12 I__602 (
            .O(N__3965),
            .I(A_c_23));
    Odrv12 I__601 (
            .O(N__3960),
            .I(A_c_23));
    InMux I__600 (
            .O(N__3955),
            .I(N__3950));
    InMux I__599 (
            .O(N__3954),
            .I(N__3947));
    InMux I__598 (
            .O(N__3953),
            .I(N__3944));
    LocalMux I__597 (
            .O(N__3950),
            .I(N__3935));
    LocalMux I__596 (
            .O(N__3947),
            .I(N__3935));
    LocalMux I__595 (
            .O(N__3944),
            .I(N__3932));
    InMux I__594 (
            .O(N__3943),
            .I(N__3929));
    InMux I__593 (
            .O(N__3942),
            .I(N__3926));
    InMux I__592 (
            .O(N__3941),
            .I(N__3921));
    InMux I__591 (
            .O(N__3940),
            .I(N__3921));
    Span4Mux_h I__590 (
            .O(N__3935),
            .I(N__3913));
    Span4Mux_v I__589 (
            .O(N__3932),
            .I(N__3913));
    LocalMux I__588 (
            .O(N__3929),
            .I(N__3913));
    LocalMux I__587 (
            .O(N__3926),
            .I(N__3908));
    LocalMux I__586 (
            .O(N__3921),
            .I(N__3908));
    InMux I__585 (
            .O(N__3920),
            .I(N__3905));
    Span4Mux_h I__584 (
            .O(N__3913),
            .I(N__3902));
    Sp12to4 I__583 (
            .O(N__3908),
            .I(N__3897));
    LocalMux I__582 (
            .O(N__3905),
            .I(N__3897));
    Span4Mux_v I__581 (
            .O(N__3902),
            .I(N__3894));
    Span12Mux_v I__580 (
            .O(N__3897),
            .I(N__3891));
    Span4Mux_v I__579 (
            .O(N__3894),
            .I(N__3888));
    Odrv12 I__578 (
            .O(N__3891),
            .I(A_c_22));
    Odrv4 I__577 (
            .O(N__3888),
            .I(A_c_22));
    IoInMux I__576 (
            .O(N__3883),
            .I(N__3880));
    LocalMux I__575 (
            .O(N__3880),
            .I(N__3877));
    Span4Mux_s3_v I__574 (
            .O(N__3877),
            .I(N__3874));
    Span4Mux_h I__573 (
            .O(N__3874),
            .I(N__3871));
    Span4Mux_h I__572 (
            .O(N__3871),
            .I(N__3868));
    Span4Mux_h I__571 (
            .O(N__3868),
            .I(N__3865));
    Span4Mux_h I__570 (
            .O(N__3865),
            .I(N__3862));
    Span4Mux_v I__569 (
            .O(N__3862),
            .I(N__3859));
    Odrv4 I__568 (
            .O(N__3859),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn_i));
    InMux I__567 (
            .O(N__3856),
            .I(N__3847));
    InMux I__566 (
            .O(N__3855),
            .I(N__3847));
    InMux I__565 (
            .O(N__3854),
            .I(N__3844));
    InMux I__564 (
            .O(N__3853),
            .I(N__3839));
    InMux I__563 (
            .O(N__3852),
            .I(N__3839));
    LocalMux I__562 (
            .O(N__3847),
            .I(N__3836));
    LocalMux I__561 (
            .O(N__3844),
            .I(N__3833));
    LocalMux I__560 (
            .O(N__3839),
            .I(N__3830));
    Span4Mux_v I__559 (
            .O(N__3836),
            .I(N__3827));
    Span4Mux_v I__558 (
            .O(N__3833),
            .I(N__3822));
    Span4Mux_h I__557 (
            .O(N__3830),
            .I(N__3822));
    Span4Mux_h I__556 (
            .O(N__3827),
            .I(N__3819));
    Span4Mux_h I__555 (
            .O(N__3822),
            .I(N__3816));
    Odrv4 I__554 (
            .O(N__3819),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0 ));
    Odrv4 I__553 (
            .O(N__3816),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0 ));
    CascadeMux I__552 (
            .O(N__3811),
            .I(N__3808));
    InMux I__551 (
            .O(N__3808),
            .I(N__3802));
    InMux I__550 (
            .O(N__3807),
            .I(N__3802));
    LocalMux I__549 (
            .O(N__3802),
            .I(N__3799));
    Span4Mux_v I__548 (
            .O(N__3799),
            .I(N__3796));
    Odrv4 I__547 (
            .O(N__3796),
            .I(\U409_ADDRESS_DECODE.un2_REGSPACEn_0_0 ));
    CascadeMux I__546 (
            .O(N__3793),
            .I(N__3789));
    InMux I__545 (
            .O(N__3792),
            .I(N__3784));
    InMux I__544 (
            .O(N__3789),
            .I(N__3784));
    LocalMux I__543 (
            .O(N__3784),
            .I(N__3781));
    Odrv4 I__542 (
            .O(N__3781),
            .I(\U409_ADDRESS_DECODE.REG_SPACE_3_0 ));
    InMux I__541 (
            .O(N__3778),
            .I(N__3772));
    InMux I__540 (
            .O(N__3777),
            .I(N__3772));
    LocalMux I__539 (
            .O(N__3772),
            .I(\U409_ADDRESS_DECODE.REG_SPACEZ0Z_2 ));
    InMux I__538 (
            .O(N__3769),
            .I(N__3766));
    LocalMux I__537 (
            .O(N__3766),
            .I(N__3762));
    InMux I__536 (
            .O(N__3765),
            .I(N__3759));
    Span4Mux_h I__535 (
            .O(N__3762),
            .I(N__3754));
    LocalMux I__534 (
            .O(N__3759),
            .I(N__3754));
    Odrv4 I__533 (
            .O(N__3754),
            .I(U409_ADDRESS_DECODE_un1_RTC_ENn));
    IoInMux I__532 (
            .O(N__3751),
            .I(N__3748));
    LocalMux I__531 (
            .O(N__3748),
            .I(N__3745));
    Span12Mux_s10_v I__530 (
            .O(N__3745),
            .I(N__3742));
    Odrv12 I__529 (
            .O(N__3742),
            .I(PORTSIZE_0_i));
    CascadeMux I__528 (
            .O(N__3739),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0_0_cascade_ ));
    CEMux I__527 (
            .O(N__3736),
            .I(N__3733));
    LocalMux I__526 (
            .O(N__3733),
            .I(N__3730));
    Span4Mux_v I__525 (
            .O(N__3730),
            .I(N__3727));
    Odrv4 I__524 (
            .O(N__3727),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_0 ));
    InMux I__523 (
            .O(N__3724),
            .I(N__3721));
    LocalMux I__522 (
            .O(N__3721),
            .I(N__3718));
    Span4Mux_v I__521 (
            .O(N__3718),
            .I(N__3715));
    IoSpan4Mux I__520 (
            .O(N__3715),
            .I(N__3712));
    Odrv4 I__519 (
            .O(N__3712),
            .I(TT_c_1));
    InMux I__518 (
            .O(N__3709),
            .I(N__3706));
    LocalMux I__517 (
            .O(N__3706),
            .I(N__3703));
    Span4Mux_h I__516 (
            .O(N__3703),
            .I(N__3700));
    Span4Mux_v I__515 (
            .O(N__3700),
            .I(N__3697));
    Odrv4 I__514 (
            .O(N__3697),
            .I(TT_c_0));
    InMux I__513 (
            .O(N__3694),
            .I(N__3691));
    LocalMux I__512 (
            .O(N__3691),
            .I(N__3688));
    Odrv12 I__511 (
            .O(N__3688),
            .I(U409_ADDRESS_DECODE_AUTOVECTOR_2));
    CascadeMux I__510 (
            .O(N__3685),
            .I(U409_ADDRESS_DECODE_LOWROM_2_cascade_));
    InMux I__509 (
            .O(N__3682),
            .I(N__3679));
    LocalMux I__508 (
            .O(N__3679),
            .I(\U409_TRANSFER_ACK.N_45 ));
    CascadeMux I__507 (
            .O(N__3676),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2Z0Z_1_cascade_ ));
    CascadeMux I__506 (
            .O(N__3673),
            .I(N__3670));
    InMux I__505 (
            .O(N__3670),
            .I(N__3667));
    LocalMux I__504 (
            .O(N__3667),
            .I(N__3663));
    InMux I__503 (
            .O(N__3666),
            .I(N__3660));
    Odrv4 I__502 (
            .O(N__3663),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2 ));
    LocalMux I__501 (
            .O(N__3660),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2 ));
    CascadeMux I__500 (
            .O(N__3655),
            .I(N__3651));
    InMux I__499 (
            .O(N__3654),
            .I(N__3648));
    InMux I__498 (
            .O(N__3651),
            .I(N__3642));
    LocalMux I__497 (
            .O(N__3648),
            .I(N__3639));
    InMux I__496 (
            .O(N__3647),
            .I(N__3634));
    InMux I__495 (
            .O(N__3646),
            .I(N__3634));
    InMux I__494 (
            .O(N__3645),
            .I(N__3631));
    LocalMux I__493 (
            .O(N__3642),
            .I(N__3628));
    Span4Mux_v I__492 (
            .O(N__3639),
            .I(N__3625));
    LocalMux I__491 (
            .O(N__3634),
            .I(N__3620));
    LocalMux I__490 (
            .O(N__3631),
            .I(N__3620));
    Span4Mux_v I__489 (
            .O(N__3628),
            .I(N__3617));
    Span4Mux_h I__488 (
            .O(N__3625),
            .I(N__3612));
    Span4Mux_v I__487 (
            .O(N__3620),
            .I(N__3612));
    Sp12to4 I__486 (
            .O(N__3617),
            .I(N__3607));
    Sp12to4 I__485 (
            .O(N__3612),
            .I(N__3607));
    Span12Mux_h I__484 (
            .O(N__3607),
            .I(N__3604));
    Span12Mux_v I__483 (
            .O(N__3604),
            .I(N__3601));
    Odrv12 I__482 (
            .O(N__3601),
            .I(A_c_18));
    InMux I__481 (
            .O(N__3598),
            .I(N__3590));
    InMux I__480 (
            .O(N__3597),
            .I(N__3590));
    InMux I__479 (
            .O(N__3596),
            .I(N__3585));
    InMux I__478 (
            .O(N__3595),
            .I(N__3585));
    LocalMux I__477 (
            .O(N__3590),
            .I(N__3580));
    LocalMux I__476 (
            .O(N__3585),
            .I(N__3576));
    InMux I__475 (
            .O(N__3584),
            .I(N__3573));
    InMux I__474 (
            .O(N__3583),
            .I(N__3570));
    Span4Mux_v I__473 (
            .O(N__3580),
            .I(N__3566));
    InMux I__472 (
            .O(N__3579),
            .I(N__3563));
    Span4Mux_v I__471 (
            .O(N__3576),
            .I(N__3560));
    LocalMux I__470 (
            .O(N__3573),
            .I(N__3557));
    LocalMux I__469 (
            .O(N__3570),
            .I(N__3554));
    InMux I__468 (
            .O(N__3569),
            .I(N__3551));
    Sp12to4 I__467 (
            .O(N__3566),
            .I(N__3546));
    LocalMux I__466 (
            .O(N__3563),
            .I(N__3546));
    Span4Mux_h I__465 (
            .O(N__3560),
            .I(N__3539));
    Span4Mux_v I__464 (
            .O(N__3557),
            .I(N__3539));
    Span4Mux_v I__463 (
            .O(N__3554),
            .I(N__3539));
    LocalMux I__462 (
            .O(N__3551),
            .I(N__3536));
    Span12Mux_h I__461 (
            .O(N__3546),
            .I(N__3529));
    Sp12to4 I__460 (
            .O(N__3539),
            .I(N__3529));
    Span12Mux_v I__459 (
            .O(N__3536),
            .I(N__3529));
    Odrv12 I__458 (
            .O(N__3529),
            .I(A_c_20));
    CascadeMux I__457 (
            .O(N__3526),
            .I(N__3522));
    InMux I__456 (
            .O(N__3525),
            .I(N__3518));
    InMux I__455 (
            .O(N__3522),
            .I(N__3515));
    InMux I__454 (
            .O(N__3521),
            .I(N__3512));
    LocalMux I__453 (
            .O(N__3518),
            .I(N__3503));
    LocalMux I__452 (
            .O(N__3515),
            .I(N__3503));
    LocalMux I__451 (
            .O(N__3512),
            .I(N__3503));
    InMux I__450 (
            .O(N__3511),
            .I(N__3500));
    CascadeMux I__449 (
            .O(N__3510),
            .I(N__3495));
    Span4Mux_v I__448 (
            .O(N__3503),
            .I(N__3492));
    LocalMux I__447 (
            .O(N__3500),
            .I(N__3489));
    InMux I__446 (
            .O(N__3499),
            .I(N__3484));
    InMux I__445 (
            .O(N__3498),
            .I(N__3484));
    InMux I__444 (
            .O(N__3495),
            .I(N__3481));
    Span4Mux_v I__443 (
            .O(N__3492),
            .I(N__3478));
    Span4Mux_h I__442 (
            .O(N__3489),
            .I(N__3471));
    LocalMux I__441 (
            .O(N__3484),
            .I(N__3471));
    LocalMux I__440 (
            .O(N__3481),
            .I(N__3471));
    Span4Mux_v I__439 (
            .O(N__3478),
            .I(N__3468));
    Span4Mux_h I__438 (
            .O(N__3471),
            .I(N__3465));
    Sp12to4 I__437 (
            .O(N__3468),
            .I(N__3462));
    Sp12to4 I__436 (
            .O(N__3465),
            .I(N__3459));
    Span12Mux_h I__435 (
            .O(N__3462),
            .I(N__3454));
    Span12Mux_v I__434 (
            .O(N__3459),
            .I(N__3454));
    Odrv12 I__433 (
            .O(N__3454),
            .I(A_c_19));
    CascadeMux I__432 (
            .O(N__3451),
            .I(N__3448));
    InMux I__431 (
            .O(N__3448),
            .I(N__3442));
    InMux I__430 (
            .O(N__3447),
            .I(N__3442));
    LocalMux I__429 (
            .O(N__3442),
            .I(N__3438));
    InMux I__428 (
            .O(N__3441),
            .I(N__3435));
    Span4Mux_v I__427 (
            .O(N__3438),
            .I(N__3432));
    LocalMux I__426 (
            .O(N__3435),
            .I(N__3429));
    Span4Mux_h I__425 (
            .O(N__3432),
            .I(N__3423));
    Span4Mux_v I__424 (
            .O(N__3429),
            .I(N__3423));
    InMux I__423 (
            .O(N__3428),
            .I(N__3420));
    Sp12to4 I__422 (
            .O(N__3423),
            .I(N__3417));
    LocalMux I__421 (
            .O(N__3420),
            .I(N__3414));
    Span12Mux_s5_h I__420 (
            .O(N__3417),
            .I(N__3409));
    Span12Mux_v I__419 (
            .O(N__3414),
            .I(N__3409));
    Span12Mux_v I__418 (
            .O(N__3409),
            .I(N__3406));
    Odrv12 I__417 (
            .O(N__3406),
            .I(A_c_17));
    InMux I__416 (
            .O(N__3403),
            .I(N__3400));
    LocalMux I__415 (
            .O(N__3400),
            .I(N__3397));
    Span4Mux_v I__414 (
            .O(N__3397),
            .I(N__3393));
    InMux I__413 (
            .O(N__3396),
            .I(N__3390));
    Odrv4 I__412 (
            .O(N__3393),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_0 ));
    LocalMux I__411 (
            .O(N__3390),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_0 ));
    CascadeMux I__410 (
            .O(N__3385),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4_cascade_ ));
    CascadeMux I__409 (
            .O(N__3382),
            .I(N__3378));
    InMux I__408 (
            .O(N__3381),
            .I(N__3373));
    InMux I__407 (
            .O(N__3378),
            .I(N__3373));
    LocalMux I__406 (
            .O(N__3373),
            .I(N__3370));
    Span4Mux_h I__405 (
            .O(N__3370),
            .I(N__3367));
    Odrv4 I__404 (
            .O(N__3367),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_4 ));
    InMux I__403 (
            .O(N__3364),
            .I(N__3358));
    InMux I__402 (
            .O(N__3363),
            .I(N__3358));
    LocalMux I__401 (
            .O(N__3358),
            .I(N__3355));
    Span4Mux_v I__400 (
            .O(N__3355),
            .I(N__3352));
    Odrv4 I__399 (
            .O(N__3352),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_5 ));
    CascadeMux I__398 (
            .O(N__3349),
            .I(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_0_cascade_ ));
    InMux I__397 (
            .O(N__3346),
            .I(N__3343));
    LocalMux I__396 (
            .O(N__3343),
            .I(N__3340));
    Span4Mux_h I__395 (
            .O(N__3340),
            .I(N__3337));
    Span4Mux_v I__394 (
            .O(N__3337),
            .I(N__3334));
    Span4Mux_v I__393 (
            .O(N__3334),
            .I(N__3331));
    Odrv4 I__392 (
            .O(N__3331),
            .I(RnW_c));
    IoInMux I__391 (
            .O(N__3328),
            .I(N__3325));
    LocalMux I__390 (
            .O(N__3325),
            .I(N__3319));
    IoInMux I__389 (
            .O(N__3324),
            .I(N__3316));
    IoInMux I__388 (
            .O(N__3323),
            .I(N__3313));
    IoInMux I__387 (
            .O(N__3322),
            .I(N__3310));
    IoSpan4Mux I__386 (
            .O(N__3319),
            .I(N__3300));
    LocalMux I__385 (
            .O(N__3316),
            .I(N__3300));
    LocalMux I__384 (
            .O(N__3313),
            .I(N__3300));
    LocalMux I__383 (
            .O(N__3310),
            .I(N__3297));
    IoInMux I__382 (
            .O(N__3309),
            .I(N__3294));
    IoInMux I__381 (
            .O(N__3308),
            .I(N__3291));
    IoInMux I__380 (
            .O(N__3307),
            .I(N__3288));
    IoSpan4Mux I__379 (
            .O(N__3300),
            .I(N__3281));
    IoSpan4Mux I__378 (
            .O(N__3297),
            .I(N__3281));
    LocalMux I__377 (
            .O(N__3294),
            .I(N__3281));
    LocalMux I__376 (
            .O(N__3291),
            .I(N__3276));
    LocalMux I__375 (
            .O(N__3288),
            .I(N__3276));
    IoSpan4Mux I__374 (
            .O(N__3281),
            .I(N__3270));
    IoSpan4Mux I__373 (
            .O(N__3276),
            .I(N__3270));
    IoInMux I__372 (
            .O(N__3275),
            .I(N__3267));
    Sp12to4 I__371 (
            .O(N__3270),
            .I(N__3262));
    LocalMux I__370 (
            .O(N__3267),
            .I(N__3262));
    Span12Mux_s3_v I__369 (
            .O(N__3262),
            .I(N__3259));
    Span12Mux_v I__368 (
            .O(N__3259),
            .I(N__3256));
    Odrv12 I__367 (
            .O(N__3256),
            .I(D_1_i));
    IoInMux I__366 (
            .O(N__3253),
            .I(N__3250));
    LocalMux I__365 (
            .O(N__3250),
            .I(N__3247));
    IoSpan4Mux I__364 (
            .O(N__3247),
            .I(N__3244));
    Span4Mux_s2_h I__363 (
            .O(N__3244),
            .I(N__3241));
    Sp12to4 I__362 (
            .O(N__3241),
            .I(N__3238));
    Span12Mux_s11_h I__361 (
            .O(N__3238),
            .I(N__3235));
    Span12Mux_h I__360 (
            .O(N__3235),
            .I(N__3232));
    Span12Mux_v I__359 (
            .O(N__3232),
            .I(N__3229));
    Odrv12 I__358 (
            .O(N__3229),
            .I(U409_ADDRESS_DECODE_un1_RTC_ENn_i));
    InMux I__357 (
            .O(N__3226),
            .I(N__3223));
    LocalMux I__356 (
            .O(N__3223),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3 ));
    CascadeMux I__355 (
            .O(N__3220),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3_cascade_ ));
    InMux I__354 (
            .O(N__3217),
            .I(N__3214));
    LocalMux I__353 (
            .O(N__3214),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_0 ));
    InMux I__352 (
            .O(N__3211),
            .I(N__3208));
    LocalMux I__351 (
            .O(N__3208),
            .I(N__3205));
    Span4Mux_v I__350 (
            .O(N__3205),
            .I(N__3202));
    Odrv4 I__349 (
            .O(N__3202),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_5 ));
    CascadeMux I__348 (
            .O(N__3199),
            .I(U409_ADDRESS_DECODE_LOWROM_3_cascade_));
    InMux I__347 (
            .O(N__3196),
            .I(N__3193));
    LocalMux I__346 (
            .O(N__3193),
            .I(N__3190));
    Odrv4 I__345 (
            .O(N__3190),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_3 ));
    CascadeMux I__344 (
            .O(N__3187),
            .I(N__3184));
    InMux I__343 (
            .O(N__3184),
            .I(N__3181));
    LocalMux I__342 (
            .O(N__3181),
            .I(N__3178));
    Span4Mux_v I__341 (
            .O(N__3178),
            .I(N__3175));
    Odrv4 I__340 (
            .O(N__3175),
            .I(U409_ADDRESS_DECODE_AUTOVECTOR_3));
    InMux I__339 (
            .O(N__3172),
            .I(N__3169));
    LocalMux I__338 (
            .O(N__3169),
            .I(N__3166));
    Odrv4 I__337 (
            .O(N__3166),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5 ));
    CascadeMux I__336 (
            .O(N__3163),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_ ));
    InMux I__335 (
            .O(N__3160),
            .I(N__3154));
    InMux I__334 (
            .O(N__3159),
            .I(N__3154));
    LocalMux I__333 (
            .O(N__3154),
            .I(N__3151));
    Span4Mux_v I__332 (
            .O(N__3151),
            .I(N__3148));
    Sp12to4 I__331 (
            .O(N__3148),
            .I(N__3145));
    Odrv12 I__330 (
            .O(N__3145),
            .I(A_c_31));
    InMux I__329 (
            .O(N__3142),
            .I(N__3136));
    InMux I__328 (
            .O(N__3141),
            .I(N__3136));
    LocalMux I__327 (
            .O(N__3136),
            .I(N__3133));
    Span4Mux_v I__326 (
            .O(N__3133),
            .I(N__3130));
    Span4Mux_h I__325 (
            .O(N__3130),
            .I(N__3127));
    Odrv4 I__324 (
            .O(N__3127),
            .I(A_c_30));
    CascadeMux I__323 (
            .O(N__3124),
            .I(N__3120));
    InMux I__322 (
            .O(N__3123),
            .I(N__3115));
    InMux I__321 (
            .O(N__3120),
            .I(N__3115));
    LocalMux I__320 (
            .O(N__3115),
            .I(N__3112));
    Span4Mux_v I__319 (
            .O(N__3112),
            .I(N__3109));
    Span4Mux_v I__318 (
            .O(N__3109),
            .I(N__3106));
    Sp12to4 I__317 (
            .O(N__3106),
            .I(N__3103));
    Odrv12 I__316 (
            .O(N__3103),
            .I(A_c_28));
    InMux I__315 (
            .O(N__3100),
            .I(N__3094));
    InMux I__314 (
            .O(N__3099),
            .I(N__3094));
    LocalMux I__313 (
            .O(N__3094),
            .I(N__3091));
    Span4Mux_h I__312 (
            .O(N__3091),
            .I(N__3088));
    Span4Mux_v I__311 (
            .O(N__3088),
            .I(N__3085));
    Odrv4 I__310 (
            .O(N__3085),
            .I(A_c_29));
    CascadeMux I__309 (
            .O(N__3082),
            .I(\U409_ADDRESS_DECODE.CIA_SPACE_0Z0Z_1_cascade_ ));
    CascadeMux I__308 (
            .O(N__3079),
            .I(N__3076));
    InMux I__307 (
            .O(N__3076),
            .I(N__3072));
    InMux I__306 (
            .O(N__3075),
            .I(N__3069));
    LocalMux I__305 (
            .O(N__3072),
            .I(N__3064));
    LocalMux I__304 (
            .O(N__3069),
            .I(N__3064));
    Span4Mux_h I__303 (
            .O(N__3064),
            .I(N__3061));
    Span4Mux_v I__302 (
            .O(N__3061),
            .I(N__3058));
    Sp12to4 I__301 (
            .O(N__3058),
            .I(N__3055));
    Span12Mux_v I__300 (
            .O(N__3055),
            .I(N__3052));
    Odrv12 I__299 (
            .O(N__3052),
            .I(A_c_16));
    CascadeMux I__298 (
            .O(N__3049),
            .I(\U409_ADDRESS_DECODE.RAN_SPACEZ0Z_0_cascade_ ));
    CascadeMux I__297 (
            .O(N__3046),
            .I(N__3043));
    InMux I__296 (
            .O(N__3043),
            .I(N__3037));
    InMux I__295 (
            .O(N__3042),
            .I(N__3037));
    LocalMux I__294 (
            .O(N__3037),
            .I(N__3034));
    Span4Mux_v I__293 (
            .O(N__3034),
            .I(N__3031));
    Span4Mux_h I__292 (
            .O(N__3031),
            .I(N__3028));
    Odrv4 I__291 (
            .O(N__3028),
            .I(A_c_27));
    CascadeMux I__290 (
            .O(N__3025),
            .I(N__3021));
    InMux I__289 (
            .O(N__3024),
            .I(N__3016));
    InMux I__288 (
            .O(N__3021),
            .I(N__3016));
    LocalMux I__287 (
            .O(N__3016),
            .I(N__3013));
    Span4Mux_v I__286 (
            .O(N__3013),
            .I(N__3010));
    Span4Mux_v I__285 (
            .O(N__3010),
            .I(N__3007));
    Sp12to4 I__284 (
            .O(N__3007),
            .I(N__3004));
    Odrv12 I__283 (
            .O(N__3004),
            .I(A_c_26));
    InMux I__282 (
            .O(N__3001),
            .I(N__2995));
    InMux I__281 (
            .O(N__3000),
            .I(N__2995));
    LocalMux I__280 (
            .O(N__2995),
            .I(N__2992));
    Span4Mux_v I__279 (
            .O(N__2992),
            .I(N__2989));
    Sp12to4 I__278 (
            .O(N__2989),
            .I(N__2986));
    Odrv12 I__277 (
            .O(N__2986),
            .I(A_c_25));
    InMux I__276 (
            .O(N__2983),
            .I(N__2980));
    LocalMux I__275 (
            .O(N__2980),
            .I(N__2976));
    InMux I__274 (
            .O(N__2979),
            .I(N__2973));
    Span4Mux_v I__273 (
            .O(N__2976),
            .I(N__2968));
    LocalMux I__272 (
            .O(N__2973),
            .I(N__2968));
    Span4Mux_h I__271 (
            .O(N__2968),
            .I(N__2965));
    Span4Mux_v I__270 (
            .O(N__2965),
            .I(N__2962));
    Odrv4 I__269 (
            .O(N__2962),
            .I(A_c_24));
    ClkMux I__268 (
            .O(N__2959),
            .I(N__2920));
    ClkMux I__267 (
            .O(N__2958),
            .I(N__2920));
    ClkMux I__266 (
            .O(N__2957),
            .I(N__2920));
    ClkMux I__265 (
            .O(N__2956),
            .I(N__2920));
    ClkMux I__264 (
            .O(N__2955),
            .I(N__2920));
    ClkMux I__263 (
            .O(N__2954),
            .I(N__2920));
    ClkMux I__262 (
            .O(N__2953),
            .I(N__2920));
    ClkMux I__261 (
            .O(N__2952),
            .I(N__2920));
    ClkMux I__260 (
            .O(N__2951),
            .I(N__2920));
    ClkMux I__259 (
            .O(N__2950),
            .I(N__2920));
    ClkMux I__258 (
            .O(N__2949),
            .I(N__2920));
    ClkMux I__257 (
            .O(N__2948),
            .I(N__2920));
    ClkMux I__256 (
            .O(N__2947),
            .I(N__2920));
    GlobalMux I__255 (
            .O(N__2920),
            .I(CLK80_OUT));
    INV \INVU409_TRANSFER_ACK.LASTCLK_0C  (
            .O(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .I(N__2957));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_1C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .I(N__2951));
    INV \INVU409_TRANSFER_ACK.CIA_ENABLED_1C  (
            .O(\INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ),
            .I(N__2948));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .I(N__2947));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .I(N__2950));
    INV \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC  (
            .O(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .I(N__2958));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .I(N__2953));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net ),
            .I(N__2949));
    INV \INVU409_TRANSFER_ACK.IRQ_TACK_EN_nesrC  (
            .O(\INVU409_TRANSFER_ACK.IRQ_TACK_EN_nesrC_net ),
            .I(N__2959));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net ),
            .I(N__2956));
    INV \INVU409_TRANSFER_ACK.TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.TACK_ENC_net ),
            .I(N__2955));
    INV \INVU409_TRANSFER_ACK.TACK_OUTnC  (
            .O(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .I(N__2954));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_EN_nerC  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_EN_nerC_net ),
            .I(N__2952));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_9_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_14_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_9_0_));
    defparam IN_MUX_bfv_14_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_10_0_ (
            .carryinitin(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .carryinitout(bfn_14_10_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_11_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_1_15_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_1_15_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_1_15_2  (
            .in0(N__3001),
            .in1(N__3024),
            .in2(N__3046),
            .in3(N__6207),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_4_LC_1_15_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_4_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_4_LC_1_15_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_4_LC_1_15_5  (
            .in0(N__2983),
            .in1(N__3042),
            .in2(N__3025),
            .in3(N__3000),
            .lcout(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_1  (
            .in0(N__3160),
            .in1(N__3142),
            .in2(_gnd_net_),
            .in3(N__2979),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_2  (
            .in0(N__3100),
            .in1(N__3172),
            .in2(N__3163),
            .in3(N__3123),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_5_LC_1_17_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_5_LC_1_17_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_5_LC_1_17_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_5_LC_1_17_5  (
            .in0(N__3159),
            .in1(N__3141),
            .in2(N__3124),
            .in3(N__3099),
            .lcout(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_0_1_LC_2_13_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_0_1_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_0_1_LC_2_13_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_0_1_LC_2_13_3  (
            .in0(N__4424),
            .in1(N__3569),
            .in2(N__3510),
            .in3(N__3645),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.CIA_SPACE_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_0_LC_2_13_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_0_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_0_LC_2_13_4 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_0_LC_2_13_4  (
            .in0(N__3075),
            .in1(_gnd_net_),
            .in2(N__3082),
            .in3(N__3428),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_5_LC_3_13_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_5_LC_3_13_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_5_LC_3_13_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_5_LC_3_13_1  (
            .in0(N__3498),
            .in1(N__3646),
            .in2(N__3079),
            .in3(N__3441),
            .lcout(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.RAN_SPACE_0_LC_3_13_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.RAN_SPACE_0_LC_3_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.RAN_SPACE_0_LC_3_13_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U409_ADDRESS_DECODE.RAN_SPACE_0_LC_3_13_4  (
            .in0(N__3953),
            .in1(N__4425),
            .in2(_gnd_net_),
            .in3(N__4012),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.RAN_SPACEZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_0_LC_3_13_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_0_LC_3_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_0_LC_3_13_5 .LUT_INIT=16'b1110111111001111;
    LogicCell40 \U409_ADDRESS_DECODE.un2_REGSPACEn_0_LC_3_13_5  (
            .in0(N__3499),
            .in1(N__3583),
            .in2(N__3049),
            .in3(N__3647),
            .lcout(\U409_ADDRESS_DECODE.un2_REGSPACEn_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_3_LC_3_14_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_3_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_3_LC_3_14_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_3_LC_3_14_2  (
            .in0(N__4389),
            .in1(N__3584),
            .in2(N__3382),
            .in3(N__3363),
            .lcout(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_0_LC_3_14_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_0_LC_3_14_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_0_LC_3_14_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_0_LC_3_14_3  (
            .in0(N__3396),
            .in1(N__3989),
            .in2(_gnd_net_),
            .in3(N__3943),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_3_LC_3_14_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_3_LC_3_14_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_3_LC_3_14_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_3_LC_3_14_4  (
            .in0(N__3381),
            .in1(N__3364),
            .in2(N__3349),
            .in3(N__6242),
            .lcout(U409_ADDRESS_DECODE_AUTOVECTOR_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.D_1_i_LC_3_16_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.D_1_i_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.D_1_i_LC_3_16_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \U409_AUTOCONFIG.D_1_i_LC_3_16_6  (
            .in0(N__3346),
            .in1(N__6326),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(D_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_5_13_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_5_13_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_5_13_2  (
            .in0(N__3941),
            .in1(N__3598),
            .in2(N__3673),
            .in3(N__3226),
            .lcout(U409_ADDRESS_DECODE_un1_RTC_ENn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_3_LC_5_13_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_3_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_3_LC_5_13_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_3_LC_5_13_5  (
            .in0(N__3511),
            .in1(N__4437),
            .in2(N__3655),
            .in3(N__3854),
            .lcout(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3 ),
            .ltout(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_5_13_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_5_13_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_5_13_6  (
            .in0(N__3940),
            .in1(N__3597),
            .in2(N__3220),
            .in3(N__3666),
            .lcout(U409_ADDRESS_DECODE_un1_RTC_ENn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_LC_5_14_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_LC_5_14_2 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_LC_5_14_2  (
            .in0(N__4045),
            .in1(N__4081),
            .in2(_gnd_net_),
            .in3(N__6243),
            .lcout(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_9_0_a2_LC_5_14_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_9_0_a2_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_9_0_a2_LC_5_14_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_9_0_a2_LC_5_14_5  (
            .in0(_gnd_net_),
            .in1(N__3993),
            .in2(_gnd_net_),
            .in3(N__3954),
            .lcout(U409_ADDRESS_DECODE_LOWROM_3),
            .ltout(U409_ADDRESS_DECODE_LOWROM_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_5_14_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_5_14_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_5_14_6  (
            .in0(N__3217),
            .in1(N__3211),
            .in2(N__3199),
            .in3(N__3196),
            .lcout(AUTOCONFIG_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_LC_5_15_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_LC_5_15_3 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_LC_5_15_3  (
            .in0(N__6244),
            .in1(N__3765),
            .in2(N__3187),
            .in3(N__3694),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_2_LC_5_20_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_2_LC_5_20_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_2_LC_5_20_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_2_LC_5_20_1  (
            .in0(_gnd_net_),
            .in1(N__3724),
            .in2(_gnd_net_),
            .in3(N__3709),
            .lcout(U409_ADDRESS_DECODE_AUTOVECTOR_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_8_0_a2_LC_6_12_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_8_0_a2_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_8_0_a2_LC_6_12_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_8_0_a2_LC_6_12_4  (
            .in0(_gnd_net_),
            .in1(N__4439),
            .in2(_gnd_net_),
            .in3(N__3579),
            .lcout(),
            .ltout(U409_ADDRESS_DECODE_LOWROM_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_LC_6_12_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_LC_6_12_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_LC_6_12_5  (
            .in0(N__3521),
            .in1(N__4308),
            .in2(N__3685),
            .in3(N__4363),
            .lcout(\U409_TRANSFER_ACK.N_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2_1_LC_6_13_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2_1_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2_1_LC_6_13_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2_1_LC_6_13_1  (
            .in0(N__3596),
            .in1(N__4438),
            .in2(_gnd_net_),
            .in3(N__3942),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_6_13_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_6_13_2 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_6_13_2  (
            .in0(N__3682),
            .in1(N__3525),
            .in2(N__3676),
            .in3(N__4015),
            .lcout(\U409_TRANSFER_ACK.N_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_2_LC_6_13_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_2_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_2_LC_6_13_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_2_LC_6_13_3  (
            .in0(N__4014),
            .in1(N__4084),
            .in2(N__3451),
            .in3(N__4051),
            .lcout(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.REG_SPACE_3_LC_6_13_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.REG_SPACE_3_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.REG_SPACE_3_LC_6_13_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.REG_SPACE_3_LC_6_13_4  (
            .in0(N__3654),
            .in1(N__3595),
            .in2(N__3526),
            .in3(N__3447),
            .lcout(\U409_ADDRESS_DECODE.REG_SPACE_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_14_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_14_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_14_1  (
            .in0(N__4046),
            .in1(N__4082),
            .in2(_gnd_net_),
            .in3(N__3994),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_14_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_14_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_14_2  (
            .in0(N__3403),
            .in1(N__3855),
            .in2(N__3385),
            .in3(N__3955),
            .lcout(CIA_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_1_LC_6_14_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_1_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_1_LC_6_14_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_1_LC_6_14_6  (
            .in0(N__4083),
            .in1(N__3856),
            .in2(_gnd_net_),
            .in3(N__4047),
            .lcout(U409_ADDRESS_DECODE_ROMEN_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.REG_SPACE_2_LC_6_15_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.REG_SPACE_2_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.REG_SPACE_2_LC_6_15_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U409_ADDRESS_DECODE.REG_SPACE_2_LC_6_15_6  (
            .in0(N__4423),
            .in1(N__4013),
            .in2(_gnd_net_),
            .in3(N__3920),
            .lcout(\U409_ADDRESS_DECODE.REG_SPACEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_16_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_16_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_16_2 .LUT_INIT=16'b0111000011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_16_2  (
            .in0(N__3778),
            .in1(N__3792),
            .in2(N__3811),
            .in3(N__3853),
            .lcout(U409_ADDRESS_DECODE_un1_REGSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_16_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_16_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_16_7 .LUT_INIT=16'b1010001000100010;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_16_7  (
            .in0(N__3852),
            .in1(N__3807),
            .in2(N__3793),
            .in3(N__3777),
            .lcout(U409_ADDRESS_DECODE_un1_REGSPACEn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_16_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_16_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_16_7  (
            .in0(N__3769),
            .in1(N__5402),
            .in2(_gnd_net_),
            .in3(N__6803),
            .lcout(PORTSIZE_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_2_LC_8_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_2_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_2_LC_8_9_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_2_LC_8_9_2  (
            .in0(N__4830),
            .in1(N__5251),
            .in2(N__4788),
            .in3(N__5150),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_8_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_8_9_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_8_9_3  (
            .in0(N__4668),
            .in1(N__5215),
            .in2(N__3739),
            .in3(N__5317),
            .lcout(\U409_TRANSFER_ACK.N_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_LC_9_6_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_LC_9_6_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_LC_9_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_LC_9_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4612),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_EN_nerC_net ),
            .ce(N__3736),
            .sr(N__4747));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_sbtinv_LC_9_7_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_sbtinv_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_sbtinv_LC_9_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_sbtinv_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4267),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_RNIIFHQ_LC_9_7_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_RNIIFHQ_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_RNIIFHQ_LC_9_7_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_RNIIFHQ_LC_9_7_2  (
            .in0(N__4276),
            .in1(N__4255),
            .in2(N__4294),
            .in3(N__4095),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER6 ),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_9_7_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_9_7_3 .LUT_INIT=16'b0000000111011101;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_9_7_3  (
            .in0(N__4180),
            .in1(N__4159),
            .in2(N__4249),
            .in3(N__4204),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_9_7_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_9_7_4 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_LC_9_7_4  (
            .in0(N__6212),
            .in1(_gnd_net_),
            .in2(N__4246),
            .in3(N__4205),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_9_7_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_9_7_5 .LUT_INIT=16'b0000100000001100;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_9_7_5  (
            .in0(N__4182),
            .in1(N__6208),
            .in2(N__4165),
            .in3(N__4140),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_9_7_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_9_7_6 .LUT_INIT=16'b0101000010100000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_9_7_6  (
            .in0(N__4160),
            .in1(_gnd_net_),
            .in2(N__6225),
            .in3(N__4181),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_7_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_7_7 .LUT_INIT=16'b1101110111101110;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_7_7  (
            .in0(N__5163),
            .in1(N__5305),
            .in2(_gnd_net_),
            .in3(N__5269),
            .lcout(\U409_TRANSFER_ACK.N_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_9_8_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_9_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_9_8_0 .LUT_INIT=16'b0111000001110001;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_LC_9_8_0  (
            .in0(N__4183),
            .in1(N__4161),
            .in2(N__6353),
            .in3(N__4141),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_ENC_net ),
            .ce(),
            .sr(N__6451));
    defparam \U409_TRANSFER_ACK.ROMENn_LC_9_8_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_9_8_3 .SEQ_MODE=4'b1001;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_9_8_3 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_LC_9_8_3  (
            .in0(N__4107),
            .in1(N__5125),
            .in2(_gnd_net_),
            .in3(N__4129),
            .lcout(ROMENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_ENC_net ),
            .ce(),
            .sr(N__6451));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_9_8_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_9_8_6 .LUT_INIT=16'b0011010100100000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_LC_9_8_6  (
            .in0(N__4576),
            .in1(N__5629),
            .in2(N__5701),
            .in3(N__4096),
            .lcout(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_ENC_net ),
            .ce(),
            .sr(N__6451));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_9_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_9_9_0 .LUT_INIT=16'b0111100011010000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_9_9_0  (
            .in0(N__5161),
            .in1(N__5219),
            .in2(N__5274),
            .in3(N__5319),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net ),
            .ce(),
            .sr(N__6434));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_9_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_9_9_3 .LUT_INIT=16'b1101111100000010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_LC_9_9_3  (
            .in0(N__4585),
            .in1(N__5320),
            .in2(N__5224),
            .in3(N__4290),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net ),
            .ce(),
            .sr(N__6434));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_9_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_9_9_7 .LUT_INIT=16'b0101101110100000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_9_9_7  (
            .in0(N__5318),
            .in1(N__5264),
            .in2(N__5223),
            .in3(N__5160),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net ),
            .ce(),
            .sr(N__6434));
    defparam RESETn_ibuf_RNIM9SF_LC_9_10_6.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_9_10_6.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_9_10_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_9_10_6 (
            .in0(N__6226),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_LC_9_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_LC_9_11_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_LC_9_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4498),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_EN_nesrC_net ),
            .ce(N__4480),
            .sr(N__6446));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI8JGQ6_4_LC_10_6_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI8JGQ6_4_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI8JGQ6_4_LC_10_6_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI8JGQ6_4_LC_10_6_1  (
            .in0(_gnd_net_),
            .in1(N__4623),
            .in2(_gnd_net_),
            .in3(N__4642),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23 ),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIEEVK7_0_LC_10_6_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIEEVK7_0_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIEEVK7_0_LC_10_6_2 .LUT_INIT=16'b0000111100000010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIEEVK7_0_LC_10_6_2  (
            .in0(N__5541),
            .in1(N__4555),
            .in2(N__4261),
            .in3(N__4996),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_6_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_6_3 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_6_3 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_6_3  (
            .in0(_gnd_net_),
            .in1(N__4924),
            .in2(N__4258),
            .in3(N__4897),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net ),
            .ce(),
            .sr(N__4746));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_7_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_7_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_7_0 .LUT_INIT=16'b0001000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_7_0  (
            .in0(N__4554),
            .in1(N__4997),
            .in2(N__5547),
            .in3(N__4624),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__4739));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_10_7_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_10_7_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_10_7_5  (
            .in0(_gnd_net_),
            .in1(N__5268),
            .in2(_gnd_net_),
            .in3(N__5162),
            .lcout(\U409_TRANSFER_ACK.N_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_10_8_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_10_8_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_10_8_4  (
            .in0(N__5697),
            .in1(N__6475),
            .in2(N__5546),
            .in3(N__6505),
            .lcout(\U409_TRANSFER_ACK.N_142 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER16_LC_10_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER16_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER16_LC_10_9_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER16_LC_10_9_1  (
            .in0(N__4532),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5496),
            .lcout(\U409_TRANSFER_ACK.N_35_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_11_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_11_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_11_0  (
            .in0(N__4497),
            .in1(N__4569),
            .in2(N__5542),
            .in3(N__4543),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNIBIO4C_LC_10_11_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNIBIO4C_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNIBIO4C_LC_10_11_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNIBIO4C_LC_10_11_3  (
            .in0(N__4570),
            .in1(N__5527),
            .in2(N__4553),
            .in3(N__4496),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_RNO_LC_10_11_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_RNO_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_RNO_LC_10_11_4 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_RNO_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4483),
            .in3(N__6408),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_10_12_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_10_12_7 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_10_12_7  (
            .in0(N__4321),
            .in1(N__4447),
            .in2(N__4829),
            .in3(N__4355),
            .lcout(U409_ADDRESS_DECODE_un1_RAMSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_10_13_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_10_13_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_10_13_0  (
            .in0(N__4811),
            .in1(N__4446),
            .in2(N__4362),
            .in3(N__4320),
            .lcout(U409_ADDRESS_DECODE_un1_RAMSPACEn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI1CKM1_5_LC_11_6_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI1CKM1_5_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI1CKM1_5_LC_11_6_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI1CKM1_5_LC_11_6_0  (
            .in0(N__4604),
            .in1(N__5026),
            .in2(N__5058),
            .in3(N__4890),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_4_LC_11_6_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_4_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_4_LC_11_6_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_4_LC_11_6_1  (
            .in0(N__4994),
            .in1(N__4861),
            .in2(N__4645),
            .in3(N__4636),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_6_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_6_2 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_6_2  (
            .in0(N__4961),
            .in1(N__4942),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_5_LC_11_6_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_5_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_5_LC_11_6_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_5_LC_11_6_5  (
            .in0(N__5027),
            .in1(N__4603),
            .in2(N__5059),
            .in3(N__4860),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_11_6_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_11_6_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_11_6_6  (
            .in0(N__4635),
            .in1(N__4993),
            .in2(N__4627),
            .in3(N__4891),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_7_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_7_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_7_0 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_7_0  (
            .in0(N__5057),
            .in1(N__4608),
            .in2(N__5089),
            .in3(N__5008),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .ce(),
            .sr(N__4721));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_7_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_7_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_7_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_7_1  (
            .in0(N__4840),
            .in1(N__5029),
            .in2(_gnd_net_),
            .in3(N__5073),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .ce(),
            .sr(N__4721));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_7_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_7_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_7_2 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_7_2  (
            .in0(N__4998),
            .in1(_gnd_net_),
            .in2(N__5087),
            .in3(N__4945),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .ce(),
            .sr(N__4721));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_7_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_7_3 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_7_3 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_7_3  (
            .in0(N__4944),
            .in1(N__4999),
            .in2(_gnd_net_),
            .in3(N__4963),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .ce(),
            .sr(N__4721));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_7_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_7_4 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_7_4 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_7_4  (
            .in0(N__4922),
            .in1(N__4898),
            .in2(N__5088),
            .in3(N__4864),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .ce(),
            .sr(N__4721));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_7_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_7_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_7_6 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(N__5007),
            .in2(N__5086),
            .in3(N__5056),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .ce(),
            .sr(N__4721));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_8_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_8_0  (
            .in0(N__4899),
            .in1(N__5028),
            .in2(N__4923),
            .in3(N__4862),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_11_8_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_11_8_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_11_8_5  (
            .in0(N__4995),
            .in1(N__4962),
            .in2(_gnd_net_),
            .in3(N__4943),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_11_8_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_11_8_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_11_8_6  (
            .in0(N__4900),
            .in1(_gnd_net_),
            .in2(N__4867),
            .in3(N__4863),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_1_0_LC_11_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_1_0_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_1_0_LC_11_9_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_1_0_LC_11_9_0  (
            .in0(N__5214),
            .in1(N__4834),
            .in2(N__4792),
            .in3(N__5273),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_11_16_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_11_16_7 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_11_16_7  (
            .in0(N__5409),
            .in1(N__5427),
            .in2(N__6232),
            .in3(N__4765),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_1_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_1_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_1_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_1_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_7_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_7_3 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_7_3  (
            .in0(N__5202),
            .in1(N__4684),
            .in2(N__4675),
            .in3(N__4654),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__6442));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_7_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_7_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_7_4  (
            .in0(_gnd_net_),
            .in1(N__5201),
            .in2(_gnd_net_),
            .in3(N__5304),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__6442));
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_12_8_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_12_8_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_TICK.COUNTER60_RNIHJU51_4_LC_12_8_0  (
            .in0(N__5111),
            .in1(N__5962),
            .in2(_gnd_net_),
            .in3(N__5362),
            .lcout(\U409_TICK.TICK603_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_1_LC_12_8_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_1_LC_12_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_1_LC_12_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER60_1_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(N__5112),
            .in2(_gnd_net_),
            .in3(N__6038),
            .lcout(\U409_TICK.COUNTER60Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6878),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_0_LC_12_8_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_0_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_0_LC_12_8_2 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U409_TICK.COUNTER60_0_LC_12_8_2  (
            .in0(N__5840),
            .in1(N__5801),
            .in2(N__5116),
            .in3(N__5767),
            .lcout(\U409_TICK.COUNTER60Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6878),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_8_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_8_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_8_4  (
            .in0(N__5303),
            .in1(N__5275),
            .in2(N__5213),
            .in3(N__5167),
            .lcout(\U409_TRANSFER_ACK.N_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_8_LC_12_8_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_8_LC_12_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_8_LC_12_8_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_8_LC_12_8_7  (
            .in0(N__5766),
            .in1(N__5841),
            .in2(N__5808),
            .in3(N__5341),
            .lcout(\U409_TICK.COUNTER60Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6878),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_12_9_0 .C_ON=1'b1;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_12_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__5110),
            .in2(N__6039),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_2_LC_12_9_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_2_LC_12_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_2_LC_12_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_2_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(N__6051),
            .in2(_gnd_net_),
            .in3(N__5095),
            .lcout(\U409_TICK.COUNTER60Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .clk(N__6881),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_3_LC_12_9_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_3_LC_12_9_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_3_LC_12_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_3_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__5982),
            .in2(_gnd_net_),
            .in3(N__5092),
            .lcout(\U409_TICK.COUNTER60Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .clk(N__6881),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_12_9_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_12_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_4_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(N__5961),
            .in2(_gnd_net_),
            .in3(N__5365),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_5_LC_12_9_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_5_LC_12_9_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_5_LC_12_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_5_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(N__5361),
            .in2(_gnd_net_),
            .in3(N__5350),
            .lcout(\U409_TICK.COUNTER60Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .clk(N__6881),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_12_9_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_12_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_6_LC_12_9_5  (
            .in0(_gnd_net_),
            .in1(N__5934),
            .in2(_gnd_net_),
            .in3(N__5347),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_7_LC_12_9_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_7_LC_12_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_7_LC_12_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_7_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(N__5874),
            .in2(_gnd_net_),
            .in3(N__5344),
            .lcout(\U409_TICK.COUNTER60Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .clk(N__6881),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_12_9_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_12_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_8_LC_12_9_7  (
            .in0(_gnd_net_),
            .in1(N__5949),
            .in2(_gnd_net_),
            .in3(N__5335),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_12_10_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_12_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_9_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__5712),
            .in2(_gnd_net_),
            .in3(N__5332),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_10_LC_12_10_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_10_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_10_LC_12_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_10_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(N__5889),
            .in2(_gnd_net_),
            .in3(N__5329),
            .lcout(\U409_TICK.COUNTER60Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .clk(N__6884),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_11_LC_12_10_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_11_LC_12_10_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_11_LC_12_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_11_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(N__6003),
            .in2(_gnd_net_),
            .in3(N__5326),
            .lcout(\U409_TICK.COUNTER60Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .clk(N__6884),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_12_LC_12_10_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_12_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_12_LC_12_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_12_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__6063),
            .in2(_gnd_net_),
            .in3(N__5323),
            .lcout(\U409_TICK.COUNTER60Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .clk(N__6884),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_13_LC_12_10_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_13_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_13_LC_12_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_13_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(N__5902),
            .in2(_gnd_net_),
            .in3(N__5440),
            .lcout(\U409_TICK.COUNTER60Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .clk(N__6884),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_12_10_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_12_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_14_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(N__5913),
            .in2(_gnd_net_),
            .in3(N__5437),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_12_10_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_12_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_15_LC_12_10_6  (
            .in0(_gnd_net_),
            .in1(N__5853),
            .in2(_gnd_net_),
            .in3(N__5434),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_16_LC_12_10_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_16_LC_12_10_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_16_LC_12_10_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER60_16_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(N__6016),
            .in2(_gnd_net_),
            .in3(N__5431),
            .lcout(\U409_TICK.COUNTER60Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6884),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_DATA_BUFFERS.un1_BUFENn_LC_12_16_4 .C_ON=1'b0;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_LC_12_16_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_DATA_BUFFERS.un1_BUFENn_LC_12_16_4  (
            .in0(N__5428),
            .in1(N__6333),
            .in2(_gnd_net_),
            .in3(N__5410),
            .lcout(BUFENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_13_6_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_13_6_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_13_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_13_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5577),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ),
            .ce(),
            .sr(N__6450));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_13_6_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_13_6_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_13_6_6  (
            .in0(N__6775),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6186),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ),
            .ce(),
            .sr(N__6450));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_13_7_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_13_7_0 .LUT_INIT=16'b0001000000011111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_13_7_0  (
            .in0(N__5575),
            .in1(N__5598),
            .in2(N__5696),
            .in3(N__5635),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.i6_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_13_7_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_13_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_13_7_1 .LUT_INIT=16'b0100110000001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_1_LC_13_7_1  (
            .in0(N__5621),
            .in1(N__6188),
            .in2(N__5368),
            .in3(N__5689),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_LC_13_7_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_LC_13_7_5 .LUT_INIT=16'b0001000000011111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_LC_13_7_5  (
            .in0(N__5599),
            .in1(N__5576),
            .in2(N__5625),
            .in3(N__5452),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.N_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_13_7_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_13_7_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_13_7_6 .LUT_INIT=16'b0100110000001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_0_LC_13_7_6  (
            .in0(N__5688),
            .in1(N__6187),
            .in2(N__5665),
            .in3(N__5554),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK60_LC_13_8_1 .C_ON=1'b0;
    defparam \U409_TICK.TICK60_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK60_LC_13_8_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK60_LC_13_8_1  (
            .in0(N__5765),
            .in1(N__5646),
            .in2(N__5809),
            .in3(N__5842),
            .lcout(TICK60_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6876),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_1_LC_13_8_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_1_LC_13_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_1_LC_13_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER50_1_LC_13_8_2  (
            .in0(_gnd_net_),
            .in1(N__6580),
            .in2(_gnd_net_),
            .in3(N__6558),
            .lcout(\U409_TICK.COUNTER50Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6876),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_13_8_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_13_8_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_13_8_5  (
            .in0(_gnd_net_),
            .in1(N__6470),
            .in2(_gnd_net_),
            .in3(N__6500),
            .lcout(\U409_TRANSFER_ACK.N_4 ),
            .ltout(\U409_TRANSFER_ACK.N_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m4_LC_13_8_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m4_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m4_LC_13_8_6 .LUT_INIT=16'b0100111000001010;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m4_LC_13_8_6  (
            .in0(N__5617),
            .in1(N__5597),
            .in2(N__5581),
            .in3(N__5578),
            .lcout(\U409_TRANSFER_ACK.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_1_LC_13_8_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_1_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_1_LC_13_8_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_1_LC_13_8_7  (
            .in0(N__5534),
            .in1(N__6471),
            .in2(_gnd_net_),
            .in3(N__6501),
            .lcout(\U409_TRANSFER_ACK.m8_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_6_LC_13_9_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_6_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_6_LC_13_9_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_6_LC_13_9_0  (
            .in0(N__5837),
            .in1(N__5798),
            .in2(N__5769),
            .in3(N__5446),
            .lcout(\U409_TICK.COUNTER60Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6877),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_11_LC_13_9_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_11_LC_13_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_11_LC_13_9_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_11_LC_13_9_1  (
            .in0(N__6941),
            .in1(N__6982),
            .in2(N__7033),
            .in3(N__6619),
            .lcout(\U409_TICK.COUNTER50Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6877),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_9_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_9_2  (
            .in0(N__6064),
            .in1(N__6052),
            .in2(N__6040),
            .in3(N__6015),
            .lcout(),
            .ltout(\U409_TICK.TICK603_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_13_9_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_13_9_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_TICK.COUNTER60_RNI335G2_11_LC_13_9_3  (
            .in0(N__6004),
            .in1(N__5992),
            .in2(N__5986),
            .in3(N__5983),
            .lcout(\U409_TICK.TICK603_14 ),
            .ltout(\U409_TICK.TICK603_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_4_LC_13_9_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_4_LC_13_9_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_4_LC_13_9_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_4_LC_13_9_4  (
            .in0(N__5836),
            .in1(N__5770),
            .in2(N__5971),
            .in3(N__5968),
            .lcout(\U409_TICK.COUNTER60Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6877),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_13_9_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_13_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_13_9_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNICDC71_14_LC_13_9_5  (
            .in0(N__5713),
            .in1(N__5950),
            .in2(N__5938),
            .in3(N__5914),
            .lcout(\U409_TICK.TICK603_9 ),
            .ltout(\U409_TICK.TICK603_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_14_LC_13_9_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_14_LC_13_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_14_LC_13_9_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_14_LC_13_9_6  (
            .in0(N__5758),
            .in1(N__5797),
            .in2(N__5923),
            .in3(N__5920),
            .lcout(\U409_TICK.COUNTER60Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6877),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_13_10_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_13_10_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_TICK.COUNTER60_RNI2USG_10_LC_13_10_3  (
            .in0(N__5901),
            .in1(N__5890),
            .in2(N__5878),
            .in3(N__5854),
            .lcout(\U409_TICK.TICK603_10 ),
            .ltout(\U409_TICK.TICK603_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_15_LC_13_10_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_15_LC_13_10_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_15_LC_13_10_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_15_LC_13_10_4  (
            .in0(N__5838),
            .in1(N__5799),
            .in2(N__5863),
            .in3(N__5860),
            .lcout(\U409_TICK.COUNTER60Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6880),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_9_LC_13_10_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_9_LC_13_10_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_9_LC_13_10_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_9_LC_13_10_6  (
            .in0(N__5839),
            .in1(N__5800),
            .in2(N__5768),
            .in3(N__5719),
            .lcout(\U409_TICK.COUNTER60Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6880),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_13_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_13_11_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_13_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_0_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7166),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .ce(),
            .sr(N__6441));
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_13_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_13_11_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_13_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_1_LC_13_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6499),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .ce(),
            .sr(N__6441));
    defparam \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_13_16_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_13_16_1 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_13_16_1  (
            .in0(N__6360),
            .in1(N__6334),
            .in2(_gnd_net_),
            .in3(N__6810),
            .lcout(TCIn_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_14_4_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_14_4_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_14_4_0 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_14_4_0  (
            .in0(N__6280),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6115),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS1n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNI692L_0_LC_14_4_1 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNI692L_0_LC_14_4_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNI692L_0_LC_14_4_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_CIA.VMA_RNI692L_0_LC_14_4_1  (
            .in0(N__6185),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6774),
            .lcout(CIA_ENABLE),
            .ltout(CIA_ENABLE_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_14_4_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_14_4_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_14_4_2 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_14_4_2  (
            .in0(N__6109),
            .in1(_gnd_net_),
            .in2(N__6091),
            .in3(_gnd_net_),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS0n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_9_LC_14_8_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_9_LC_14_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_9_LC_14_8_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_9_LC_14_8_0  (
            .in0(N__6975),
            .in1(N__6946),
            .in2(N__7030),
            .in3(N__6661),
            .lcout(\U409_TICK.COUNTER50Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6879),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_8_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_8_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_8_1  (
            .in0(N__6835),
            .in1(N__6538),
            .in2(N__6697),
            .in3(N__6557),
            .lcout(),
            .ltout(\U409_TICK.TICK503_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_14_8_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_14_8_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_TICK.COUNTER50_RNITU182_10_LC_14_8_2  (
            .in0(N__6610),
            .in1(N__6589),
            .in2(N__6067),
            .in3(N__6649),
            .lcout(\U409_TICK.TICK503_14 ),
            .ltout(\U409_TICK.TICK503_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_5_LC_14_8_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_5_LC_14_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_5_LC_14_8_3 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \U409_TICK.COUNTER50_5_LC_14_8_3  (
            .in0(N__6736),
            .in1(N__6976),
            .in2(N__6592),
            .in3(N__7018),
            .lcout(\U409_TICK.COUNTER50Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6879),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_14_8_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_14_8_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_TICK.COUNTER50_RNID6CP_3_LC_14_8_4  (
            .in0(N__6748),
            .in1(N__6523),
            .in2(_gnd_net_),
            .in3(N__6578),
            .lcout(\U409_TICK.TICK503_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_14_8_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_14_8_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNIH14V_11_LC_14_8_5  (
            .in0(N__6631),
            .in1(N__6724),
            .in2(N__6679),
            .in3(N__7092),
            .lcout(\U409_TICK.TICK503_9 ),
            .ltout(\U409_TICK.TICK503_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_0_LC_14_8_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_0_LC_14_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_0_LC_14_8_6 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \U409_TICK.COUNTER50_0_LC_14_8_6  (
            .in0(N__7014),
            .in1(N__6945),
            .in2(N__6583),
            .in3(N__6579),
            .lcout(\U409_TICK.COUNTER50Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6879),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_6_LC_14_8_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_6_LC_14_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_6_LC_14_8_7 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_6_LC_14_8_7  (
            .in0(N__6944),
            .in1(N__6977),
            .in2(N__6712),
            .in3(N__7019),
            .lcout(\U409_TICK.COUNTER50Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6879),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_9_0 .C_ON=1'b1;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_9_0  (
            .in0(_gnd_net_),
            .in1(N__6577),
            .in2(N__6559),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_9_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_2_LC_14_9_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_2_LC_14_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_2_LC_14_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_2_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(N__6537),
            .in2(_gnd_net_),
            .in3(N__6526),
            .lcout(\U409_TICK.COUNTER50Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .clk(N__6882),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_3_LC_14_9_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_3_LC_14_9_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_3_LC_14_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_3_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(N__6522),
            .in2(_gnd_net_),
            .in3(N__6511),
            .lcout(\U409_TICK.COUNTER50Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .clk(N__6882),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_4_LC_14_9_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_4_LC_14_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_4_LC_14_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_4_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(N__7059),
            .in2(_gnd_net_),
            .in3(N__6508),
            .lcout(\U409_TICK.COUNTER50Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .clk(N__6882),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_14_9_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_14_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_5_LC_14_9_4  (
            .in0(_gnd_net_),
            .in1(N__6747),
            .in2(_gnd_net_),
            .in3(N__6727),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_14_9_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_14_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_6_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(N__6723),
            .in2(_gnd_net_),
            .in3(N__6703),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_7_LC_14_9_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_7_LC_14_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_7_LC_14_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_7_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(N__7044),
            .in2(_gnd_net_),
            .in3(N__6700),
            .lcout(\U409_TICK.COUNTER50Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .clk(N__6882),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_8_LC_14_9_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_8_LC_14_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_8_LC_14_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_8_LC_14_9_7  (
            .in0(_gnd_net_),
            .in1(N__6693),
            .in2(_gnd_net_),
            .in3(N__6682),
            .lcout(\U409_TICK.COUNTER50Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .clk(N__6882),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_14_10_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_14_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_9_LC_14_10_0  (
            .in0(_gnd_net_),
            .in1(N__6678),
            .in2(_gnd_net_),
            .in3(N__6652),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_14_10_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_10_LC_14_10_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_10_LC_14_10_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_10_LC_14_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_10_LC_14_10_1  (
            .in0(_gnd_net_),
            .in1(N__6645),
            .in2(_gnd_net_),
            .in3(N__6634),
            .lcout(\U409_TICK.COUNTER50Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .clk(N__6885),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_14_10_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_14_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_11_LC_14_10_2  (
            .in0(_gnd_net_),
            .in1(N__6630),
            .in2(_gnd_net_),
            .in3(N__6613),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_12_LC_14_10_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_12_LC_14_10_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_12_LC_14_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_12_LC_14_10_3  (
            .in0(_gnd_net_),
            .in1(N__6606),
            .in2(_gnd_net_),
            .in3(N__6595),
            .lcout(\U409_TICK.COUNTER50Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .clk(N__6885),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_14_10_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_14_10_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_13_LC_14_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7096),
            .in3(N__6847),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_14_10_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_14_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_14_LC_14_10_5  (
            .in0(_gnd_net_),
            .in1(N__7071),
            .in2(_gnd_net_),
            .in3(N__6844),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_14_10_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_14_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_15_LC_14_10_6  (
            .in0(_gnd_net_),
            .in1(N__6897),
            .in2(_gnd_net_),
            .in3(N__6841),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_16_LC_14_10_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_16_LC_14_10_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_16_LC_14_10_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER50_16_LC_14_10_7  (
            .in0(_gnd_net_),
            .in1(N__6834),
            .in2(_gnd_net_),
            .in3(N__6838),
            .lcout(\U409_TICK.COUNTER50Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6885),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_14_11_0 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_14_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_0_LC_14_11_0  (
            .in0(N__7455),
            .in1(N__7414),
            .in2(N__7330),
            .in3(N__7431),
            .lcout(),
            .ltout(\U409_CIA.CLK_CIA6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_LC_14_11_1 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_LC_14_11_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CLK_CIA_LC_14_11_1 .LUT_INIT=16'b1001101010101010;
    LogicCell40 \U409_CIA.CLK_CIA_LC_14_11_1  (
            .in0(N__7165),
            .in1(N__7213),
            .in2(N__6820),
            .in3(N__7144),
            .lcout(CLK_CIA_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7383),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_1_LC_14_11_2 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_1_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_1_LC_14_11_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_CIA.VMA_RNO_1_LC_14_11_2  (
            .in0(N__7271),
            .in1(N__7295),
            .in2(N__7218),
            .in3(N__7413),
            .lcout(),
            .ltout(\U409_CIA.un1_CIA_CLK_COUNT_3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_0_LC_14_11_3 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_0_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_0_LC_14_11_3 .LUT_INIT=16'b0100000010000000;
    LogicCell40 \U409_CIA.VMA_RNO_0_LC_14_11_3  (
            .in0(N__7325),
            .in1(N__7346),
            .in2(N__6817),
            .in3(N__7242),
            .lcout(),
            .ltout(\U409_CIA.VMA_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_LC_14_11_4 .C_ON=1'b0;
    defparam \U409_CIA.VMA_LC_14_11_4 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.VMA_LC_14_11_4 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \U409_CIA.VMA_LC_14_11_4  (
            .in0(N__6814),
            .in1(N__6764),
            .in2(N__6778),
            .in3(N__7326),
            .lcout(\U409_CIA.VMAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7383),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_14_11_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_14_11_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_14_11_6  (
            .in0(_gnd_net_),
            .in1(N__7430),
            .in2(_gnd_net_),
            .in3(N__7454),
            .lcout(\U409_CIA.CLK_CIA6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_14_11_7 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_14_11_7 .LUT_INIT=16'b0000010000010000;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_1_LC_14_11_7  (
            .in0(N__7296),
            .in1(N__7243),
            .in2(N__7170),
            .in3(N__7272),
            .lcout(\U409_CIA.CLK_CIA_r_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK50_LC_15_8_1 .C_ON=1'b0;
    defparam \U409_TICK.TICK50_LC_15_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK50_LC_15_8_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \U409_TICK.TICK50_LC_15_8_1  (
            .in0(N__6939),
            .in1(N__6979),
            .in2(N__7031),
            .in3(N__7122),
            .lcout(TICK50_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6883),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_13_LC_15_8_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_13_LC_15_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_13_LC_15_8_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_13_LC_15_8_2  (
            .in0(N__6978),
            .in1(N__6940),
            .in2(N__7111),
            .in3(N__7023),
            .lcout(\U409_TICK.COUNTER50Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6883),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_14_LC_15_9_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_14_LC_15_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_14_LC_15_9_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_14_LC_15_9_3  (
            .in0(N__6980),
            .in1(N__6942),
            .in2(N__7032),
            .in3(N__7078),
            .lcout(\U409_TICK.COUNTER50Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6886),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_15_9_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_15_9_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNII24V_14_LC_15_9_6  (
            .in0(N__7072),
            .in1(N__7060),
            .in2(N__7048),
            .in3(N__6898),
            .lcout(\U409_TICK.TICK503_10 ),
            .ltout(\U409_TICK.TICK503_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_15_LC_15_9_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_15_LC_15_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_15_LC_15_9_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_15_LC_15_9_7  (
            .in0(N__6981),
            .in1(N__6943),
            .in2(N__6907),
            .in3(N__6904),
            .lcout(\U409_TICK.COUNTER50Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6886),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_15_10_0 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_15_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_15_10_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_5_LC_15_10_0  (
            .in0(N__7348),
            .in1(N__7369),
            .in2(N__7363),
            .in3(N__7192),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7384),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_15_10_2 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_15_10_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_15_10_2  (
            .in0(N__7273),
            .in1(N__7297),
            .in2(N__7219),
            .in3(N__7415),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_15_10_3 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_15_10_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_15_10_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_1_LC_15_10_3  (
            .in0(N__7324),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7416),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7384),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNI9DRM_4_LC_15_10_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNI9DRM_4_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNI9DRM_4_LC_15_10_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNI9DRM_4_LC_15_10_4  (
            .in0(N__7241),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7323),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_2 ),
            .ltout(\U409_CIA.CIA_CLK_COUNT11_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_15_10_5 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_15_10_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_15_10_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_3_LC_15_10_5  (
            .in0(N__7359),
            .in1(N__7347),
            .in2(N__7333),
            .in3(N__7252),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7384),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_15_11_0 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_15_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(N__7322),
            .in2(N__7417),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_11_0_),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_15_11_1 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_15_11_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_15_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_2_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__7294),
            .in2(_gnd_net_),
            .in3(N__7276),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .clk(N__7382),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_3_LC_15_11_2 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_3_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_3_LC_15_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNO_0_3_LC_15_11_2  (
            .in0(_gnd_net_),
            .in1(N__7270),
            .in2(_gnd_net_),
            .in3(N__7246),
            .lcout(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_15_11_3 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_15_11_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_15_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_4_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(N__7240),
            .in2(_gnd_net_),
            .in3(N__7222),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .clk(N__7382),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_15_11_4 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_15_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_15_11_4  (
            .in0(_gnd_net_),
            .in1(N__7214),
            .in2(_gnd_net_),
            .in3(N__7186),
            .lcout(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_15_11_5 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_15_11_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_15_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_6_LC_15_11_5  (
            .in0(_gnd_net_),
            .in1(N__7456),
            .in2(_gnd_net_),
            .in3(N__7438),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ),
            .clk(N__7382),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_15_11_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_15_11_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_15_11_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_7_LC_15_11_6  (
            .in0(_gnd_net_),
            .in1(N__7432),
            .in2(_gnd_net_),
            .in3(N__7435),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7382),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_15_11_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_15_11_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_15_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_0_LC_15_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7412),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7382),
            .ce(),
            .sr(_gnd_net_));
endmodule // U409_TOP

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     May 16 2025 17:23:40

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    DA : out std_logic_vector(2 downto 0);
    A : in std_logic_vector(20 downto 0);
    DBRn : in std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    TCIn : out std_logic;
    TBIn : out std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__12697\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12382\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12211\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12146\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7827\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_6_6_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_CHIP_RAM.N_489_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_1\ : std_logic;
signal \U712_CHIP_RAM.N_413_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_159_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_413\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_cascade_\ : std_logic;
signal \LATCH_CLK_c\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.N_462\ : std_logic;
signal \U712_CHIP_RAM.N_443\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_1_2\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_1_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_3\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_7\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_383\ : std_logic;
signal \U712_REG_SM.N_339\ : std_logic;
signal \U712_REG_SM.N_339_cascade_\ : std_logic;
signal \U712_REG_SM.N_350\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_REG_SM.N_573\ : std_logic;
signal \U712_REG_SM.N_573_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_4\ : std_logic;
signal \U712_REG_SM.N_426\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_463_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_485_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_325\ : std_logic;
signal \U712_CHIP_RAM.N_329_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_389\ : std_logic;
signal \U712_CHIP_RAM.N_489\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_a2_1\ : std_logic;
signal \U712_CHIP_RAM.N_441_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a7_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.N_475_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0\ : std_logic;
signal \U712_CHIP_RAM.DBENn_8_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CYCLE_TERM.N_466_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\ : std_logic;
signal \DBR_SYNC_i_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3\ : std_logic;
signal \U712_REG_SM.N_337_cascade_\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_5_iv_0_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_424\ : std_logic;
signal \U712_REG_SM.N_338_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_5\ : std_logic;
signal \U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_6\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_7\ : std_logic;
signal \U712_REG_SM.REGENn_e_1\ : std_logic;
signal \REGENn_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_463\ : std_logic;
signal \U712_CHIP_RAM.N_461\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.N_47\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.N_574_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_475\ : std_logic;
signal \U712_CHIP_RAM.N_328\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto7_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lt7\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3\ : std_logic;
signal \U712_CHIP_RAM.N_327\ : std_logic;
signal \TSn_c\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_CYCLE_TERM.N_340\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_416\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.START_RSTZ0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_8\ : std_logic;
signal \U712_REG_SM.STATE_COUNTsr_0\ : std_logic;
signal \U712_REG_SM.N_338\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \UDSn_c\ : std_logic;
signal \U712_REG_SM.N_435\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \U712_CHIP_RAM.N_320\ : std_logic;
signal \U712_CHIP_RAM.N_480\ : std_logic;
signal \U712_CHIP_RAM.N_571_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.N_326\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_i_a2_0_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_572\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER19\ : std_logic;
signal \U712_CHIP_RAM.N_574\ : std_logic;
signal \U712_CHIP_RAM.N_571\ : std_logic;
signal \U712_CHIP_RAM.N_566\ : std_logic;
signal \U712_CHIP_RAM.N_477\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_555\ : std_logic;
signal \U712_CHIP_RAM.N_349\ : std_logic;
signal \U712_CHIP_RAM.N_447\ : std_logic;
signal \U712_CHIP_RAM.N_444_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0\ : std_logic;
signal \U712_CHIP_RAM.N_410\ : std_logic;
signal \U712_CHIP_RAM.N_411\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_476\ : std_logic;
signal \U712_CHIP_RAM.N_446\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_i_i_a2_1_0\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_431\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_471\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_5\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ1Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ1Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3_cascade_\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_433\ : std_logic;
signal \LDSn_c\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_i_i_0\ : std_logic;
signal \U712_CHIP_RAM.N_408\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.N_151\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_4\ : std_logic;
signal \N_217_i\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \N_182_i\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_434\ : std_logic;
signal \N_198_i\ : std_logic;
signal \N_343_i\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_374\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA25_0_i_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.N_368\ : std_logic;
signal \U712_CHIP_RAM.N_330_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\ : std_logic;
signal \U712_BYTE_ENABLE.N_454_cascade_\ : std_logic;
signal \N_215_i\ : std_logic;
signal \N_213_i\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \U712_BYTE_ENABLE.N_450_cascade_\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \N_211_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_456\ : std_logic;
signal \U712_BYTE_ENABLE.N_315_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_452\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_3\ : std_logic;
signal \N_322\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \N_342_i\ : std_logic;
signal \N_345_i\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \A_c_1\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \N_344_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_i_0_9\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.N_330\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA25_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_171\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \WEn_c\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.N_171_0\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_1\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_0\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \RnW_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \DMA_WRITE_CYCLE\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \N_385\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \DA_wire\ : std_logic_vector(2 downto 0);
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    TBIn <= \TBIn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    ASn <= \ASn_wire\;
    DA <= \DA_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    TCIn <= \TCIn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__4380\,
            RESETB => \N__6342\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12697\,
            DIN => \N__12696\,
            DOUT => \N__12695\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12697\,
            PADOUT => \N__12696\,
            PADIN => \N__12695\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8484\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12688\,
            DIN => \N__12687\,
            DOUT => \N__12686\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12688\,
            PADOUT => \N__12687\,
            PADIN => \N__12686\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12679\,
            DIN => \N__12678\,
            DOUT => \N__12677\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12679\,
            PADOUT => \N__12678\,
            PADIN => \N__12677\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8235\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12670\,
            DIN => \N__12669\,
            DOUT => \N__12668\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12670\,
            PADOUT => \N__12669\,
            PADIN => \N__12668\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11724\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12661\,
            DIN => \N__12660\,
            DOUT => \N__12659\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12661\,
            PADOUT => \N__12660\,
            PADIN => \N__12659\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12652\,
            DIN => \N__12651\,
            DOUT => \N__12650\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12652\,
            PADOUT => \N__12651\,
            PADIN => \N__12650\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12643\,
            DIN => \N__12642\,
            DOUT => \N__12641\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12643\,
            PADOUT => \N__12642\,
            PADIN => \N__12641\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12634\,
            DIN => \N__12633\,
            DOUT => \N__12632\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12634\,
            PADOUT => \N__12633\,
            PADIN => \N__12632\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12625\,
            DIN => \N__12624\,
            DOUT => \N__12623\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12625\,
            PADOUT => \N__12624\,
            PADIN => \N__12623\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12616\,
            DIN => \N__12615\,
            DOUT => \N__12614\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12616\,
            PADOUT => \N__12615\,
            PADIN => \N__12614\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12607\,
            DIN => \N__12606\,
            DOUT => \N__12605\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12607\,
            PADOUT => \N__12606\,
            PADIN => \N__12605\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12598\,
            DIN => \N__12597\,
            DOUT => \N__12596\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12598\,
            PADOUT => \N__12597\,
            PADIN => \N__12596\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9411\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12589\,
            DIN => \N__12588\,
            DOUT => \N__12587\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12589\,
            PADOUT => \N__12588\,
            PADIN => \N__12587\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9168\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12580\,
            DIN => \N__12579\,
            DOUT => \N__12578\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12580\,
            PADOUT => \N__12579\,
            PADIN => \N__12578\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12571\,
            DIN => \N__12570\,
            DOUT => \N__12569\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12571\,
            PADOUT => \N__12570\,
            PADIN => \N__12569\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12562\,
            DIN => \N__12561\,
            DOUT => \N__12560\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12562\,
            PADOUT => \N__12561\,
            PADIN => \N__12560\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12553\,
            DIN => \N__12552\,
            DOUT => \N__12551\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12553\,
            PADOUT => \N__12552\,
            PADIN => \N__12551\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5262\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12544\,
            DIN => \N__12543\,
            DOUT => \N__12542\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12544\,
            PADOUT => \N__12543\,
            PADIN => \N__12542\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12535\,
            DIN => \N__12534\,
            DOUT => \N__12533\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12535\,
            PADOUT => \N__12534\,
            PADIN => \N__12533\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12526\,
            DIN => \N__12525\,
            DOUT => \N__12524\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12526\,
            PADOUT => \N__12525\,
            PADIN => \N__12524\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8712\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12517\,
            DIN => \N__12516\,
            DOUT => \N__12515\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12517\,
            PADOUT => \N__12516\,
            PADIN => \N__12515\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12508\,
            DIN => \N__12507\,
            DOUT => \N__12506\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12508\,
            PADOUT => \N__12507\,
            PADIN => \N__12506\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8736\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12499\,
            DIN => \N__12498\,
            DOUT => \N__12497\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12499\,
            PADOUT => \N__12498\,
            PADIN => \N__12497\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12490\,
            DIN => \N__12489\,
            DOUT => \N__12488\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12490\,
            PADOUT => \N__12489\,
            PADIN => \N__12488\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9180\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12481\,
            DIN => \N__12480\,
            DOUT => \N__12479\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12481\,
            PADOUT => \N__12480\,
            PADIN => \N__12479\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5612\,
            DIN0 => OPEN,
            DOUT0 => \N__5679\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12472\,
            DIN => \N__12471\,
            DOUT => \N__12470\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12472\,
            PADOUT => \N__12471\,
            PADIN => \N__12470\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12463\,
            DIN => \N__12462\,
            DOUT => \N__12461\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12463\,
            PADOUT => \N__12462\,
            PADIN => \N__12461\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12454\,
            DIN => \N__12453\,
            DOUT => \N__12452\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12454\,
            PADOUT => \N__12453\,
            PADIN => \N__12452\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12445\,
            DIN => \N__12444\,
            DOUT => \N__12443\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12445\,
            PADOUT => \N__12444\,
            PADIN => \N__12443\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12436\,
            DIN => \N__12435\,
            DOUT => \N__12434\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12436\,
            PADOUT => \N__12435\,
            PADIN => \N__12434\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12427\,
            DIN => \N__12426\,
            DOUT => \N__12425\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12427\,
            PADOUT => \N__12426\,
            PADIN => \N__12425\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8001\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12418\,
            DIN => \N__12417\,
            DOUT => \N__12416\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12418\,
            PADOUT => \N__12417\,
            PADIN => \N__12416\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12409\,
            DIN => \N__12408\,
            DOUT => \N__12407\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12409\,
            PADOUT => \N__12408\,
            PADIN => \N__12407\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12400\,
            DIN => \N__12399\,
            DOUT => \N__12398\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12400\,
            PADOUT => \N__12399\,
            PADIN => \N__12398\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12391\,
            DIN => \N__12390\,
            DOUT => \N__12389\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12391\,
            PADOUT => \N__12390\,
            PADIN => \N__12389\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12382\,
            DIN => \N__12381\,
            DOUT => \N__12380\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12382\,
            PADOUT => \N__12381\,
            PADIN => \N__12380\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12373\,
            DIN => \N__12372\,
            DOUT => \N__12371\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12373\,
            PADOUT => \N__12372\,
            PADIN => \N__12371\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9801\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12364\,
            DIN => \N__12363\,
            DOUT => \N__12362\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12364\,
            PADOUT => \N__12363\,
            PADIN => \N__12362\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12355\,
            DIN => \N__12354\,
            DOUT => \N__12353\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12355\,
            PADOUT => \N__12354\,
            PADIN => \N__12353\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12346\,
            DIN => \N__12345\,
            DOUT => \N__12344\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12346\,
            PADOUT => \N__12345\,
            PADIN => \N__12344\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11202\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12337\,
            DIN => \N__12336\,
            DOUT => \N__12335\,
            PACKAGEPIN => \DA_wire\(0)
        );

    \DA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12337\,
            PADOUT => \N__12336\,
            PADIN => \N__12335\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7455\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12328\,
            DIN => \N__12327\,
            DOUT => \N__12326\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12328\,
            PADOUT => \N__12327\,
            PADIN => \N__12326\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12319\,
            DIN => \N__12318\,
            DOUT => \N__12317\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12319\,
            PADOUT => \N__12318\,
            PADIN => \N__12317\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8178\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12310\,
            DIN => \N__12309\,
            DOUT => \N__12308\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12310\,
            PADOUT => \N__12309\,
            PADIN => \N__12308\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9474\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12301\,
            DIN => \N__12300\,
            DOUT => \N__12299\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12301\,
            PADOUT => \N__12300\,
            PADIN => \N__12299\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5364\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12292\,
            DIN => \N__12291\,
            DOUT => \N__12290\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12292\,
            PADOUT => \N__12291\,
            PADIN => \N__12290\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12283\,
            DIN => \N__12282\,
            DOUT => \N__12281\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12283\,
            PADOUT => \N__12282\,
            PADIN => \N__12281\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12274\,
            DIN => \N__12273\,
            DOUT => \N__12272\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12274\,
            PADOUT => \N__12273\,
            PADIN => \N__12272\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8520\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12265\,
            DIN => \N__12264\,
            DOUT => \N__12263\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12265\,
            PADOUT => \N__12264\,
            PADIN => \N__12263\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5616\,
            DIN0 => OPEN,
            DOUT0 => \N__5678\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12256\,
            DIN => \N__12255\,
            DOUT => \N__12254\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12256\,
            PADOUT => \N__12255\,
            PADIN => \N__12254\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11646\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12247\,
            DIN => \N__12246\,
            DOUT => \N__12245\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12247\,
            PADOUT => \N__12246\,
            PADIN => \N__12245\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5703\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12238\,
            DIN => \N__12237\,
            DOUT => \N__12236\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12238\,
            PADOUT => \N__12237\,
            PADIN => \N__12236\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8505\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12229\,
            DIN => \N__12228\,
            DOUT => \N__12227\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12229\,
            PADOUT => \N__12228\,
            PADIN => \N__12227\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12220\,
            DIN => \N__12219\,
            DOUT => \N__12218\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12220\,
            PADOUT => \N__12219\,
            PADIN => \N__12218\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12211\,
            DIN => \N__12210\,
            DOUT => \N__12209\,
            PACKAGEPIN => \DA_wire\(2)
        );

    \DA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12211\,
            PADOUT => \N__12210\,
            PADIN => \N__12209\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6891\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12202\,
            DIN => \N__12201\,
            DOUT => \N__12200\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12202\,
            PADOUT => \N__12201\,
            PADIN => \N__12200\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12193\,
            DIN => \N__12192\,
            DOUT => \N__12191\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12193\,
            PADOUT => \N__12192\,
            PADIN => \N__12191\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12184\,
            DIN => \N__12183\,
            DOUT => \N__12182\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12184\,
            PADOUT => \N__12183\,
            PADIN => \N__12182\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8160\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12175\,
            DIN => \N__12174\,
            DOUT => \N__12173\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12175\,
            PADOUT => \N__12174\,
            PADIN => \N__12173\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8796\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12166\,
            DIN => \N__12165\,
            DOUT => \N__12164\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12166\,
            PADOUT => \N__12165\,
            PADIN => \N__12164\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12157\,
            DIN => \N__12156\,
            DOUT => \N__12155\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12157\,
            PADOUT => \N__12156\,
            PADIN => \N__12155\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8376\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12148\,
            DIN => \N__12147\,
            DOUT => \N__12146\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12148\,
            PADOUT => \N__12147\,
            PADIN => \N__12146\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5602\,
            DIN0 => OPEN,
            DOUT0 => \N__5671\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12139\,
            DIN => \N__12138\,
            DOUT => \N__12137\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12139\,
            PADOUT => \N__12138\,
            PADIN => \N__12137\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7956\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12130\,
            DIN => \N__12129\,
            DOUT => \N__12128\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12130\,
            PADOUT => \N__12129\,
            PADIN => \N__12128\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12121\,
            DIN => \N__12120\,
            DOUT => \N__12119\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12121\,
            PADOUT => \N__12120\,
            PADIN => \N__12119\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12112\,
            DIN => \N__12111\,
            DOUT => \N__12110\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12112\,
            PADOUT => \N__12111\,
            PADIN => \N__12110\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9285\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12103\,
            DIN => \N__12102\,
            DOUT => \N__12101\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12103\,
            PADOUT => \N__12102\,
            PADIN => \N__12101\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12094\,
            DIN => \N__12093\,
            DOUT => \N__12092\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12094\,
            PADOUT => \N__12093\,
            PADIN => \N__12092\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12085\,
            DIN => \N__12084\,
            DOUT => \N__12083\,
            PACKAGEPIN => \DA_wire\(1)
        );

    \DA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12085\,
            PADOUT => \N__12084\,
            PADIN => \N__12083\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7878\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12076\,
            DIN => \N__12075\,
            DOUT => \N__12074\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12076\,
            PADOUT => \N__12075\,
            PADIN => \N__12074\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12067\,
            DIN => \N__12066\,
            DOUT => \N__12065\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12067\,
            PADOUT => \N__12066\,
            PADIN => \N__12065\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12058\,
            DIN => \N__12057\,
            DOUT => \N__12056\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12058\,
            PADOUT => \N__12057\,
            PADIN => \N__12056\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8202\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12049\,
            DIN => \N__12048\,
            DOUT => \N__12047\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12049\,
            PADOUT => \N__12048\,
            PADIN => \N__12047\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6378\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12040\,
            DIN => \N__12039\,
            DOUT => \N__12038\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12040\,
            PADOUT => \N__12039\,
            PADIN => \N__12038\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7989\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12031\,
            DIN => \N__12030\,
            DOUT => \N__12029\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12031\,
            PADOUT => \N__12030\,
            PADIN => \N__12029\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4461\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12022\,
            DIN => \N__12021\,
            DOUT => \N__12020\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12022\,
            PADOUT => \N__12021\,
            PADIN => \N__12020\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12013\,
            DIN => \N__12012\,
            DOUT => \N__12011\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12013\,
            PADOUT => \N__12012\,
            PADIN => \N__12011\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12004\,
            DIN => \N__12003\,
            DOUT => \N__12002\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12004\,
            PADOUT => \N__12003\,
            PADIN => \N__12002\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9444\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11995\,
            DIN => \N__11994\,
            DOUT => \N__11993\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11995\,
            PADOUT => \N__11994\,
            PADIN => \N__11993\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11986\,
            DIN => \N__11985\,
            DOUT => \N__11984\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11986\,
            PADOUT => \N__11985\,
            PADIN => \N__11984\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11977\,
            DIN => \N__11976\,
            DOUT => \N__11975\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11977\,
            PADOUT => \N__11976\,
            PADIN => \N__11975\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4734\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11968\,
            DIN => \N__11967\,
            DOUT => \N__11966\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11968\,
            PADOUT => \N__11967\,
            PADIN => \N__11966\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7485\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11959\,
            DIN => \N__11958\,
            DOUT => \N__11957\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11959\,
            PADOUT => \N__11958\,
            PADIN => \N__11957\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6141\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11950\,
            DIN => \N__11949\,
            DOUT => \N__11948\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11950\,
            PADOUT => \N__11949\,
            PADIN => \N__11948\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11941\,
            DIN => \N__11940\,
            DOUT => \N__11939\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11941\,
            PADOUT => \N__11940\,
            PADIN => \N__11939\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6137\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11932\,
            DIN => \N__11931\,
            DOUT => \N__11930\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11932\,
            PADOUT => \N__11931\,
            PADIN => \N__11930\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4407\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11923\,
            DIN => \N__11922\,
            DOUT => \N__11921\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11923\,
            PADOUT => \N__11922\,
            PADIN => \N__11921\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9501\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11914\,
            DIN => \N__11913\,
            DOUT => \N__11912\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11914\,
            PADOUT => \N__11913\,
            PADIN => \N__11912\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11905\,
            DIN => \N__11904\,
            DOUT => \N__11903\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11905\,
            PADOUT => \N__11904\,
            PADIN => \N__11903\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11896\,
            DIN => \N__11895\,
            DOUT => \N__11894\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11896\,
            PADOUT => \N__11895\,
            PADIN => \N__11894\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11887\,
            DIN => \N__11886\,
            DOUT => \N__11885\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11887\,
            PADOUT => \N__11886\,
            PADIN => \N__11885\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11878\,
            DIN => \N__11877\,
            DOUT => \N__11876\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11878\,
            PADOUT => \N__11877\,
            PADIN => \N__11876\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6125\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11869\,
            DIN => \N__11868\,
            DOUT => \N__11867\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11869\,
            PADOUT => \N__11868\,
            PADIN => \N__11867\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8037\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11860\,
            DIN => \N__11859\,
            DOUT => \N__11858\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11860\,
            PADOUT => \N__11859\,
            PADIN => \N__11858\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8088\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11851\,
            DIN => \N__11850\,
            DOUT => \N__11849\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11851\,
            PADOUT => \N__11850\,
            PADIN => \N__11849\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9528\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2866\ : CascadeMux
    port map (
            O => \N__11832\,
            I => \N__11828\
        );

    \I__2865\ : InMux
    port map (
            O => \N__11831\,
            I => \N__11825\
        );

    \I__2864\ : InMux
    port map (
            O => \N__11828\,
            I => \N__11822\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__11825\,
            I => \N__11819\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__11822\,
            I => \N__11816\
        );

    \I__2861\ : Span4Mux_h
    port map (
            O => \N__11819\,
            I => \N__11813\
        );

    \I__2860\ : Span12Mux_h
    port map (
            O => \N__11816\,
            I => \N__11810\
        );

    \I__2859\ : Span4Mux_v
    port map (
            O => \N__11813\,
            I => \N__11807\
        );

    \I__2858\ : Span12Mux_v
    port map (
            O => \N__11810\,
            I => \N__11803\
        );

    \I__2857\ : Sp12to4
    port map (
            O => \N__11807\,
            I => \N__11800\
        );

    \I__2856\ : InMux
    port map (
            O => \N__11806\,
            I => \N__11797\
        );

    \I__2855\ : Odrv12
    port map (
            O => \N__11803\,
            I => \DMA_WRITE_CYCLE\
        );

    \I__2854\ : Odrv12
    port map (
            O => \N__11800\,
            I => \DMA_WRITE_CYCLE\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__11797\,
            I => \DMA_WRITE_CYCLE\
        );

    \I__2852\ : CascadeMux
    port map (
            O => \N__11790\,
            I => \N__11785\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__11789\,
            I => \N__11782\
        );

    \I__2850\ : InMux
    port map (
            O => \N__11788\,
            I => \N__11779\
        );

    \I__2849\ : InMux
    port map (
            O => \N__11785\,
            I => \N__11776\
        );

    \I__2848\ : InMux
    port map (
            O => \N__11782\,
            I => \N__11773\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__11779\,
            I => \N__11766\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__11776\,
            I => \N__11766\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__11773\,
            I => \N__11763\
        );

    \I__2844\ : InMux
    port map (
            O => \N__11772\,
            I => \N__11760\
        );

    \I__2843\ : InMux
    port map (
            O => \N__11771\,
            I => \N__11757\
        );

    \I__2842\ : Span4Mux_v
    port map (
            O => \N__11766\,
            I => \N__11750\
        );

    \I__2841\ : Span4Mux_h
    port map (
            O => \N__11763\,
            I => \N__11750\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__11760\,
            I => \N__11750\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__11757\,
            I => \N__11747\
        );

    \I__2838\ : Sp12to4
    port map (
            O => \N__11750\,
            I => \N__11741\
        );

    \I__2837\ : Sp12to4
    port map (
            O => \N__11747\,
            I => \N__11741\
        );

    \I__2836\ : InMux
    port map (
            O => \N__11746\,
            I => \N__11738\
        );

    \I__2835\ : Span12Mux_v
    port map (
            O => \N__11741\,
            I => \N__11735\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__11738\,
            I => \N__11732\
        );

    \I__2833\ : Span12Mux_h
    port map (
            O => \N__11735\,
            I => \N__11727\
        );

    \I__2832\ : Span12Mux_v
    port map (
            O => \N__11732\,
            I => \N__11727\
        );

    \I__2831\ : Odrv12
    port map (
            O => \N__11727\,
            I => \CASLn_c\
        );

    \I__2830\ : IoInMux
    port map (
            O => \N__11724\,
            I => \N__11721\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__11721\,
            I => \N__11718\
        );

    \I__2828\ : IoSpan4Mux
    port map (
            O => \N__11718\,
            I => \N__11715\
        );

    \I__2827\ : Span4Mux_s3_v
    port map (
            O => \N__11715\,
            I => \N__11712\
        );

    \I__2826\ : Span4Mux_v
    port map (
            O => \N__11712\,
            I => \N__11709\
        );

    \I__2825\ : Odrv4
    port map (
            O => \N__11709\,
            I => \N_385\
        );

    \I__2824\ : InMux
    port map (
            O => \N__11706\,
            I => \N__11700\
        );

    \I__2823\ : InMux
    port map (
            O => \N__11705\,
            I => \N__11700\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__11700\,
            I => \N__11697\
        );

    \I__2821\ : Odrv12
    port map (
            O => \N__11697\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2820\ : InMux
    port map (
            O => \N__11694\,
            I => \N__11689\
        );

    \I__2819\ : InMux
    port map (
            O => \N__11693\,
            I => \N__11686\
        );

    \I__2818\ : InMux
    port map (
            O => \N__11692\,
            I => \N__11683\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__11689\,
            I => \N__11676\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__11686\,
            I => \N__11676\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__11683\,
            I => \N__11676\
        );

    \I__2814\ : Odrv12
    port map (
            O => \N__11676\,
            I => \U712_REG_SM.N_171\
        );

    \I__2813\ : InMux
    port map (
            O => \N__11673\,
            I => \N__11670\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__11670\,
            I => \N__11663\
        );

    \I__2811\ : InMux
    port map (
            O => \N__11669\,
            I => \N__11658\
        );

    \I__2810\ : InMux
    port map (
            O => \N__11668\,
            I => \N__11658\
        );

    \I__2809\ : InMux
    port map (
            O => \N__11667\,
            I => \N__11653\
        );

    \I__2808\ : InMux
    port map (
            O => \N__11666\,
            I => \N__11653\
        );

    \I__2807\ : Odrv12
    port map (
            O => \N__11663\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__11658\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__11653\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2804\ : IoInMux
    port map (
            O => \N__11646\,
            I => \N__11643\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__11643\,
            I => \N__11640\
        );

    \I__2802\ : Span4Mux_s1_h
    port map (
            O => \N__11640\,
            I => \N__11637\
        );

    \I__2801\ : Span4Mux_h
    port map (
            O => \N__11637\,
            I => \N__11634\
        );

    \I__2800\ : Sp12to4
    port map (
            O => \N__11634\,
            I => \N__11631\
        );

    \I__2799\ : Span12Mux_s11_v
    port map (
            O => \N__11631\,
            I => \N__11628\
        );

    \I__2798\ : Odrv12
    port map (
            O => \N__11628\,
            I => \WEn_c\
        );

    \I__2797\ : InMux
    port map (
            O => \N__11625\,
            I => \N__11621\
        );

    \I__2796\ : InMux
    port map (
            O => \N__11624\,
            I => \N__11618\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__11621\,
            I => \N__11612\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__11618\,
            I => \N__11612\
        );

    \I__2793\ : InMux
    port map (
            O => \N__11617\,
            I => \N__11609\
        );

    \I__2792\ : Span4Mux_h
    port map (
            O => \N__11612\,
            I => \N__11604\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__11609\,
            I => \N__11604\
        );

    \I__2790\ : Span4Mux_v
    port map (
            O => \N__11604\,
            I => \N__11600\
        );

    \I__2789\ : InMux
    port map (
            O => \N__11603\,
            I => \N__11597\
        );

    \I__2788\ : Sp12to4
    port map (
            O => \N__11600\,
            I => \N__11594\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__11597\,
            I => \N__11591\
        );

    \I__2786\ : Span12Mux_h
    port map (
            O => \N__11594\,
            I => \N__11588\
        );

    \I__2785\ : Span12Mux_v
    port map (
            O => \N__11591\,
            I => \N__11585\
        );

    \I__2784\ : Span12Mux_v
    port map (
            O => \N__11588\,
            I => \N__11582\
        );

    \I__2783\ : Span12Mux_v
    port map (
            O => \N__11585\,
            I => \N__11579\
        );

    \I__2782\ : Odrv12
    port map (
            O => \N__11582\,
            I => \DRA_c_9\
        );

    \I__2781\ : Odrv12
    port map (
            O => \N__11579\,
            I => \DRA_c_9\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__11574\,
            I => \N__11571\
        );

    \I__2779\ : InMux
    port map (
            O => \N__11571\,
            I => \N__11568\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__11568\,
            I => \N__11561\
        );

    \I__2777\ : InMux
    port map (
            O => \N__11567\,
            I => \N__11558\
        );

    \I__2776\ : CascadeMux
    port map (
            O => \N__11566\,
            I => \N__11553\
        );

    \I__2775\ : CascadeMux
    port map (
            O => \N__11565\,
            I => \N__11548\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__11564\,
            I => \N__11538\
        );

    \I__2773\ : Span4Mux_h
    port map (
            O => \N__11561\,
            I => \N__11534\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__11558\,
            I => \N__11531\
        );

    \I__2771\ : InMux
    port map (
            O => \N__11557\,
            I => \N__11528\
        );

    \I__2770\ : InMux
    port map (
            O => \N__11556\,
            I => \N__11524\
        );

    \I__2769\ : InMux
    port map (
            O => \N__11553\,
            I => \N__11517\
        );

    \I__2768\ : InMux
    port map (
            O => \N__11552\,
            I => \N__11517\
        );

    \I__2767\ : InMux
    port map (
            O => \N__11551\,
            I => \N__11517\
        );

    \I__2766\ : InMux
    port map (
            O => \N__11548\,
            I => \N__11510\
        );

    \I__2765\ : InMux
    port map (
            O => \N__11547\,
            I => \N__11510\
        );

    \I__2764\ : InMux
    port map (
            O => \N__11546\,
            I => \N__11510\
        );

    \I__2763\ : InMux
    port map (
            O => \N__11545\,
            I => \N__11505\
        );

    \I__2762\ : InMux
    port map (
            O => \N__11544\,
            I => \N__11505\
        );

    \I__2761\ : InMux
    port map (
            O => \N__11543\,
            I => \N__11499\
        );

    \I__2760\ : InMux
    port map (
            O => \N__11542\,
            I => \N__11499\
        );

    \I__2759\ : InMux
    port map (
            O => \N__11541\,
            I => \N__11496\
        );

    \I__2758\ : InMux
    port map (
            O => \N__11538\,
            I => \N__11491\
        );

    \I__2757\ : InMux
    port map (
            O => \N__11537\,
            I => \N__11491\
        );

    \I__2756\ : Span4Mux_h
    port map (
            O => \N__11534\,
            I => \N__11484\
        );

    \I__2755\ : Span4Mux_v
    port map (
            O => \N__11531\,
            I => \N__11484\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__11528\,
            I => \N__11484\
        );

    \I__2753\ : InMux
    port map (
            O => \N__11527\,
            I => \N__11481\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__11524\,
            I => \N__11478\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__11517\,
            I => \N__11471\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__11510\,
            I => \N__11471\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__11505\,
            I => \N__11468\
        );

    \I__2748\ : InMux
    port map (
            O => \N__11504\,
            I => \N__11465\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__11499\,
            I => \N__11458\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__11496\,
            I => \N__11458\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__11491\,
            I => \N__11458\
        );

    \I__2744\ : Span4Mux_h
    port map (
            O => \N__11484\,
            I => \N__11453\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__11481\,
            I => \N__11453\
        );

    \I__2742\ : Span4Mux_v
    port map (
            O => \N__11478\,
            I => \N__11450\
        );

    \I__2741\ : InMux
    port map (
            O => \N__11477\,
            I => \N__11447\
        );

    \I__2740\ : InMux
    port map (
            O => \N__11476\,
            I => \N__11444\
        );

    \I__2739\ : Span4Mux_v
    port map (
            O => \N__11471\,
            I => \N__11437\
        );

    \I__2738\ : Span4Mux_h
    port map (
            O => \N__11468\,
            I => \N__11437\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__11465\,
            I => \N__11437\
        );

    \I__2736\ : Span4Mux_v
    port map (
            O => \N__11458\,
            I => \N__11432\
        );

    \I__2735\ : Span4Mux_v
    port map (
            O => \N__11453\,
            I => \N__11432\
        );

    \I__2734\ : Sp12to4
    port map (
            O => \N__11450\,
            I => \N__11429\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__11447\,
            I => \N__11424\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__11444\,
            I => \N__11424\
        );

    \I__2731\ : Sp12to4
    port map (
            O => \N__11437\,
            I => \N__11421\
        );

    \I__2730\ : Sp12to4
    port map (
            O => \N__11432\,
            I => \N__11418\
        );

    \I__2729\ : Span12Mux_h
    port map (
            O => \N__11429\,
            I => \N__11415\
        );

    \I__2728\ : Span12Mux_v
    port map (
            O => \N__11424\,
            I => \N__11412\
        );

    \I__2727\ : Span12Mux_v
    port map (
            O => \N__11421\,
            I => \N__11409\
        );

    \I__2726\ : Span12Mux_h
    port map (
            O => \N__11418\,
            I => \N__11406\
        );

    \I__2725\ : Span12Mux_v
    port map (
            O => \N__11415\,
            I => \N__11403\
        );

    \I__2724\ : Span12Mux_h
    port map (
            O => \N__11412\,
            I => \N__11400\
        );

    \I__2723\ : Span12Mux_h
    port map (
            O => \N__11409\,
            I => \N__11395\
        );

    \I__2722\ : Span12Mux_v
    port map (
            O => \N__11406\,
            I => \N__11395\
        );

    \I__2721\ : Odrv12
    port map (
            O => \N__11403\,
            I => \AGNUS_REV_c\
        );

    \I__2720\ : Odrv12
    port map (
            O => \N__11400\,
            I => \AGNUS_REV_c\
        );

    \I__2719\ : Odrv12
    port map (
            O => \N__11395\,
            I => \AGNUS_REV_c\
        );

    \I__2718\ : InMux
    port map (
            O => \N__11388\,
            I => \N__11385\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__11385\,
            I => \N__11382\
        );

    \I__2716\ : Span4Mux_v
    port map (
            O => \N__11382\,
            I => \N__11379\
        );

    \I__2715\ : Span4Mux_h
    port map (
            O => \N__11379\,
            I => \N__11376\
        );

    \I__2714\ : Odrv4
    port map (
            O => \N__11376\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2713\ : ClkMux
    port map (
            O => \N__11373\,
            I => \N__11355\
        );

    \I__2712\ : ClkMux
    port map (
            O => \N__11372\,
            I => \N__11355\
        );

    \I__2711\ : ClkMux
    port map (
            O => \N__11371\,
            I => \N__11355\
        );

    \I__2710\ : ClkMux
    port map (
            O => \N__11370\,
            I => \N__11355\
        );

    \I__2709\ : ClkMux
    port map (
            O => \N__11369\,
            I => \N__11355\
        );

    \I__2708\ : ClkMux
    port map (
            O => \N__11368\,
            I => \N__11355\
        );

    \I__2707\ : GlobalMux
    port map (
            O => \N__11355\,
            I => \N__11352\
        );

    \I__2706\ : gio2CtrlBuf
    port map (
            O => \N__11352\,
            I => \C3_c_g\
        );

    \I__2705\ : CEMux
    port map (
            O => \N__11349\,
            I => \N__11316\
        );

    \I__2704\ : CEMux
    port map (
            O => \N__11348\,
            I => \N__11316\
        );

    \I__2703\ : CEMux
    port map (
            O => \N__11347\,
            I => \N__11316\
        );

    \I__2702\ : CEMux
    port map (
            O => \N__11346\,
            I => \N__11316\
        );

    \I__2701\ : CEMux
    port map (
            O => \N__11345\,
            I => \N__11316\
        );

    \I__2700\ : CEMux
    port map (
            O => \N__11344\,
            I => \N__11316\
        );

    \I__2699\ : CEMux
    port map (
            O => \N__11343\,
            I => \N__11316\
        );

    \I__2698\ : CEMux
    port map (
            O => \N__11342\,
            I => \N__11316\
        );

    \I__2697\ : CEMux
    port map (
            O => \N__11341\,
            I => \N__11316\
        );

    \I__2696\ : CEMux
    port map (
            O => \N__11340\,
            I => \N__11316\
        );

    \I__2695\ : CEMux
    port map (
            O => \N__11339\,
            I => \N__11316\
        );

    \I__2694\ : GlobalMux
    port map (
            O => \N__11316\,
            I => \N__11313\
        );

    \I__2693\ : gio2CtrlBuf
    port map (
            O => \N__11313\,
            I => \DBRn_c_i_0_g\
        );

    \I__2692\ : InMux
    port map (
            O => \N__11310\,
            I => \N__11307\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__11307\,
            I => \N__11304\
        );

    \I__2690\ : Span4Mux_h
    port map (
            O => \N__11304\,
            I => \N__11301\
        );

    \I__2689\ : Odrv4
    port map (
            O => \N__11301\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\
        );

    \I__2688\ : CascadeMux
    port map (
            O => \N__11298\,
            I => \N__11295\
        );

    \I__2687\ : InMux
    port map (
            O => \N__11295\,
            I => \N__11289\
        );

    \I__2686\ : InMux
    port map (
            O => \N__11294\,
            I => \N__11286\
        );

    \I__2685\ : CascadeMux
    port map (
            O => \N__11293\,
            I => \N__11280\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__11292\,
            I => \N__11276\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__11289\,
            I => \N__11273\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__11286\,
            I => \N__11270\
        );

    \I__2681\ : CascadeMux
    port map (
            O => \N__11285\,
            I => \N__11266\
        );

    \I__2680\ : InMux
    port map (
            O => \N__11284\,
            I => \N__11262\
        );

    \I__2679\ : InMux
    port map (
            O => \N__11283\,
            I => \N__11257\
        );

    \I__2678\ : InMux
    port map (
            O => \N__11280\,
            I => \N__11257\
        );

    \I__2677\ : InMux
    port map (
            O => \N__11279\,
            I => \N__11250\
        );

    \I__2676\ : InMux
    port map (
            O => \N__11276\,
            I => \N__11247\
        );

    \I__2675\ : Span4Mux_h
    port map (
            O => \N__11273\,
            I => \N__11244\
        );

    \I__2674\ : Span12Mux_h
    port map (
            O => \N__11270\,
            I => \N__11241\
        );

    \I__2673\ : InMux
    port map (
            O => \N__11269\,
            I => \N__11238\
        );

    \I__2672\ : InMux
    port map (
            O => \N__11266\,
            I => \N__11233\
        );

    \I__2671\ : InMux
    port map (
            O => \N__11265\,
            I => \N__11233\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__11262\,
            I => \N__11228\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__11257\,
            I => \N__11228\
        );

    \I__2668\ : InMux
    port map (
            O => \N__11256\,
            I => \N__11219\
        );

    \I__2667\ : InMux
    port map (
            O => \N__11255\,
            I => \N__11219\
        );

    \I__2666\ : InMux
    port map (
            O => \N__11254\,
            I => \N__11219\
        );

    \I__2665\ : InMux
    port map (
            O => \N__11253\,
            I => \N__11219\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__11250\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__11247\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2662\ : Odrv4
    port map (
            O => \N__11244\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2661\ : Odrv12
    port map (
            O => \N__11241\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__11238\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__11233\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2658\ : Odrv4
    port map (
            O => \N__11228\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__11219\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2656\ : IoInMux
    port map (
            O => \N__11202\,
            I => \N__11199\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__11199\,
            I => \N__11196\
        );

    \I__2654\ : Span4Mux_s1_v
    port map (
            O => \N__11196\,
            I => \N__11193\
        );

    \I__2653\ : Sp12to4
    port map (
            O => \N__11193\,
            I => \N__11190\
        );

    \I__2652\ : Span12Mux_h
    port map (
            O => \N__11190\,
            I => \N__11187\
        );

    \I__2651\ : Span12Mux_v
    port map (
            O => \N__11187\,
            I => \N__11184\
        );

    \I__2650\ : Odrv12
    port map (
            O => \N__11184\,
            I => \ASn_c\
        );

    \I__2649\ : CEMux
    port map (
            O => \N__11181\,
            I => \N__11178\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__11178\,
            I => \U712_REG_SM.N_171_0\
        );

    \I__2647\ : InMux
    port map (
            O => \N__11175\,
            I => \N__11166\
        );

    \I__2646\ : InMux
    port map (
            O => \N__11174\,
            I => \N__11163\
        );

    \I__2645\ : InMux
    port map (
            O => \N__11173\,
            I => \N__11158\
        );

    \I__2644\ : InMux
    port map (
            O => \N__11172\,
            I => \N__11158\
        );

    \I__2643\ : InMux
    port map (
            O => \N__11171\,
            I => \N__11155\
        );

    \I__2642\ : InMux
    port map (
            O => \N__11170\,
            I => \N__11152\
        );

    \I__2641\ : InMux
    port map (
            O => \N__11169\,
            I => \N__11149\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__11166\,
            I => \N__11141\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__11163\,
            I => \N__11138\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__11158\,
            I => \N__11135\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__11155\,
            I => \N__11123\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__11152\,
            I => \N__11106\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__11149\,
            I => \N__11103\
        );

    \I__2634\ : SRMux
    port map (
            O => \N__11148\,
            I => \N__11001\
        );

    \I__2633\ : SRMux
    port map (
            O => \N__11147\,
            I => \N__11001\
        );

    \I__2632\ : SRMux
    port map (
            O => \N__11146\,
            I => \N__11001\
        );

    \I__2631\ : SRMux
    port map (
            O => \N__11145\,
            I => \N__11001\
        );

    \I__2630\ : SRMux
    port map (
            O => \N__11144\,
            I => \N__11001\
        );

    \I__2629\ : Glb2LocalMux
    port map (
            O => \N__11141\,
            I => \N__11001\
        );

    \I__2628\ : Glb2LocalMux
    port map (
            O => \N__11138\,
            I => \N__11001\
        );

    \I__2627\ : Glb2LocalMux
    port map (
            O => \N__11135\,
            I => \N__11001\
        );

    \I__2626\ : SRMux
    port map (
            O => \N__11134\,
            I => \N__11001\
        );

    \I__2625\ : SRMux
    port map (
            O => \N__11133\,
            I => \N__11001\
        );

    \I__2624\ : SRMux
    port map (
            O => \N__11132\,
            I => \N__11001\
        );

    \I__2623\ : SRMux
    port map (
            O => \N__11131\,
            I => \N__11001\
        );

    \I__2622\ : SRMux
    port map (
            O => \N__11130\,
            I => \N__11001\
        );

    \I__2621\ : SRMux
    port map (
            O => \N__11129\,
            I => \N__11001\
        );

    \I__2620\ : SRMux
    port map (
            O => \N__11128\,
            I => \N__11001\
        );

    \I__2619\ : SRMux
    port map (
            O => \N__11127\,
            I => \N__11001\
        );

    \I__2618\ : SRMux
    port map (
            O => \N__11126\,
            I => \N__11001\
        );

    \I__2617\ : Glb2LocalMux
    port map (
            O => \N__11123\,
            I => \N__11001\
        );

    \I__2616\ : SRMux
    port map (
            O => \N__11122\,
            I => \N__11001\
        );

    \I__2615\ : SRMux
    port map (
            O => \N__11121\,
            I => \N__11001\
        );

    \I__2614\ : SRMux
    port map (
            O => \N__11120\,
            I => \N__11001\
        );

    \I__2613\ : SRMux
    port map (
            O => \N__11119\,
            I => \N__11001\
        );

    \I__2612\ : SRMux
    port map (
            O => \N__11118\,
            I => \N__11001\
        );

    \I__2611\ : SRMux
    port map (
            O => \N__11117\,
            I => \N__11001\
        );

    \I__2610\ : SRMux
    port map (
            O => \N__11116\,
            I => \N__11001\
        );

    \I__2609\ : SRMux
    port map (
            O => \N__11115\,
            I => \N__11001\
        );

    \I__2608\ : SRMux
    port map (
            O => \N__11114\,
            I => \N__11001\
        );

    \I__2607\ : SRMux
    port map (
            O => \N__11113\,
            I => \N__11001\
        );

    \I__2606\ : SRMux
    port map (
            O => \N__11112\,
            I => \N__11001\
        );

    \I__2605\ : SRMux
    port map (
            O => \N__11111\,
            I => \N__11001\
        );

    \I__2604\ : SRMux
    port map (
            O => \N__11110\,
            I => \N__11001\
        );

    \I__2603\ : SRMux
    port map (
            O => \N__11109\,
            I => \N__11001\
        );

    \I__2602\ : Glb2LocalMux
    port map (
            O => \N__11106\,
            I => \N__11001\
        );

    \I__2601\ : Glb2LocalMux
    port map (
            O => \N__11103\,
            I => \N__11001\
        );

    \I__2600\ : SRMux
    port map (
            O => \N__11102\,
            I => \N__11001\
        );

    \I__2599\ : SRMux
    port map (
            O => \N__11101\,
            I => \N__11001\
        );

    \I__2598\ : SRMux
    port map (
            O => \N__11100\,
            I => \N__11001\
        );

    \I__2597\ : SRMux
    port map (
            O => \N__11099\,
            I => \N__11001\
        );

    \I__2596\ : SRMux
    port map (
            O => \N__11098\,
            I => \N__11001\
        );

    \I__2595\ : SRMux
    port map (
            O => \N__11097\,
            I => \N__11001\
        );

    \I__2594\ : SRMux
    port map (
            O => \N__11096\,
            I => \N__11001\
        );

    \I__2593\ : SRMux
    port map (
            O => \N__11095\,
            I => \N__11001\
        );

    \I__2592\ : SRMux
    port map (
            O => \N__11094\,
            I => \N__11001\
        );

    \I__2591\ : SRMux
    port map (
            O => \N__11093\,
            I => \N__11001\
        );

    \I__2590\ : SRMux
    port map (
            O => \N__11092\,
            I => \N__11001\
        );

    \I__2589\ : GlobalMux
    port map (
            O => \N__11001\,
            I => \N__10998\
        );

    \I__2588\ : gio2CtrlBuf
    port map (
            O => \N__10998\,
            I => \RESETn_c_i_g\
        );

    \I__2587\ : InMux
    port map (
            O => \N__10995\,
            I => \N__10992\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__10992\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__2585\ : CascadeMux
    port map (
            O => \N__10989\,
            I => \N__10982\
        );

    \I__2584\ : CascadeMux
    port map (
            O => \N__10988\,
            I => \N__10963\
        );

    \I__2583\ : CascadeMux
    port map (
            O => \N__10987\,
            I => \N__10960\
        );

    \I__2582\ : InMux
    port map (
            O => \N__10986\,
            I => \N__10955\
        );

    \I__2581\ : InMux
    port map (
            O => \N__10985\,
            I => \N__10952\
        );

    \I__2580\ : InMux
    port map (
            O => \N__10982\,
            I => \N__10941\
        );

    \I__2579\ : InMux
    port map (
            O => \N__10981\,
            I => \N__10941\
        );

    \I__2578\ : InMux
    port map (
            O => \N__10980\,
            I => \N__10941\
        );

    \I__2577\ : InMux
    port map (
            O => \N__10979\,
            I => \N__10941\
        );

    \I__2576\ : InMux
    port map (
            O => \N__10978\,
            I => \N__10941\
        );

    \I__2575\ : CascadeMux
    port map (
            O => \N__10977\,
            I => \N__10935\
        );

    \I__2574\ : InMux
    port map (
            O => \N__10976\,
            I => \N__10926\
        );

    \I__2573\ : InMux
    port map (
            O => \N__10975\,
            I => \N__10926\
        );

    \I__2572\ : InMux
    port map (
            O => \N__10974\,
            I => \N__10926\
        );

    \I__2571\ : InMux
    port map (
            O => \N__10973\,
            I => \N__10926\
        );

    \I__2570\ : InMux
    port map (
            O => \N__10972\,
            I => \N__10923\
        );

    \I__2569\ : InMux
    port map (
            O => \N__10971\,
            I => \N__10918\
        );

    \I__2568\ : InMux
    port map (
            O => \N__10970\,
            I => \N__10918\
        );

    \I__2567\ : InMux
    port map (
            O => \N__10969\,
            I => \N__10904\
        );

    \I__2566\ : InMux
    port map (
            O => \N__10968\,
            I => \N__10904\
        );

    \I__2565\ : InMux
    port map (
            O => \N__10967\,
            I => \N__10904\
        );

    \I__2564\ : InMux
    port map (
            O => \N__10966\,
            I => \N__10901\
        );

    \I__2563\ : InMux
    port map (
            O => \N__10963\,
            I => \N__10894\
        );

    \I__2562\ : InMux
    port map (
            O => \N__10960\,
            I => \N__10894\
        );

    \I__2561\ : InMux
    port map (
            O => \N__10959\,
            I => \N__10894\
        );

    \I__2560\ : InMux
    port map (
            O => \N__10958\,
            I => \N__10891\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__10955\,
            I => \N__10883\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__10952\,
            I => \N__10883\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__10941\,
            I => \N__10883\
        );

    \I__2556\ : InMux
    port map (
            O => \N__10940\,
            I => \N__10874\
        );

    \I__2555\ : InMux
    port map (
            O => \N__10939\,
            I => \N__10874\
        );

    \I__2554\ : InMux
    port map (
            O => \N__10938\,
            I => \N__10874\
        );

    \I__2553\ : InMux
    port map (
            O => \N__10935\,
            I => \N__10874\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__10926\,
            I => \N__10868\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__10923\,
            I => \N__10868\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__10918\,
            I => \N__10865\
        );

    \I__2549\ : InMux
    port map (
            O => \N__10917\,
            I => \N__10862\
        );

    \I__2548\ : InMux
    port map (
            O => \N__10916\,
            I => \N__10853\
        );

    \I__2547\ : InMux
    port map (
            O => \N__10915\,
            I => \N__10853\
        );

    \I__2546\ : InMux
    port map (
            O => \N__10914\,
            I => \N__10853\
        );

    \I__2545\ : InMux
    port map (
            O => \N__10913\,
            I => \N__10853\
        );

    \I__2544\ : InMux
    port map (
            O => \N__10912\,
            I => \N__10850\
        );

    \I__2543\ : InMux
    port map (
            O => \N__10911\,
            I => \N__10847\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__10904\,
            I => \N__10843\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__10901\,
            I => \N__10836\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__10894\,
            I => \N__10836\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__10891\,
            I => \N__10836\
        );

    \I__2538\ : InMux
    port map (
            O => \N__10890\,
            I => \N__10833\
        );

    \I__2537\ : Span4Mux_v
    port map (
            O => \N__10883\,
            I => \N__10828\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__10874\,
            I => \N__10828\
        );

    \I__2535\ : InMux
    port map (
            O => \N__10873\,
            I => \N__10825\
        );

    \I__2534\ : Span4Mux_v
    port map (
            O => \N__10868\,
            I => \N__10822\
        );

    \I__2533\ : Span4Mux_v
    port map (
            O => \N__10865\,
            I => \N__10811\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__10862\,
            I => \N__10811\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__10853\,
            I => \N__10811\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__10850\,
            I => \N__10811\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__10847\,
            I => \N__10811\
        );

    \I__2528\ : CascadeMux
    port map (
            O => \N__10846\,
            I => \N__10804\
        );

    \I__2527\ : Span4Mux_v
    port map (
            O => \N__10843\,
            I => \N__10799\
        );

    \I__2526\ : Span4Mux_v
    port map (
            O => \N__10836\,
            I => \N__10799\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__10833\,
            I => \N__10796\
        );

    \I__2524\ : Span4Mux_h
    port map (
            O => \N__10828\,
            I => \N__10791\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__10825\,
            I => \N__10791\
        );

    \I__2522\ : Span4Mux_h
    port map (
            O => \N__10822\,
            I => \N__10785\
        );

    \I__2521\ : Span4Mux_v
    port map (
            O => \N__10811\,
            I => \N__10785\
        );

    \I__2520\ : InMux
    port map (
            O => \N__10810\,
            I => \N__10782\
        );

    \I__2519\ : InMux
    port map (
            O => \N__10809\,
            I => \N__10777\
        );

    \I__2518\ : InMux
    port map (
            O => \N__10808\,
            I => \N__10777\
        );

    \I__2517\ : InMux
    port map (
            O => \N__10807\,
            I => \N__10774\
        );

    \I__2516\ : InMux
    port map (
            O => \N__10804\,
            I => \N__10771\
        );

    \I__2515\ : Span4Mux_h
    port map (
            O => \N__10799\,
            I => \N__10764\
        );

    \I__2514\ : Span4Mux_v
    port map (
            O => \N__10796\,
            I => \N__10764\
        );

    \I__2513\ : Span4Mux_v
    port map (
            O => \N__10791\,
            I => \N__10764\
        );

    \I__2512\ : InMux
    port map (
            O => \N__10790\,
            I => \N__10761\
        );

    \I__2511\ : Span4Mux_h
    port map (
            O => \N__10785\,
            I => \N__10758\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__10782\,
            I => \N__10753\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__10777\,
            I => \N__10753\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__10774\,
            I => \N__10744\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__10771\,
            I => \N__10744\
        );

    \I__2506\ : Sp12to4
    port map (
            O => \N__10764\,
            I => \N__10744\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__10761\,
            I => \N__10744\
        );

    \I__2504\ : Span4Mux_h
    port map (
            O => \N__10758\,
            I => \N__10739\
        );

    \I__2503\ : Span4Mux_v
    port map (
            O => \N__10753\,
            I => \N__10739\
        );

    \I__2502\ : Span12Mux_h
    port map (
            O => \N__10744\,
            I => \N__10734\
        );

    \I__2501\ : Sp12to4
    port map (
            O => \N__10739\,
            I => \N__10734\
        );

    \I__2500\ : Odrv12
    port map (
            O => \N__10734\,
            I => \RESETn_c\
        );

    \I__2499\ : InMux
    port map (
            O => \N__10731\,
            I => \N__10728\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__10728\,
            I => \N__10725\
        );

    \I__2497\ : Span12Mux_h
    port map (
            O => \N__10725\,
            I => \N__10722\
        );

    \I__2496\ : Odrv12
    port map (
            O => \N__10722\,
            I => \RAS1n_c\
        );

    \I__2495\ : InMux
    port map (
            O => \N__10719\,
            I => \N__10716\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__10716\,
            I => \N__10713\
        );

    \I__2493\ : Span4Mux_v
    port map (
            O => \N__10713\,
            I => \N__10709\
        );

    \I__2492\ : InMux
    port map (
            O => \N__10712\,
            I => \N__10706\
        );

    \I__2491\ : Sp12to4
    port map (
            O => \N__10709\,
            I => \N__10701\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__10706\,
            I => \N__10701\
        );

    \I__2489\ : Odrv12
    port map (
            O => \N__10701\,
            I => \RAS0n_c\
        );

    \I__2488\ : InMux
    port map (
            O => \N__10698\,
            I => \N__10695\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__10695\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2486\ : InMux
    port map (
            O => \N__10692\,
            I => \N__10689\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__10689\,
            I => \N__10645\
        );

    \I__2484\ : ClkMux
    port map (
            O => \N__10688\,
            I => \N__10536\
        );

    \I__2483\ : ClkMux
    port map (
            O => \N__10687\,
            I => \N__10536\
        );

    \I__2482\ : ClkMux
    port map (
            O => \N__10686\,
            I => \N__10536\
        );

    \I__2481\ : ClkMux
    port map (
            O => \N__10685\,
            I => \N__10536\
        );

    \I__2480\ : ClkMux
    port map (
            O => \N__10684\,
            I => \N__10536\
        );

    \I__2479\ : ClkMux
    port map (
            O => \N__10683\,
            I => \N__10536\
        );

    \I__2478\ : ClkMux
    port map (
            O => \N__10682\,
            I => \N__10536\
        );

    \I__2477\ : ClkMux
    port map (
            O => \N__10681\,
            I => \N__10536\
        );

    \I__2476\ : ClkMux
    port map (
            O => \N__10680\,
            I => \N__10536\
        );

    \I__2475\ : ClkMux
    port map (
            O => \N__10679\,
            I => \N__10536\
        );

    \I__2474\ : ClkMux
    port map (
            O => \N__10678\,
            I => \N__10536\
        );

    \I__2473\ : ClkMux
    port map (
            O => \N__10677\,
            I => \N__10536\
        );

    \I__2472\ : ClkMux
    port map (
            O => \N__10676\,
            I => \N__10536\
        );

    \I__2471\ : ClkMux
    port map (
            O => \N__10675\,
            I => \N__10536\
        );

    \I__2470\ : ClkMux
    port map (
            O => \N__10674\,
            I => \N__10536\
        );

    \I__2469\ : ClkMux
    port map (
            O => \N__10673\,
            I => \N__10536\
        );

    \I__2468\ : ClkMux
    port map (
            O => \N__10672\,
            I => \N__10536\
        );

    \I__2467\ : ClkMux
    port map (
            O => \N__10671\,
            I => \N__10536\
        );

    \I__2466\ : ClkMux
    port map (
            O => \N__10670\,
            I => \N__10536\
        );

    \I__2465\ : ClkMux
    port map (
            O => \N__10669\,
            I => \N__10536\
        );

    \I__2464\ : ClkMux
    port map (
            O => \N__10668\,
            I => \N__10536\
        );

    \I__2463\ : ClkMux
    port map (
            O => \N__10667\,
            I => \N__10536\
        );

    \I__2462\ : ClkMux
    port map (
            O => \N__10666\,
            I => \N__10536\
        );

    \I__2461\ : ClkMux
    port map (
            O => \N__10665\,
            I => \N__10536\
        );

    \I__2460\ : ClkMux
    port map (
            O => \N__10664\,
            I => \N__10536\
        );

    \I__2459\ : ClkMux
    port map (
            O => \N__10663\,
            I => \N__10536\
        );

    \I__2458\ : ClkMux
    port map (
            O => \N__10662\,
            I => \N__10536\
        );

    \I__2457\ : ClkMux
    port map (
            O => \N__10661\,
            I => \N__10536\
        );

    \I__2456\ : ClkMux
    port map (
            O => \N__10660\,
            I => \N__10536\
        );

    \I__2455\ : ClkMux
    port map (
            O => \N__10659\,
            I => \N__10536\
        );

    \I__2454\ : ClkMux
    port map (
            O => \N__10658\,
            I => \N__10536\
        );

    \I__2453\ : ClkMux
    port map (
            O => \N__10657\,
            I => \N__10536\
        );

    \I__2452\ : ClkMux
    port map (
            O => \N__10656\,
            I => \N__10536\
        );

    \I__2451\ : ClkMux
    port map (
            O => \N__10655\,
            I => \N__10536\
        );

    \I__2450\ : ClkMux
    port map (
            O => \N__10654\,
            I => \N__10536\
        );

    \I__2449\ : ClkMux
    port map (
            O => \N__10653\,
            I => \N__10536\
        );

    \I__2448\ : ClkMux
    port map (
            O => \N__10652\,
            I => \N__10536\
        );

    \I__2447\ : ClkMux
    port map (
            O => \N__10651\,
            I => \N__10536\
        );

    \I__2446\ : ClkMux
    port map (
            O => \N__10650\,
            I => \N__10536\
        );

    \I__2445\ : ClkMux
    port map (
            O => \N__10649\,
            I => \N__10536\
        );

    \I__2444\ : ClkMux
    port map (
            O => \N__10648\,
            I => \N__10536\
        );

    \I__2443\ : Glb2LocalMux
    port map (
            O => \N__10645\,
            I => \N__10536\
        );

    \I__2442\ : ClkMux
    port map (
            O => \N__10644\,
            I => \N__10536\
        );

    \I__2441\ : ClkMux
    port map (
            O => \N__10643\,
            I => \N__10536\
        );

    \I__2440\ : ClkMux
    port map (
            O => \N__10642\,
            I => \N__10536\
        );

    \I__2439\ : ClkMux
    port map (
            O => \N__10641\,
            I => \N__10536\
        );

    \I__2438\ : ClkMux
    port map (
            O => \N__10640\,
            I => \N__10536\
        );

    \I__2437\ : ClkMux
    port map (
            O => \N__10639\,
            I => \N__10536\
        );

    \I__2436\ : ClkMux
    port map (
            O => \N__10638\,
            I => \N__10536\
        );

    \I__2435\ : ClkMux
    port map (
            O => \N__10637\,
            I => \N__10536\
        );

    \I__2434\ : GlobalMux
    port map (
            O => \N__10536\,
            I => \CLK80_PLL\
        );

    \I__2433\ : InMux
    port map (
            O => \N__10533\,
            I => \N__10529\
        );

    \I__2432\ : InMux
    port map (
            O => \N__10532\,
            I => \N__10525\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__10529\,
            I => \N__10522\
        );

    \I__2430\ : InMux
    port map (
            O => \N__10528\,
            I => \N__10519\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__10525\,
            I => \N__10516\
        );

    \I__2428\ : Span4Mux_v
    port map (
            O => \N__10522\,
            I => \N__10512\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__10519\,
            I => \N__10509\
        );

    \I__2426\ : Span4Mux_v
    port map (
            O => \N__10516\,
            I => \N__10505\
        );

    \I__2425\ : InMux
    port map (
            O => \N__10515\,
            I => \N__10502\
        );

    \I__2424\ : Span4Mux_v
    port map (
            O => \N__10512\,
            I => \N__10499\
        );

    \I__2423\ : Span4Mux_v
    port map (
            O => \N__10509\,
            I => \N__10496\
        );

    \I__2422\ : InMux
    port map (
            O => \N__10508\,
            I => \N__10493\
        );

    \I__2421\ : Sp12to4
    port map (
            O => \N__10505\,
            I => \N__10490\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__10502\,
            I => \N__10487\
        );

    \I__2419\ : Sp12to4
    port map (
            O => \N__10499\,
            I => \N__10480\
        );

    \I__2418\ : Sp12to4
    port map (
            O => \N__10496\,
            I => \N__10480\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__10493\,
            I => \N__10480\
        );

    \I__2416\ : Span12Mux_h
    port map (
            O => \N__10490\,
            I => \N__10475\
        );

    \I__2415\ : Span12Mux_v
    port map (
            O => \N__10487\,
            I => \N__10475\
        );

    \I__2414\ : Span12Mux_h
    port map (
            O => \N__10480\,
            I => \N__10472\
        );

    \I__2413\ : Span12Mux_h
    port map (
            O => \N__10475\,
            I => \N__10469\
        );

    \I__2412\ : Span12Mux_v
    port map (
            O => \N__10472\,
            I => \N__10466\
        );

    \I__2411\ : Odrv12
    port map (
            O => \N__10469\,
            I => \RnW_c\
        );

    \I__2410\ : Odrv12
    port map (
            O => \N__10466\,
            I => \RnW_c\
        );

    \I__2409\ : InMux
    port map (
            O => \N__10461\,
            I => \N__10456\
        );

    \I__2408\ : InMux
    port map (
            O => \N__10460\,
            I => \N__10453\
        );

    \I__2407\ : InMux
    port map (
            O => \N__10459\,
            I => \N__10450\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__10456\,
            I => \N__10443\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__10453\,
            I => \N__10443\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__10450\,
            I => \N__10443\
        );

    \I__2403\ : Span4Mux_v
    port map (
            O => \N__10443\,
            I => \N__10439\
        );

    \I__2402\ : InMux
    port map (
            O => \N__10442\,
            I => \N__10436\
        );

    \I__2401\ : Span4Mux_v
    port map (
            O => \N__10439\,
            I => \N__10433\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__10436\,
            I => \N__10430\
        );

    \I__2399\ : Span4Mux_v
    port map (
            O => \N__10433\,
            I => \N__10425\
        );

    \I__2398\ : Span4Mux_h
    port map (
            O => \N__10430\,
            I => \N__10425\
        );

    \I__2397\ : Span4Mux_h
    port map (
            O => \N__10425\,
            I => \N__10421\
        );

    \I__2396\ : InMux
    port map (
            O => \N__10424\,
            I => \N__10417\
        );

    \I__2395\ : Span4Mux_h
    port map (
            O => \N__10421\,
            I => \N__10414\
        );

    \I__2394\ : InMux
    port map (
            O => \N__10420\,
            I => \N__10411\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__10417\,
            I => \N__10408\
        );

    \I__2392\ : Span4Mux_h
    port map (
            O => \N__10414\,
            I => \N__10403\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__10411\,
            I => \N__10403\
        );

    \I__2390\ : Span12Mux_h
    port map (
            O => \N__10408\,
            I => \N__10400\
        );

    \I__2389\ : Span4Mux_h
    port map (
            O => \N__10403\,
            I => \N__10397\
        );

    \I__2388\ : Span12Mux_v
    port map (
            O => \N__10400\,
            I => \N__10394\
        );

    \I__2387\ : Span4Mux_v
    port map (
            O => \N__10397\,
            I => \N__10391\
        );

    \I__2386\ : Odrv12
    port map (
            O => \N__10394\,
            I => \CASUn_c\
        );

    \I__2385\ : Odrv4
    port map (
            O => \N__10391\,
            I => \CASUn_c\
        );

    \I__2384\ : InMux
    port map (
            O => \N__10386\,
            I => \N__10383\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__10383\,
            I => \N__10380\
        );

    \I__2382\ : Span4Mux_h
    port map (
            O => \N__10380\,
            I => \N__10377\
        );

    \I__2381\ : Span4Mux_h
    port map (
            O => \N__10377\,
            I => \N__10374\
        );

    \I__2380\ : Odrv4
    port map (
            O => \N__10374\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2379\ : InMux
    port map (
            O => \N__10371\,
            I => \N__10367\
        );

    \I__2378\ : InMux
    port map (
            O => \N__10370\,
            I => \N__10364\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__10367\,
            I => \N__10359\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__10364\,
            I => \N__10359\
        );

    \I__2375\ : Span4Mux_v
    port map (
            O => \N__10359\,
            I => \N__10356\
        );

    \I__2374\ : Sp12to4
    port map (
            O => \N__10356\,
            I => \N__10353\
        );

    \I__2373\ : Span12Mux_h
    port map (
            O => \N__10353\,
            I => \N__10350\
        );

    \I__2372\ : Span12Mux_v
    port map (
            O => \N__10350\,
            I => \N__10347\
        );

    \I__2371\ : Odrv12
    port map (
            O => \N__10347\,
            I => \DRA_c_0\
        );

    \I__2370\ : InMux
    port map (
            O => \N__10344\,
            I => \N__10341\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__10341\,
            I => \N__10338\
        );

    \I__2368\ : Span4Mux_h
    port map (
            O => \N__10338\,
            I => \N__10335\
        );

    \I__2367\ : Odrv4
    port map (
            O => \N__10335\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__10332\,
            I => \N__10329\
        );

    \I__2365\ : InMux
    port map (
            O => \N__10329\,
            I => \N__10326\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__10326\,
            I => \N__10323\
        );

    \I__2363\ : Span4Mux_v
    port map (
            O => \N__10323\,
            I => \N__10320\
        );

    \I__2362\ : Odrv4
    port map (
            O => \N__10320\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2361\ : InMux
    port map (
            O => \N__10317\,
            I => \N__10312\
        );

    \I__2360\ : InMux
    port map (
            O => \N__10316\,
            I => \N__10309\
        );

    \I__2359\ : InMux
    port map (
            O => \N__10315\,
            I => \N__10305\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__10312\,
            I => \N__10300\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__10309\,
            I => \N__10300\
        );

    \I__2356\ : InMux
    port map (
            O => \N__10308\,
            I => \N__10297\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__10305\,
            I => \N__10290\
        );

    \I__2354\ : Sp12to4
    port map (
            O => \N__10300\,
            I => \N__10290\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__10297\,
            I => \N__10290\
        );

    \I__2352\ : Span12Mux_v
    port map (
            O => \N__10290\,
            I => \N__10287\
        );

    \I__2351\ : Span12Mux_h
    port map (
            O => \N__10287\,
            I => \N__10284\
        );

    \I__2350\ : Odrv12
    port map (
            O => \N__10284\,
            I => \DRA_c_6\
        );

    \I__2349\ : CascadeMux
    port map (
            O => \N__10281\,
            I => \N__10278\
        );

    \I__2348\ : InMux
    port map (
            O => \N__10278\,
            I => \N__10272\
        );

    \I__2347\ : InMux
    port map (
            O => \N__10277\,
            I => \N__10272\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__10272\,
            I => \N__10267\
        );

    \I__2345\ : InMux
    port map (
            O => \N__10271\,
            I => \N__10264\
        );

    \I__2344\ : InMux
    port map (
            O => \N__10270\,
            I => \N__10261\
        );

    \I__2343\ : Sp12to4
    port map (
            O => \N__10267\,
            I => \N__10254\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__10264\,
            I => \N__10254\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__10261\,
            I => \N__10254\
        );

    \I__2340\ : Span12Mux_v
    port map (
            O => \N__10254\,
            I => \N__10251\
        );

    \I__2339\ : Span12Mux_h
    port map (
            O => \N__10251\,
            I => \N__10248\
        );

    \I__2338\ : Odrv12
    port map (
            O => \N__10248\,
            I => \DRA_c_5\
        );

    \I__2337\ : InMux
    port map (
            O => \N__10245\,
            I => \N__10242\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__10242\,
            I => \N__10239\
        );

    \I__2335\ : Span4Mux_h
    port map (
            O => \N__10239\,
            I => \N__10236\
        );

    \I__2334\ : Odrv4
    port map (
            O => \N__10236\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2333\ : InMux
    port map (
            O => \N__10233\,
            I => \N__10230\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__10230\,
            I => \N__10227\
        );

    \I__2331\ : Span4Mux_h
    port map (
            O => \N__10227\,
            I => \N__10224\
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__10224\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__2329\ : InMux
    port map (
            O => \N__10221\,
            I => \N__10218\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__10218\,
            I => \N__10215\
        );

    \I__2327\ : Span4Mux_h
    port map (
            O => \N__10215\,
            I => \N__10212\
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__10212\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__2325\ : InMux
    port map (
            O => \N__10209\,
            I => \N__10203\
        );

    \I__2324\ : InMux
    port map (
            O => \N__10208\,
            I => \N__10200\
        );

    \I__2323\ : InMux
    port map (
            O => \N__10207\,
            I => \N__10197\
        );

    \I__2322\ : InMux
    port map (
            O => \N__10206\,
            I => \N__10194\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__10203\,
            I => \N__10191\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__10200\,
            I => \N__10184\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__10197\,
            I => \N__10184\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__10194\,
            I => \N__10184\
        );

    \I__2317\ : Span4Mux_v
    port map (
            O => \N__10191\,
            I => \N__10181\
        );

    \I__2316\ : Span4Mux_v
    port map (
            O => \N__10184\,
            I => \N__10178\
        );

    \I__2315\ : Sp12to4
    port map (
            O => \N__10181\,
            I => \N__10173\
        );

    \I__2314\ : Sp12to4
    port map (
            O => \N__10178\,
            I => \N__10173\
        );

    \I__2313\ : Span12Mux_h
    port map (
            O => \N__10173\,
            I => \N__10170\
        );

    \I__2312\ : Odrv12
    port map (
            O => \N__10170\,
            I => \DRA_c_8\
        );

    \I__2311\ : InMux
    port map (
            O => \N__10167\,
            I => \N__10164\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__10164\,
            I => \N__10161\
        );

    \I__2309\ : Span4Mux_v
    port map (
            O => \N__10161\,
            I => \N__10158\
        );

    \I__2308\ : Odrv4
    port map (
            O => \N__10158\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2307\ : InMux
    port map (
            O => \N__10155\,
            I => \N__10152\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__10152\,
            I => \N__10147\
        );

    \I__2305\ : InMux
    port map (
            O => \N__10151\,
            I => \N__10144\
        );

    \I__2304\ : InMux
    port map (
            O => \N__10150\,
            I => \N__10140\
        );

    \I__2303\ : Span4Mux_h
    port map (
            O => \N__10147\,
            I => \N__10135\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__10144\,
            I => \N__10135\
        );

    \I__2301\ : InMux
    port map (
            O => \N__10143\,
            I => \N__10132\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__10140\,
            I => \N__10129\
        );

    \I__2299\ : Span4Mux_v
    port map (
            O => \N__10135\,
            I => \N__10126\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__10132\,
            I => \N__10121\
        );

    \I__2297\ : Sp12to4
    port map (
            O => \N__10129\,
            I => \N__10121\
        );

    \I__2296\ : Span4Mux_v
    port map (
            O => \N__10126\,
            I => \N__10118\
        );

    \I__2295\ : Span12Mux_v
    port map (
            O => \N__10121\,
            I => \N__10113\
        );

    \I__2294\ : Sp12to4
    port map (
            O => \N__10118\,
            I => \N__10113\
        );

    \I__2293\ : Span12Mux_h
    port map (
            O => \N__10113\,
            I => \N__10110\
        );

    \I__2292\ : Odrv12
    port map (
            O => \N__10110\,
            I => \DRA_c_3\
        );

    \I__2291\ : InMux
    port map (
            O => \N__10107\,
            I => \N__10102\
        );

    \I__2290\ : InMux
    port map (
            O => \N__10106\,
            I => \N__10099\
        );

    \I__2289\ : InMux
    port map (
            O => \N__10105\,
            I => \N__10096\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__10102\,
            I => \N__10092\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__10099\,
            I => \N__10089\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__10096\,
            I => \N__10086\
        );

    \I__2285\ : InMux
    port map (
            O => \N__10095\,
            I => \N__10083\
        );

    \I__2284\ : Span4Mux_v
    port map (
            O => \N__10092\,
            I => \N__10080\
        );

    \I__2283\ : Span4Mux_v
    port map (
            O => \N__10089\,
            I => \N__10077\
        );

    \I__2282\ : Span4Mux_h
    port map (
            O => \N__10086\,
            I => \N__10074\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__10083\,
            I => \N__10071\
        );

    \I__2280\ : Span4Mux_v
    port map (
            O => \N__10080\,
            I => \N__10068\
        );

    \I__2279\ : Span4Mux_v
    port map (
            O => \N__10077\,
            I => \N__10065\
        );

    \I__2278\ : Sp12to4
    port map (
            O => \N__10074\,
            I => \N__10060\
        );

    \I__2277\ : Sp12to4
    port map (
            O => \N__10071\,
            I => \N__10060\
        );

    \I__2276\ : Sp12to4
    port map (
            O => \N__10068\,
            I => \N__10057\
        );

    \I__2275\ : Sp12to4
    port map (
            O => \N__10065\,
            I => \N__10052\
        );

    \I__2274\ : Span12Mux_v
    port map (
            O => \N__10060\,
            I => \N__10052\
        );

    \I__2273\ : Span12Mux_h
    port map (
            O => \N__10057\,
            I => \N__10049\
        );

    \I__2272\ : Span12Mux_h
    port map (
            O => \N__10052\,
            I => \N__10046\
        );

    \I__2271\ : Odrv12
    port map (
            O => \N__10049\,
            I => \DRA_c_4\
        );

    \I__2270\ : Odrv12
    port map (
            O => \N__10046\,
            I => \DRA_c_4\
        );

    \I__2269\ : InMux
    port map (
            O => \N__10041\,
            I => \N__10038\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__10038\,
            I => \N__10035\
        );

    \I__2267\ : Span4Mux_h
    port map (
            O => \N__10035\,
            I => \N__10032\
        );

    \I__2266\ : Odrv4
    port map (
            O => \N__10032\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2265\ : InMux
    port map (
            O => \N__10029\,
            I => \N__10025\
        );

    \I__2264\ : InMux
    port map (
            O => \N__10028\,
            I => \N__10022\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__10025\,
            I => \N__10017\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__10022\,
            I => \N__10014\
        );

    \I__2261\ : InMux
    port map (
            O => \N__10021\,
            I => \N__10011\
        );

    \I__2260\ : InMux
    port map (
            O => \N__10020\,
            I => \N__10008\
        );

    \I__2259\ : Span4Mux_v
    port map (
            O => \N__10017\,
            I => \N__10005\
        );

    \I__2258\ : Span4Mux_v
    port map (
            O => \N__10014\,
            I => \N__10002\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__10011\,
            I => \N__9997\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__10008\,
            I => \N__9997\
        );

    \I__2255\ : Sp12to4
    port map (
            O => \N__10005\,
            I => \N__9994\
        );

    \I__2254\ : Span4Mux_v
    port map (
            O => \N__10002\,
            I => \N__9991\
        );

    \I__2253\ : Span4Mux_h
    port map (
            O => \N__9997\,
            I => \N__9988\
        );

    \I__2252\ : Span12Mux_h
    port map (
            O => \N__9994\,
            I => \N__9985\
        );

    \I__2251\ : Span4Mux_v
    port map (
            O => \N__9991\,
            I => \N__9982\
        );

    \I__2250\ : Sp12to4
    port map (
            O => \N__9988\,
            I => \N__9979\
        );

    \I__2249\ : Span12Mux_v
    port map (
            O => \N__9985\,
            I => \N__9976\
        );

    \I__2248\ : Sp12to4
    port map (
            O => \N__9982\,
            I => \N__9971\
        );

    \I__2247\ : Span12Mux_v
    port map (
            O => \N__9979\,
            I => \N__9971\
        );

    \I__2246\ : Odrv12
    port map (
            O => \N__9976\,
            I => \DRA_c_2\
        );

    \I__2245\ : Odrv12
    port map (
            O => \N__9971\,
            I => \DRA_c_2\
        );

    \I__2244\ : InMux
    port map (
            O => \N__9966\,
            I => \N__9961\
        );

    \I__2243\ : InMux
    port map (
            O => \N__9965\,
            I => \N__9958\
        );

    \I__2242\ : InMux
    port map (
            O => \N__9964\,
            I => \N__9955\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__9961\,
            I => \N__9952\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__9958\,
            I => \N__9949\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__9955\,
            I => \N__9945\
        );

    \I__2238\ : Span4Mux_v
    port map (
            O => \N__9952\,
            I => \N__9942\
        );

    \I__2237\ : Span4Mux_v
    port map (
            O => \N__9949\,
            I => \N__9939\
        );

    \I__2236\ : InMux
    port map (
            O => \N__9948\,
            I => \N__9936\
        );

    \I__2235\ : Sp12to4
    port map (
            O => \N__9945\,
            I => \N__9933\
        );

    \I__2234\ : Sp12to4
    port map (
            O => \N__9942\,
            I => \N__9926\
        );

    \I__2233\ : Sp12to4
    port map (
            O => \N__9939\,
            I => \N__9926\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__9936\,
            I => \N__9926\
        );

    \I__2231\ : Span12Mux_v
    port map (
            O => \N__9933\,
            I => \N__9923\
        );

    \I__2230\ : Span12Mux_h
    port map (
            O => \N__9926\,
            I => \N__9920\
        );

    \I__2229\ : Span12Mux_h
    port map (
            O => \N__9923\,
            I => \N__9915\
        );

    \I__2228\ : Span12Mux_v
    port map (
            O => \N__9920\,
            I => \N__9915\
        );

    \I__2227\ : Odrv12
    port map (
            O => \N__9915\,
            I => \DRA_c_1\
        );

    \I__2226\ : InMux
    port map (
            O => \N__9912\,
            I => \N__9909\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__9909\,
            I => \N__9906\
        );

    \I__2224\ : Span4Mux_h
    port map (
            O => \N__9906\,
            I => \N__9903\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__9903\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__2222\ : InMux
    port map (
            O => \N__9900\,
            I => \N__9897\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__9897\,
            I => \N__9894\
        );

    \I__2220\ : Span4Mux_h
    port map (
            O => \N__9894\,
            I => \N__9891\
        );

    \I__2219\ : Odrv4
    port map (
            O => \N__9891\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2218\ : CascadeMux
    port map (
            O => \N__9888\,
            I => \N__9885\
        );

    \I__2217\ : InMux
    port map (
            O => \N__9885\,
            I => \N__9882\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__9882\,
            I => \N__9879\
        );

    \I__2215\ : Span4Mux_v
    port map (
            O => \N__9879\,
            I => \N__9875\
        );

    \I__2214\ : InMux
    port map (
            O => \N__9878\,
            I => \N__9872\
        );

    \I__2213\ : Span4Mux_h
    port map (
            O => \N__9875\,
            I => \N__9869\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__9872\,
            I => \N__9866\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__9869\,
            I => \DBRn_c_i\
        );

    \I__2210\ : Odrv4
    port map (
            O => \N__9866\,
            I => \DBRn_c_i\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__9861\,
            I => \N__9858\
        );

    \I__2208\ : InMux
    port map (
            O => \N__9858\,
            I => \N__9854\
        );

    \I__2207\ : InMux
    port map (
            O => \N__9857\,
            I => \N__9851\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__9854\,
            I => \N__9848\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__9851\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__2204\ : Odrv4
    port map (
            O => \N__9848\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__2203\ : InMux
    port map (
            O => \N__9843\,
            I => \N__9840\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__9840\,
            I => \N__9834\
        );

    \I__2201\ : InMux
    port map (
            O => \N__9839\,
            I => \N__9828\
        );

    \I__2200\ : InMux
    port map (
            O => \N__9838\,
            I => \N__9828\
        );

    \I__2199\ : InMux
    port map (
            O => \N__9837\,
            I => \N__9825\
        );

    \I__2198\ : Span4Mux_h
    port map (
            O => \N__9834\,
            I => \N__9821\
        );

    \I__2197\ : InMux
    port map (
            O => \N__9833\,
            I => \N__9818\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__9828\,
            I => \N__9813\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__9825\,
            I => \N__9813\
        );

    \I__2194\ : InMux
    port map (
            O => \N__9824\,
            I => \N__9810\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__9821\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__9818\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2191\ : Odrv4
    port map (
            O => \N__9813\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__9810\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2189\ : IoInMux
    port map (
            O => \N__9801\,
            I => \N__9798\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__9798\,
            I => \N__9795\
        );

    \I__2187\ : IoSpan4Mux
    port map (
            O => \N__9795\,
            I => \N__9792\
        );

    \I__2186\ : Sp12to4
    port map (
            O => \N__9792\,
            I => \N__9789\
        );

    \I__2185\ : Span12Mux_s9_v
    port map (
            O => \N__9789\,
            I => \N__9786\
        );

    \I__2184\ : Odrv12
    port map (
            O => \N__9786\,
            I => \RASn_c\
        );

    \I__2183\ : InMux
    port map (
            O => \N__9783\,
            I => \N__9780\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__9780\,
            I => \N__9777\
        );

    \I__2181\ : Span4Mux_v
    port map (
            O => \N__9777\,
            I => \N__9774\
        );

    \I__2180\ : Odrv4
    port map (
            O => \N__9774\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__2179\ : InMux
    port map (
            O => \N__9771\,
            I => \N__9768\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__9768\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2177\ : InMux
    port map (
            O => \N__9765\,
            I => \N__9757\
        );

    \I__2176\ : InMux
    port map (
            O => \N__9764\,
            I => \N__9757\
        );

    \I__2175\ : InMux
    port map (
            O => \N__9763\,
            I => \N__9754\
        );

    \I__2174\ : InMux
    port map (
            O => \N__9762\,
            I => \N__9751\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__9757\,
            I => \N__9748\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__9754\,
            I => \N__9743\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__9751\,
            I => \N__9743\
        );

    \I__2170\ : Span4Mux_v
    port map (
            O => \N__9748\,
            I => \N__9740\
        );

    \I__2169\ : Span4Mux_v
    port map (
            O => \N__9743\,
            I => \N__9737\
        );

    \I__2168\ : Sp12to4
    port map (
            O => \N__9740\,
            I => \N__9732\
        );

    \I__2167\ : Sp12to4
    port map (
            O => \N__9737\,
            I => \N__9732\
        );

    \I__2166\ : Span12Mux_h
    port map (
            O => \N__9732\,
            I => \N__9729\
        );

    \I__2165\ : Odrv12
    port map (
            O => \N__9729\,
            I => \DRA_c_7\
        );

    \I__2164\ : InMux
    port map (
            O => \N__9726\,
            I => \N__9723\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__9723\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2162\ : InMux
    port map (
            O => \N__9720\,
            I => \N__9717\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__9717\,
            I => \N__9714\
        );

    \I__2160\ : Span4Mux_v
    port map (
            O => \N__9714\,
            I => \N__9711\
        );

    \I__2159\ : Odrv4
    port map (
            O => \N__9711\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__2158\ : InMux
    port map (
            O => \N__9708\,
            I => \N__9705\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__9705\,
            I => \U712_CHIP_RAM.CMA_5_i_0_9\
        );

    \I__2156\ : InMux
    port map (
            O => \N__9702\,
            I => \N__9699\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__9699\,
            I => \N__9696\
        );

    \I__2154\ : Span4Mux_v
    port map (
            O => \N__9696\,
            I => \N__9693\
        );

    \I__2153\ : Span4Mux_v
    port map (
            O => \N__9693\,
            I => \N__9690\
        );

    \I__2152\ : Sp12to4
    port map (
            O => \N__9690\,
            I => \N__9687\
        );

    \I__2151\ : Span12Mux_h
    port map (
            O => \N__9687\,
            I => \N__9684\
        );

    \I__2150\ : Odrv12
    port map (
            O => \N__9684\,
            I => \A_c_19\
        );

    \I__2149\ : CascadeMux
    port map (
            O => \N__9681\,
            I => \N__9672\
        );

    \I__2148\ : CascadeMux
    port map (
            O => \N__9680\,
            I => \N__9666\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9679\,
            I => \N__9657\
        );

    \I__2146\ : InMux
    port map (
            O => \N__9678\,
            I => \N__9657\
        );

    \I__2145\ : InMux
    port map (
            O => \N__9677\,
            I => \N__9657\
        );

    \I__2144\ : InMux
    port map (
            O => \N__9676\,
            I => \N__9652\
        );

    \I__2143\ : InMux
    port map (
            O => \N__9675\,
            I => \N__9652\
        );

    \I__2142\ : InMux
    port map (
            O => \N__9672\,
            I => \N__9648\
        );

    \I__2141\ : InMux
    port map (
            O => \N__9671\,
            I => \N__9645\
        );

    \I__2140\ : InMux
    port map (
            O => \N__9670\,
            I => \N__9636\
        );

    \I__2139\ : InMux
    port map (
            O => \N__9669\,
            I => \N__9636\
        );

    \I__2138\ : InMux
    port map (
            O => \N__9666\,
            I => \N__9636\
        );

    \I__2137\ : InMux
    port map (
            O => \N__9665\,
            I => \N__9636\
        );

    \I__2136\ : InMux
    port map (
            O => \N__9664\,
            I => \N__9626\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__9657\,
            I => \N__9621\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__9652\,
            I => \N__9621\
        );

    \I__2133\ : InMux
    port map (
            O => \N__9651\,
            I => \N__9618\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__9648\,
            I => \N__9613\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__9645\,
            I => \N__9613\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__9636\,
            I => \N__9610\
        );

    \I__2129\ : InMux
    port map (
            O => \N__9635\,
            I => \N__9607\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9634\,
            I => \N__9603\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9633\,
            I => \N__9600\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9632\,
            I => \N__9592\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9631\,
            I => \N__9592\
        );

    \I__2124\ : InMux
    port map (
            O => \N__9630\,
            I => \N__9592\
        );

    \I__2123\ : InMux
    port map (
            O => \N__9629\,
            I => \N__9589\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__9626\,
            I => \N__9586\
        );

    \I__2121\ : Span4Mux_v
    port map (
            O => \N__9621\,
            I => \N__9577\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__9618\,
            I => \N__9577\
        );

    \I__2119\ : Span4Mux_v
    port map (
            O => \N__9613\,
            I => \N__9577\
        );

    \I__2118\ : Span4Mux_v
    port map (
            O => \N__9610\,
            I => \N__9577\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__9607\,
            I => \N__9574\
        );

    \I__2116\ : InMux
    port map (
            O => \N__9606\,
            I => \N__9571\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__9603\,
            I => \N__9566\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__9600\,
            I => \N__9566\
        );

    \I__2113\ : InMux
    port map (
            O => \N__9599\,
            I => \N__9561\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__9592\,
            I => \N__9556\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__9589\,
            I => \N__9556\
        );

    \I__2110\ : Span4Mux_v
    port map (
            O => \N__9586\,
            I => \N__9551\
        );

    \I__2109\ : Span4Mux_h
    port map (
            O => \N__9577\,
            I => \N__9551\
        );

    \I__2108\ : Span4Mux_v
    port map (
            O => \N__9574\,
            I => \N__9544\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__9571\,
            I => \N__9544\
        );

    \I__2106\ : Span4Mux_v
    port map (
            O => \N__9566\,
            I => \N__9544\
        );

    \I__2105\ : InMux
    port map (
            O => \N__9565\,
            I => \N__9539\
        );

    \I__2104\ : InMux
    port map (
            O => \N__9564\,
            I => \N__9539\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__9561\,
            I => \CPU_CYCLEm\
        );

    \I__2102\ : Odrv12
    port map (
            O => \N__9556\,
            I => \CPU_CYCLEm\
        );

    \I__2101\ : Odrv4
    port map (
            O => \N__9551\,
            I => \CPU_CYCLEm\
        );

    \I__2100\ : Odrv4
    port map (
            O => \N__9544\,
            I => \CPU_CYCLEm\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__9539\,
            I => \CPU_CYCLEm\
        );

    \I__2098\ : IoInMux
    port map (
            O => \N__9528\,
            I => \N__9525\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__9525\,
            I => \N__9522\
        );

    \I__2096\ : IoSpan4Mux
    port map (
            O => \N__9522\,
            I => \N__9519\
        );

    \I__2095\ : IoSpan4Mux
    port map (
            O => \N__9519\,
            I => \N__9516\
        );

    \I__2094\ : Span4Mux_s2_h
    port map (
            O => \N__9516\,
            I => \N__9513\
        );

    \I__2093\ : Sp12to4
    port map (
            O => \N__9513\,
            I => \N__9510\
        );

    \I__2092\ : Odrv12
    port map (
            O => \N__9510\,
            I => \CMA_c_9\
        );

    \I__2091\ : InMux
    port map (
            O => \N__9507\,
            I => \N__9504\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__9504\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__2089\ : IoInMux
    port map (
            O => \N__9501\,
            I => \N__9498\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__9498\,
            I => \N__9495\
        );

    \I__2087\ : IoSpan4Mux
    port map (
            O => \N__9495\,
            I => \N__9492\
        );

    \I__2086\ : Sp12to4
    port map (
            O => \N__9492\,
            I => \N__9489\
        );

    \I__2085\ : Span12Mux_s7_h
    port map (
            O => \N__9489\,
            I => \N__9486\
        );

    \I__2084\ : Span12Mux_v
    port map (
            O => \N__9486\,
            I => \N__9483\
        );

    \I__2083\ : Odrv12
    port map (
            O => \N__9483\,
            I => \CMA_c_3\
        );

    \I__2082\ : InMux
    port map (
            O => \N__9480\,
            I => \N__9477\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__9477\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__2080\ : IoInMux
    port map (
            O => \N__9474\,
            I => \N__9471\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__9471\,
            I => \N__9468\
        );

    \I__2078\ : Span4Mux_s3_h
    port map (
            O => \N__9468\,
            I => \N__9465\
        );

    \I__2077\ : Sp12to4
    port map (
            O => \N__9465\,
            I => \N__9462\
        );

    \I__2076\ : Span12Mux_s9_v
    port map (
            O => \N__9462\,
            I => \N__9459\
        );

    \I__2075\ : Span12Mux_h
    port map (
            O => \N__9459\,
            I => \N__9456\
        );

    \I__2074\ : Odrv12
    port map (
            O => \N__9456\,
            I => \CMA_c_4\
        );

    \I__2073\ : InMux
    port map (
            O => \N__9453\,
            I => \N__9450\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__9450\,
            I => \N__9447\
        );

    \I__2071\ : Odrv4
    port map (
            O => \N__9447\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__2070\ : IoInMux
    port map (
            O => \N__9444\,
            I => \N__9441\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__9441\,
            I => \N__9438\
        );

    \I__2068\ : IoSpan4Mux
    port map (
            O => \N__9438\,
            I => \N__9435\
        );

    \I__2067\ : IoSpan4Mux
    port map (
            O => \N__9435\,
            I => \N__9432\
        );

    \I__2066\ : Span4Mux_s2_h
    port map (
            O => \N__9432\,
            I => \N__9429\
        );

    \I__2065\ : Sp12to4
    port map (
            O => \N__9429\,
            I => \N__9426\
        );

    \I__2064\ : Span12Mux_h
    port map (
            O => \N__9426\,
            I => \N__9423\
        );

    \I__2063\ : Odrv12
    port map (
            O => \N__9423\,
            I => \CMA_c_6\
        );

    \I__2062\ : CascadeMux
    port map (
            O => \N__9420\,
            I => \N__9417\
        );

    \I__2061\ : InMux
    port map (
            O => \N__9417\,
            I => \N__9414\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__9414\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__2059\ : IoInMux
    port map (
            O => \N__9411\,
            I => \N__9408\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__9408\,
            I => \N__9405\
        );

    \I__2057\ : Span4Mux_s3_h
    port map (
            O => \N__9405\,
            I => \N__9402\
        );

    \I__2056\ : Sp12to4
    port map (
            O => \N__9402\,
            I => \N__9399\
        );

    \I__2055\ : Span12Mux_s11_v
    port map (
            O => \N__9399\,
            I => \N__9396\
        );

    \I__2054\ : Span12Mux_h
    port map (
            O => \N__9396\,
            I => \N__9393\
        );

    \I__2053\ : Odrv12
    port map (
            O => \N__9393\,
            I => \CMA_c_7\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__9390\,
            I => \N__9381\
        );

    \I__2051\ : CascadeMux
    port map (
            O => \N__9389\,
            I => \N__9378\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__9388\,
            I => \N__9375\
        );

    \I__2049\ : InMux
    port map (
            O => \N__9387\,
            I => \N__9369\
        );

    \I__2048\ : InMux
    port map (
            O => \N__9386\,
            I => \N__9358\
        );

    \I__2047\ : InMux
    port map (
            O => \N__9385\,
            I => \N__9358\
        );

    \I__2046\ : InMux
    port map (
            O => \N__9384\,
            I => \N__9358\
        );

    \I__2045\ : InMux
    port map (
            O => \N__9381\,
            I => \N__9358\
        );

    \I__2044\ : InMux
    port map (
            O => \N__9378\,
            I => \N__9358\
        );

    \I__2043\ : InMux
    port map (
            O => \N__9375\,
            I => \N__9355\
        );

    \I__2042\ : InMux
    port map (
            O => \N__9374\,
            I => \N__9352\
        );

    \I__2041\ : InMux
    port map (
            O => \N__9373\,
            I => \N__9349\
        );

    \I__2040\ : InMux
    port map (
            O => \N__9372\,
            I => \N__9346\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__9369\,
            I => \U712_CHIP_RAM.N_330\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__9358\,
            I => \U712_CHIP_RAM.N_330\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__9355\,
            I => \U712_CHIP_RAM.N_330\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__9352\,
            I => \U712_CHIP_RAM.N_330\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__9349\,
            I => \U712_CHIP_RAM.N_330\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__9346\,
            I => \U712_CHIP_RAM.N_330\
        );

    \I__2033\ : InMux
    port map (
            O => \N__9333\,
            I => \N__9329\
        );

    \I__2032\ : InMux
    port map (
            O => \N__9332\,
            I => \N__9326\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__9329\,
            I => \N__9318\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__9326\,
            I => \N__9315\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9325\,
            I => \N__9308\
        );

    \I__2028\ : InMux
    port map (
            O => \N__9324\,
            I => \N__9308\
        );

    \I__2027\ : InMux
    port map (
            O => \N__9323\,
            I => \N__9308\
        );

    \I__2026\ : InMux
    port map (
            O => \N__9322\,
            I => \N__9303\
        );

    \I__2025\ : InMux
    port map (
            O => \N__9321\,
            I => \N__9303\
        );

    \I__2024\ : Odrv4
    port map (
            O => \N__9318\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__9315\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__9308\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__9303\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__2020\ : CascadeMux
    port map (
            O => \N__9294\,
            I => \N__9291\
        );

    \I__2019\ : InMux
    port map (
            O => \N__9291\,
            I => \N__9288\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__9288\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\
        );

    \I__2017\ : IoInMux
    port map (
            O => \N__9285\,
            I => \N__9282\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__9282\,
            I => \N__9279\
        );

    \I__2015\ : Span4Mux_s3_h
    port map (
            O => \N__9279\,
            I => \N__9276\
        );

    \I__2014\ : Sp12to4
    port map (
            O => \N__9276\,
            I => \N__9273\
        );

    \I__2013\ : Span12Mux_v
    port map (
            O => \N__9273\,
            I => \N__9270\
        );

    \I__2012\ : Span12Mux_h
    port map (
            O => \N__9270\,
            I => \N__9267\
        );

    \I__2011\ : Odrv12
    port map (
            O => \N__9267\,
            I => \CMA_c_8\
        );

    \I__2010\ : CEMux
    port map (
            O => \N__9264\,
            I => \N__9257\
        );

    \I__2009\ : CEMux
    port map (
            O => \N__9263\,
            I => \N__9254\
        );

    \I__2008\ : CEMux
    port map (
            O => \N__9262\,
            I => \N__9251\
        );

    \I__2007\ : CEMux
    port map (
            O => \N__9261\,
            I => \N__9248\
        );

    \I__2006\ : CEMux
    port map (
            O => \N__9260\,
            I => \N__9245\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__9257\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__9254\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__9251\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__9248\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__9245\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__2000\ : InMux
    port map (
            O => \N__9234\,
            I => \N__9231\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__9231\,
            I => \N__9228\
        );

    \I__1998\ : Span4Mux_h
    port map (
            O => \N__9228\,
            I => \N__9225\
        );

    \I__1997\ : Odrv4
    port map (
            O => \N__9225\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1996\ : InMux
    port map (
            O => \N__9222\,
            I => \N__9219\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__9219\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__1994\ : InMux
    port map (
            O => \N__9216\,
            I => \N__9213\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__9213\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__1992\ : InMux
    port map (
            O => \N__9210\,
            I => \N__9207\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__9207\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\
        );

    \I__1990\ : InMux
    port map (
            O => \N__9204\,
            I => \N__9198\
        );

    \I__1989\ : InMux
    port map (
            O => \N__9203\,
            I => \N__9198\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__9198\,
            I => \N__9195\
        );

    \I__1987\ : Odrv4
    port map (
            O => \N__9195\,
            I => \N_322\
        );

    \I__1986\ : IoInMux
    port map (
            O => \N__9192\,
            I => \N__9189\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__9189\,
            I => \N__9186\
        );

    \I__1984\ : Span12Mux_s5_v
    port map (
            O => \N__9186\,
            I => \N__9183\
        );

    \I__1983\ : Odrv12
    port map (
            O => \N__9183\,
            I => \RESETn_c_i\
        );

    \I__1982\ : IoInMux
    port map (
            O => \N__9180\,
            I => \N__9177\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__9177\,
            I => \N__9174\
        );

    \I__1980\ : Span12Mux_s7_v
    port map (
            O => \N__9174\,
            I => \N__9171\
        );

    \I__1979\ : Odrv12
    port map (
            O => \N__9171\,
            I => \N_342_i\
        );

    \I__1978\ : IoInMux
    port map (
            O => \N__9168\,
            I => \N__9165\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__9165\,
            I => \N__9162\
        );

    \I__1976\ : Span4Mux_s2_v
    port map (
            O => \N__9162\,
            I => \N__9159\
        );

    \I__1975\ : Span4Mux_v
    port map (
            O => \N__9159\,
            I => \N__9156\
        );

    \I__1974\ : Odrv4
    port map (
            O => \N__9156\,
            I => \N_345_i\
        );

    \I__1973\ : InMux
    port map (
            O => \N__9153\,
            I => \N__9145\
        );

    \I__1972\ : InMux
    port map (
            O => \N__9152\,
            I => \N__9141\
        );

    \I__1971\ : InMux
    port map (
            O => \N__9151\,
            I => \N__9136\
        );

    \I__1970\ : InMux
    port map (
            O => \N__9150\,
            I => \N__9136\
        );

    \I__1969\ : InMux
    port map (
            O => \N__9149\,
            I => \N__9132\
        );

    \I__1968\ : CascadeMux
    port map (
            O => \N__9148\,
            I => \N__9129\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__9145\,
            I => \N__9126\
        );

    \I__1966\ : InMux
    port map (
            O => \N__9144\,
            I => \N__9123\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__9141\,
            I => \N__9120\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__9136\,
            I => \N__9117\
        );

    \I__1963\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9114\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__9132\,
            I => \N__9111\
        );

    \I__1961\ : InMux
    port map (
            O => \N__9129\,
            I => \N__9108\
        );

    \I__1960\ : Span4Mux_v
    port map (
            O => \N__9126\,
            I => \N__9105\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__9123\,
            I => \N__9102\
        );

    \I__1958\ : Span4Mux_v
    port map (
            O => \N__9120\,
            I => \N__9095\
        );

    \I__1957\ : Span4Mux_h
    port map (
            O => \N__9117\,
            I => \N__9095\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__9114\,
            I => \N__9095\
        );

    \I__1955\ : Span4Mux_v
    port map (
            O => \N__9111\,
            I => \N__9092\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__9108\,
            I => \N__9089\
        );

    \I__1953\ : Span4Mux_h
    port map (
            O => \N__9105\,
            I => \N__9084\
        );

    \I__1952\ : Span4Mux_v
    port map (
            O => \N__9102\,
            I => \N__9084\
        );

    \I__1951\ : Span4Mux_h
    port map (
            O => \N__9095\,
            I => \N__9081\
        );

    \I__1950\ : Sp12to4
    port map (
            O => \N__9092\,
            I => \N__9074\
        );

    \I__1949\ : Span12Mux_h
    port map (
            O => \N__9089\,
            I => \N__9074\
        );

    \I__1948\ : Sp12to4
    port map (
            O => \N__9084\,
            I => \N__9074\
        );

    \I__1947\ : Span4Mux_v
    port map (
            O => \N__9081\,
            I => \N__9071\
        );

    \I__1946\ : Span12Mux_h
    port map (
            O => \N__9074\,
            I => \N__9068\
        );

    \I__1945\ : Span4Mux_h
    port map (
            O => \N__9071\,
            I => \N__9065\
        );

    \I__1944\ : Span12Mux_v
    port map (
            O => \N__9068\,
            I => \N__9062\
        );

    \I__1943\ : Span4Mux_h
    port map (
            O => \N__9065\,
            I => \N__9059\
        );

    \I__1942\ : Odrv12
    port map (
            O => \N__9062\,
            I => \SIZ_c_1\
        );

    \I__1941\ : Odrv4
    port map (
            O => \N__9059\,
            I => \SIZ_c_1\
        );

    \I__1940\ : CascadeMux
    port map (
            O => \N__9054\,
            I => \N__9048\
        );

    \I__1939\ : CascadeMux
    port map (
            O => \N__9053\,
            I => \N__9045\
        );

    \I__1938\ : InMux
    port map (
            O => \N__9052\,
            I => \N__9039\
        );

    \I__1937\ : InMux
    port map (
            O => \N__9051\,
            I => \N__9036\
        );

    \I__1936\ : InMux
    port map (
            O => \N__9048\,
            I => \N__9029\
        );

    \I__1935\ : InMux
    port map (
            O => \N__9045\,
            I => \N__9029\
        );

    \I__1934\ : InMux
    port map (
            O => \N__9044\,
            I => \N__9029\
        );

    \I__1933\ : InMux
    port map (
            O => \N__9043\,
            I => \N__9024\
        );

    \I__1932\ : InMux
    port map (
            O => \N__9042\,
            I => \N__9024\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__9039\,
            I => \N__9021\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__9036\,
            I => \N__9015\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__9029\,
            I => \N__9015\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__9024\,
            I => \N__9012\
        );

    \I__1927\ : Span4Mux_v
    port map (
            O => \N__9021\,
            I => \N__9009\
        );

    \I__1926\ : InMux
    port map (
            O => \N__9020\,
            I => \N__9006\
        );

    \I__1925\ : Span12Mux_v
    port map (
            O => \N__9015\,
            I => \N__9001\
        );

    \I__1924\ : Span12Mux_s7_v
    port map (
            O => \N__9012\,
            I => \N__9001\
        );

    \I__1923\ : Span4Mux_h
    port map (
            O => \N__9009\,
            I => \N__8998\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__9006\,
            I => \N__8995\
        );

    \I__1921\ : Span12Mux_h
    port map (
            O => \N__9001\,
            I => \N__8992\
        );

    \I__1920\ : Sp12to4
    port map (
            O => \N__8998\,
            I => \N__8987\
        );

    \I__1919\ : Span12Mux_h
    port map (
            O => \N__8995\,
            I => \N__8987\
        );

    \I__1918\ : Odrv12
    port map (
            O => \N__8992\,
            I => \A_c_1\
        );

    \I__1917\ : Odrv12
    port map (
            O => \N__8987\,
            I => \A_c_1\
        );

    \I__1916\ : InMux
    port map (
            O => \N__8982\,
            I => \N__8977\
        );

    \I__1915\ : InMux
    port map (
            O => \N__8981\,
            I => \N__8970\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__8980\,
            I => \N__8966\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__8977\,
            I => \N__8963\
        );

    \I__1912\ : InMux
    port map (
            O => \N__8976\,
            I => \N__8960\
        );

    \I__1911\ : CascadeMux
    port map (
            O => \N__8975\,
            I => \N__8957\
        );

    \I__1910\ : CascadeMux
    port map (
            O => \N__8974\,
            I => \N__8954\
        );

    \I__1909\ : CascadeMux
    port map (
            O => \N__8973\,
            I => \N__8951\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8970\,
            I => \N__8948\
        );

    \I__1907\ : InMux
    port map (
            O => \N__8969\,
            I => \N__8945\
        );

    \I__1906\ : InMux
    port map (
            O => \N__8966\,
            I => \N__8941\
        );

    \I__1905\ : Span4Mux_v
    port map (
            O => \N__8963\,
            I => \N__8938\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__8960\,
            I => \N__8935\
        );

    \I__1903\ : InMux
    port map (
            O => \N__8957\,
            I => \N__8930\
        );

    \I__1902\ : InMux
    port map (
            O => \N__8954\,
            I => \N__8930\
        );

    \I__1901\ : InMux
    port map (
            O => \N__8951\,
            I => \N__8927\
        );

    \I__1900\ : Span4Mux_v
    port map (
            O => \N__8948\,
            I => \N__8922\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__8945\,
            I => \N__8922\
        );

    \I__1898\ : InMux
    port map (
            O => \N__8944\,
            I => \N__8919\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__8941\,
            I => \N__8916\
        );

    \I__1896\ : Span4Mux_v
    port map (
            O => \N__8938\,
            I => \N__8913\
        );

    \I__1895\ : Span4Mux_v
    port map (
            O => \N__8935\,
            I => \N__8910\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__8930\,
            I => \N__8905\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__8927\,
            I => \N__8905\
        );

    \I__1892\ : Span4Mux_h
    port map (
            O => \N__8922\,
            I => \N__8900\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__8919\,
            I => \N__8900\
        );

    \I__1890\ : Span12Mux_v
    port map (
            O => \N__8916\,
            I => \N__8891\
        );

    \I__1889\ : Sp12to4
    port map (
            O => \N__8913\,
            I => \N__8891\
        );

    \I__1888\ : Sp12to4
    port map (
            O => \N__8910\,
            I => \N__8891\
        );

    \I__1887\ : Span12Mux_s10_v
    port map (
            O => \N__8905\,
            I => \N__8891\
        );

    \I__1886\ : Span4Mux_v
    port map (
            O => \N__8900\,
            I => \N__8888\
        );

    \I__1885\ : Span12Mux_h
    port map (
            O => \N__8891\,
            I => \N__8885\
        );

    \I__1884\ : Sp12to4
    port map (
            O => \N__8888\,
            I => \N__8882\
        );

    \I__1883\ : Odrv12
    port map (
            O => \N__8885\,
            I => \A_c_0\
        );

    \I__1882\ : Odrv12
    port map (
            O => \N__8882\,
            I => \A_c_0\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__8877\,
            I => \N__8873\
        );

    \I__1880\ : InMux
    port map (
            O => \N__8876\,
            I => \N__8868\
        );

    \I__1879\ : InMux
    port map (
            O => \N__8873\,
            I => \N__8865\
        );

    \I__1878\ : InMux
    port map (
            O => \N__8872\,
            I => \N__8862\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__8871\,
            I => \N__8857\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__8868\,
            I => \N__8854\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__8865\,
            I => \N__8850\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__8862\,
            I => \N__8847\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8861\,
            I => \N__8842\
        );

    \I__1872\ : InMux
    port map (
            O => \N__8860\,
            I => \N__8842\
        );

    \I__1871\ : InMux
    port map (
            O => \N__8857\,
            I => \N__8839\
        );

    \I__1870\ : Span4Mux_v
    port map (
            O => \N__8854\,
            I => \N__8836\
        );

    \I__1869\ : InMux
    port map (
            O => \N__8853\,
            I => \N__8833\
        );

    \I__1868\ : Span4Mux_v
    port map (
            O => \N__8850\,
            I => \N__8830\
        );

    \I__1867\ : Span4Mux_v
    port map (
            O => \N__8847\,
            I => \N__8823\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__8842\,
            I => \N__8823\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__8839\,
            I => \N__8823\
        );

    \I__1864\ : Sp12to4
    port map (
            O => \N__8836\,
            I => \N__8818\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__8833\,
            I => \N__8818\
        );

    \I__1862\ : Span4Mux_v
    port map (
            O => \N__8830\,
            I => \N__8813\
        );

    \I__1861\ : Span4Mux_h
    port map (
            O => \N__8823\,
            I => \N__8813\
        );

    \I__1860\ : Span12Mux_h
    port map (
            O => \N__8818\,
            I => \N__8810\
        );

    \I__1859\ : Span4Mux_v
    port map (
            O => \N__8813\,
            I => \N__8807\
        );

    \I__1858\ : Span12Mux_v
    port map (
            O => \N__8810\,
            I => \N__8804\
        );

    \I__1857\ : Sp12to4
    port map (
            O => \N__8807\,
            I => \N__8801\
        );

    \I__1856\ : Odrv12
    port map (
            O => \N__8804\,
            I => \SIZ_c_0\
        );

    \I__1855\ : Odrv12
    port map (
            O => \N__8801\,
            I => \SIZ_c_0\
        );

    \I__1854\ : IoInMux
    port map (
            O => \N__8796\,
            I => \N__8793\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__8793\,
            I => \N__8790\
        );

    \I__1852\ : Span4Mux_s3_v
    port map (
            O => \N__8790\,
            I => \N__8787\
        );

    \I__1851\ : Span4Mux_h
    port map (
            O => \N__8787\,
            I => \N__8784\
        );

    \I__1850\ : Odrv4
    port map (
            O => \N__8784\,
            I => \N_344_i\
        );

    \I__1849\ : InMux
    port map (
            O => \N__8781\,
            I => \N__8778\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__8778\,
            I => \N__8774\
        );

    \I__1847\ : InMux
    port map (
            O => \N__8777\,
            I => \N__8771\
        );

    \I__1846\ : Span4Mux_v
    port map (
            O => \N__8774\,
            I => \N__8764\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__8771\,
            I => \N__8764\
        );

    \I__1844\ : InMux
    port map (
            O => \N__8770\,
            I => \N__8760\
        );

    \I__1843\ : CascadeMux
    port map (
            O => \N__8769\,
            I => \N__8757\
        );

    \I__1842\ : Span4Mux_h
    port map (
            O => \N__8764\,
            I => \N__8754\
        );

    \I__1841\ : InMux
    port map (
            O => \N__8763\,
            I => \N__8751\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__8760\,
            I => \N__8748\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8757\,
            I => \N__8745\
        );

    \I__1838\ : Odrv4
    port map (
            O => \N__8754\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__8751\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1836\ : Odrv12
    port map (
            O => \N__8748\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__8745\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1834\ : IoInMux
    port map (
            O => \N__8736\,
            I => \N__8733\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__8733\,
            I => \N__8730\
        );

    \I__1832\ : Span4Mux_s3_v
    port map (
            O => \N__8730\,
            I => \N__8727\
        );

    \I__1831\ : Sp12to4
    port map (
            O => \N__8727\,
            I => \N__8724\
        );

    \I__1830\ : Span12Mux_h
    port map (
            O => \N__8724\,
            I => \N__8721\
        );

    \I__1829\ : Odrv12
    port map (
            O => \N__8721\,
            I => \CRCSn_c\
        );

    \I__1828\ : InMux
    port map (
            O => \N__8718\,
            I => \N__8715\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8715\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__1826\ : IoInMux
    port map (
            O => \N__8712\,
            I => \N__8709\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__8709\,
            I => \N__8706\
        );

    \I__1824\ : Span4Mux_s3_v
    port map (
            O => \N__8706\,
            I => \N__8703\
        );

    \I__1823\ : Span4Mux_v
    port map (
            O => \N__8703\,
            I => \N__8700\
        );

    \I__1822\ : Span4Mux_h
    port map (
            O => \N__8700\,
            I => \N__8697\
        );

    \I__1821\ : Odrv4
    port map (
            O => \N__8697\,
            I => \CMA_c_0\
        );

    \I__1820\ : InMux
    port map (
            O => \N__8694\,
            I => \N__8691\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__8691\,
            I => \N__8688\
        );

    \I__1818\ : Odrv12
    port map (
            O => \N__8688\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8685\,
            I => \N__8682\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__8682\,
            I => \N__8679\
        );

    \I__1815\ : Span4Mux_v
    port map (
            O => \N__8679\,
            I => \N__8676\
        );

    \I__1814\ : Sp12to4
    port map (
            O => \N__8676\,
            I => \N__8673\
        );

    \I__1813\ : Span12Mux_h
    port map (
            O => \N__8673\,
            I => \N__8670\
        );

    \I__1812\ : Odrv12
    port map (
            O => \N__8670\,
            I => \A_c_12\
        );

    \I__1811\ : CascadeMux
    port map (
            O => \N__8667\,
            I => \N__8660\
        );

    \I__1810\ : CascadeMux
    port map (
            O => \N__8666\,
            I => \N__8656\
        );

    \I__1809\ : CascadeMux
    port map (
            O => \N__8665\,
            I => \N__8648\
        );

    \I__1808\ : CascadeMux
    port map (
            O => \N__8664\,
            I => \N__8645\
        );

    \I__1807\ : InMux
    port map (
            O => \N__8663\,
            I => \N__8638\
        );

    \I__1806\ : InMux
    port map (
            O => \N__8660\,
            I => \N__8635\
        );

    \I__1805\ : CascadeMux
    port map (
            O => \N__8659\,
            I => \N__8632\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8656\,
            I => \N__8625\
        );

    \I__1803\ : InMux
    port map (
            O => \N__8655\,
            I => \N__8620\
        );

    \I__1802\ : InMux
    port map (
            O => \N__8654\,
            I => \N__8620\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8653\,
            I => \N__8611\
        );

    \I__1800\ : InMux
    port map (
            O => \N__8652\,
            I => \N__8611\
        );

    \I__1799\ : InMux
    port map (
            O => \N__8651\,
            I => \N__8603\
        );

    \I__1798\ : InMux
    port map (
            O => \N__8648\,
            I => \N__8603\
        );

    \I__1797\ : InMux
    port map (
            O => \N__8645\,
            I => \N__8600\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8644\,
            I => \N__8591\
        );

    \I__1795\ : InMux
    port map (
            O => \N__8643\,
            I => \N__8591\
        );

    \I__1794\ : InMux
    port map (
            O => \N__8642\,
            I => \N__8591\
        );

    \I__1793\ : InMux
    port map (
            O => \N__8641\,
            I => \N__8591\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__8638\,
            I => \N__8586\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__8635\,
            I => \N__8586\
        );

    \I__1790\ : InMux
    port map (
            O => \N__8632\,
            I => \N__8583\
        );

    \I__1789\ : InMux
    port map (
            O => \N__8631\,
            I => \N__8574\
        );

    \I__1788\ : InMux
    port map (
            O => \N__8630\,
            I => \N__8574\
        );

    \I__1787\ : InMux
    port map (
            O => \N__8629\,
            I => \N__8574\
        );

    \I__1786\ : InMux
    port map (
            O => \N__8628\,
            I => \N__8574\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__8625\,
            I => \N__8569\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__8620\,
            I => \N__8569\
        );

    \I__1783\ : InMux
    port map (
            O => \N__8619\,
            I => \N__8566\
        );

    \I__1782\ : InMux
    port map (
            O => \N__8618\,
            I => \N__8559\
        );

    \I__1781\ : InMux
    port map (
            O => \N__8617\,
            I => \N__8559\
        );

    \I__1780\ : InMux
    port map (
            O => \N__8616\,
            I => \N__8559\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__8611\,
            I => \N__8556\
        );

    \I__1778\ : InMux
    port map (
            O => \N__8610\,
            I => \N__8549\
        );

    \I__1777\ : InMux
    port map (
            O => \N__8609\,
            I => \N__8549\
        );

    \I__1776\ : InMux
    port map (
            O => \N__8608\,
            I => \N__8549\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__8603\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__8600\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__8591\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1772\ : Odrv4
    port map (
            O => \N__8586\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__8583\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__8574\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1769\ : Odrv4
    port map (
            O => \N__8569\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__8566\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__8559\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1766\ : Odrv4
    port map (
            O => \N__8556\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__8549\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1764\ : CascadeMux
    port map (
            O => \N__8526\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\
        );

    \I__1763\ : CascadeMux
    port map (
            O => \N__8523\,
            I => \U712_BYTE_ENABLE.N_454_cascade_\
        );

    \I__1762\ : IoInMux
    port map (
            O => \N__8520\,
            I => \N__8517\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__8517\,
            I => \N__8514\
        );

    \I__1760\ : Span12Mux_s6_h
    port map (
            O => \N__8514\,
            I => \N__8511\
        );

    \I__1759\ : Span12Mux_v
    port map (
            O => \N__8511\,
            I => \N__8508\
        );

    \I__1758\ : Odrv12
    port map (
            O => \N__8508\,
            I => \N_215_i\
        );

    \I__1757\ : IoInMux
    port map (
            O => \N__8505\,
            I => \N__8502\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__8502\,
            I => \N__8499\
        );

    \I__1755\ : Span4Mux_s3_h
    port map (
            O => \N__8499\,
            I => \N__8496\
        );

    \I__1754\ : Sp12to4
    port map (
            O => \N__8496\,
            I => \N__8493\
        );

    \I__1753\ : Span12Mux_v
    port map (
            O => \N__8493\,
            I => \N__8490\
        );

    \I__1752\ : Span12Mux_h
    port map (
            O => \N__8490\,
            I => \N__8487\
        );

    \I__1751\ : Odrv12
    port map (
            O => \N__8487\,
            I => \N_213_i\
        );

    \I__1750\ : IoInMux
    port map (
            O => \N__8484\,
            I => \N__8481\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__8481\,
            I => \N__8478\
        );

    \I__1748\ : Span4Mux_s2_v
    port map (
            O => \N__8478\,
            I => \N__8471\
        );

    \I__1747\ : InMux
    port map (
            O => \N__8477\,
            I => \N__8468\
        );

    \I__1746\ : InMux
    port map (
            O => \N__8476\,
            I => \N__8465\
        );

    \I__1745\ : InMux
    port map (
            O => \N__8475\,
            I => \N__8460\
        );

    \I__1744\ : InMux
    port map (
            O => \N__8474\,
            I => \N__8460\
        );

    \I__1743\ : Span4Mux_h
    port map (
            O => \N__8471\,
            I => \N__8457\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__8468\,
            I => \N__8450\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__8465\,
            I => \N__8450\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__8460\,
            I => \N__8450\
        );

    \I__1739\ : Sp12to4
    port map (
            O => \N__8457\,
            I => \N__8446\
        );

    \I__1738\ : Span4Mux_v
    port map (
            O => \N__8450\,
            I => \N__8443\
        );

    \I__1737\ : InMux
    port map (
            O => \N__8449\,
            I => \N__8440\
        );

    \I__1736\ : Odrv12
    port map (
            O => \N__8446\,
            I => \DBENn_c\
        );

    \I__1735\ : Odrv4
    port map (
            O => \N__8443\,
            I => \DBENn_c\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__8440\,
            I => \DBENn_c\
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__8433\,
            I => \U712_BYTE_ENABLE.N_450_cascade_\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__8430\,
            I => \N__8426\
        );

    \I__1731\ : InMux
    port map (
            O => \N__8429\,
            I => \N__8421\
        );

    \I__1730\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8418\
        );

    \I__1729\ : InMux
    port map (
            O => \N__8425\,
            I => \N__8413\
        );

    \I__1728\ : InMux
    port map (
            O => \N__8424\,
            I => \N__8413\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__8421\,
            I => \N__8405\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__8418\,
            I => \N__8405\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__8413\,
            I => \N__8405\
        );

    \I__1724\ : InMux
    port map (
            O => \N__8412\,
            I => \N__8401\
        );

    \I__1723\ : Span4Mux_v
    port map (
            O => \N__8405\,
            I => \N__8396\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8404\,
            I => \N__8393\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__8401\,
            I => \N__8390\
        );

    \I__1720\ : InMux
    port map (
            O => \N__8400\,
            I => \N__8385\
        );

    \I__1719\ : InMux
    port map (
            O => \N__8399\,
            I => \N__8385\
        );

    \I__1718\ : Odrv4
    port map (
            O => \N__8396\,
            I => \DMA_CYCLEm\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__8393\,
            I => \DMA_CYCLEm\
        );

    \I__1716\ : Odrv4
    port map (
            O => \N__8390\,
            I => \DMA_CYCLEm\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__8385\,
            I => \DMA_CYCLEm\
        );

    \I__1714\ : IoInMux
    port map (
            O => \N__8376\,
            I => \N__8373\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__8373\,
            I => \N__8370\
        );

    \I__1712\ : Span4Mux_s2_h
    port map (
            O => \N__8370\,
            I => \N__8367\
        );

    \I__1711\ : Span4Mux_v
    port map (
            O => \N__8367\,
            I => \N__8364\
        );

    \I__1710\ : Sp12to4
    port map (
            O => \N__8364\,
            I => \N__8361\
        );

    \I__1709\ : Span12Mux_h
    port map (
            O => \N__8361\,
            I => \N__8358\
        );

    \I__1708\ : Odrv12
    port map (
            O => \N__8358\,
            I => \N_211_i\
        );

    \I__1707\ : InMux
    port map (
            O => \N__8355\,
            I => \N__8352\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__8352\,
            I => \U712_BYTE_ENABLE.N_456\
        );

    \I__1705\ : CascadeMux
    port map (
            O => \N__8349\,
            I => \N__8343\
        );

    \I__1704\ : InMux
    port map (
            O => \N__8348\,
            I => \N__8340\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8347\,
            I => \N__8333\
        );

    \I__1702\ : InMux
    port map (
            O => \N__8346\,
            I => \N__8333\
        );

    \I__1701\ : InMux
    port map (
            O => \N__8343\,
            I => \N__8333\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8340\,
            I => \N__8330\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__8333\,
            I => \N__8327\
        );

    \I__1698\ : Odrv4
    port map (
            O => \N__8330\,
            I => \U712_BYTE_ENABLE.N_315_i\
        );

    \I__1697\ : Odrv4
    port map (
            O => \N__8327\,
            I => \U712_BYTE_ENABLE.N_315_i\
        );

    \I__1696\ : InMux
    port map (
            O => \N__8322\,
            I => \N__8319\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8319\,
            I => \U712_BYTE_ENABLE.N_452\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8316\,
            I => \N__8313\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__8313\,
            I => \N__8310\
        );

    \I__1692\ : Span4Mux_h
    port map (
            O => \N__8310\,
            I => \N__8307\
        );

    \I__1691\ : Sp12to4
    port map (
            O => \N__8307\,
            I => \N__8304\
        );

    \I__1690\ : Span12Mux_v
    port map (
            O => \N__8304\,
            I => \N__8301\
        );

    \I__1689\ : Span12Mux_h
    port map (
            O => \N__8301\,
            I => \N__8298\
        );

    \I__1688\ : Odrv12
    port map (
            O => \N__8298\,
            I => \A_c_14\
        );

    \I__1687\ : InMux
    port map (
            O => \N__8295\,
            I => \N__8292\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__8292\,
            I => \U712_CHIP_RAM.N_368\
        );

    \I__1685\ : CascadeMux
    port map (
            O => \N__8289\,
            I => \U712_CHIP_RAM.N_330_cascade_\
        );

    \I__1684\ : InMux
    port map (
            O => \N__8286\,
            I => \N__8283\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__8283\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__1682\ : InMux
    port map (
            O => \N__8280\,
            I => \N__8277\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__8277\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__1680\ : InMux
    port map (
            O => \N__8274\,
            I => \N__8271\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__8271\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8\
        );

    \I__1678\ : InMux
    port map (
            O => \N__8268\,
            I => \N__8265\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__8265\,
            I => \N__8262\
        );

    \I__1676\ : Span12Mux_v
    port map (
            O => \N__8262\,
            I => \N__8259\
        );

    \I__1675\ : Span12Mux_h
    port map (
            O => \N__8259\,
            I => \N__8256\
        );

    \I__1674\ : Odrv12
    port map (
            O => \N__8256\,
            I => \A_c_13\
        );

    \I__1673\ : InMux
    port map (
            O => \N__8253\,
            I => \N__8250\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__8250\,
            I => \N__8247\
        );

    \I__1671\ : Span4Mux_h
    port map (
            O => \N__8247\,
            I => \N__8244\
        );

    \I__1670\ : Span4Mux_h
    port map (
            O => \N__8244\,
            I => \N__8241\
        );

    \I__1669\ : Odrv4
    port map (
            O => \N__8241\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\
        );

    \I__1668\ : CascadeMux
    port map (
            O => \N__8238\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\
        );

    \I__1667\ : IoInMux
    port map (
            O => \N__8235\,
            I => \N__8232\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__8232\,
            I => \N__8229\
        );

    \I__1665\ : Span12Mux_s9_v
    port map (
            O => \N__8229\,
            I => \N__8226\
        );

    \I__1664\ : Span12Mux_h
    port map (
            O => \N__8226\,
            I => \N__8223\
        );

    \I__1663\ : Odrv12
    port map (
            O => \N__8223\,
            I => \CASn_c\
        );

    \I__1662\ : InMux
    port map (
            O => \N__8220\,
            I => \N__8217\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__8217\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__1660\ : InMux
    port map (
            O => \N__8214\,
            I => \N__8211\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__8211\,
            I => \N__8208\
        );

    \I__1658\ : Span4Mux_h
    port map (
            O => \N__8208\,
            I => \N__8205\
        );

    \I__1657\ : Odrv4
    port map (
            O => \N__8205\,
            I => \U712_CHIP_RAM.N_374\
        );

    \I__1656\ : IoInMux
    port map (
            O => \N__8202\,
            I => \N__8199\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__8199\,
            I => \N__8196\
        );

    \I__1654\ : Span4Mux_s3_h
    port map (
            O => \N__8196\,
            I => \N__8193\
        );

    \I__1653\ : Span4Mux_v
    port map (
            O => \N__8193\,
            I => \N__8190\
        );

    \I__1652\ : Span4Mux_h
    port map (
            O => \N__8190\,
            I => \N__8187\
        );

    \I__1651\ : Span4Mux_h
    port map (
            O => \N__8187\,
            I => \N__8184\
        );

    \I__1650\ : Span4Mux_h
    port map (
            O => \N__8184\,
            I => \N__8181\
        );

    \I__1649\ : Odrv4
    port map (
            O => \N__8181\,
            I => \CMA_c_5\
        );

    \I__1648\ : IoInMux
    port map (
            O => \N__8178\,
            I => \N__8175\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__8175\,
            I => \N__8172\
        );

    \I__1646\ : Span4Mux_s3_v
    port map (
            O => \N__8172\,
            I => \N__8169\
        );

    \I__1645\ : Sp12to4
    port map (
            O => \N__8169\,
            I => \N__8166\
        );

    \I__1644\ : Span12Mux_h
    port map (
            O => \N__8166\,
            I => \N__8163\
        );

    \I__1643\ : Odrv12
    port map (
            O => \N__8163\,
            I => \CMA_c_10\
        );

    \I__1642\ : IoInMux
    port map (
            O => \N__8160\,
            I => \N__8157\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__8157\,
            I => \N__8154\
        );

    \I__1640\ : Span12Mux_s5_v
    port map (
            O => \N__8154\,
            I => \N__8151\
        );

    \I__1639\ : Odrv12
    port map (
            O => \N__8151\,
            I => \CMA_c_1\
        );

    \I__1638\ : CascadeMux
    port map (
            O => \N__8148\,
            I => \N__8145\
        );

    \I__1637\ : InMux
    port map (
            O => \N__8145\,
            I => \N__8142\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__8142\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\
        );

    \I__1635\ : CascadeMux
    port map (
            O => \N__8139\,
            I => \N__8136\
        );

    \I__1634\ : InMux
    port map (
            O => \N__8136\,
            I => \N__8133\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__8133\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\
        );

    \I__1632\ : SRMux
    port map (
            O => \N__8130\,
            I => \N__8126\
        );

    \I__1631\ : InMux
    port map (
            O => \N__8129\,
            I => \N__8123\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__8126\,
            I => \N__8120\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__8123\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1628\ : Odrv12
    port map (
            O => \N__8120\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__8115\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_cascade_\
        );

    \I__1626\ : InMux
    port map (
            O => \N__8112\,
            I => \N__8109\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__8109\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__1624\ : InMux
    port map (
            O => \N__8106\,
            I => \N__8103\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__8103\,
            I => \N__8100\
        );

    \I__1622\ : Odrv12
    port map (
            O => \N__8100\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\
        );

    \I__1621\ : InMux
    port map (
            O => \N__8097\,
            I => \N__8091\
        );

    \I__1620\ : InMux
    port map (
            O => \N__8096\,
            I => \N__8091\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__8091\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\
        );

    \I__1618\ : IoInMux
    port map (
            O => \N__8088\,
            I => \N__8085\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__8085\,
            I => \N__8082\
        );

    \I__1616\ : IoSpan4Mux
    port map (
            O => \N__8082\,
            I => \N__8079\
        );

    \I__1615\ : Span4Mux_s2_v
    port map (
            O => \N__8079\,
            I => \N__8076\
        );

    \I__1614\ : Sp12to4
    port map (
            O => \N__8076\,
            I => \N__8073\
        );

    \I__1613\ : Odrv12
    port map (
            O => \N__8073\,
            I => \N_217_i\
        );

    \I__1612\ : InMux
    port map (
            O => \N__8070\,
            I => \N__8067\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__8067\,
            I => \N__8064\
        );

    \I__1610\ : Span4Mux_h
    port map (
            O => \N__8064\,
            I => \N__8060\
        );

    \I__1609\ : InMux
    port map (
            O => \N__8063\,
            I => \N__8057\
        );

    \I__1608\ : Span4Mux_v
    port map (
            O => \N__8060\,
            I => \N__8052\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__8057\,
            I => \N__8052\
        );

    \I__1606\ : Span4Mux_v
    port map (
            O => \N__8052\,
            I => \N__8047\
        );

    \I__1605\ : InMux
    port map (
            O => \N__8051\,
            I => \N__8042\
        );

    \I__1604\ : InMux
    port map (
            O => \N__8050\,
            I => \N__8042\
        );

    \I__1603\ : Odrv4
    port map (
            O => \N__8047\,
            I => \REG_CYCLEm\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__8042\,
            I => \REG_CYCLEm\
        );

    \I__1601\ : IoInMux
    port map (
            O => \N__8037\,
            I => \N__8034\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__8034\,
            I => \N__8031\
        );

    \I__1599\ : IoSpan4Mux
    port map (
            O => \N__8031\,
            I => \N__8028\
        );

    \I__1598\ : Span4Mux_s2_v
    port map (
            O => \N__8028\,
            I => \N__8025\
        );

    \I__1597\ : Span4Mux_v
    port map (
            O => \N__8025\,
            I => \N__8022\
        );

    \I__1596\ : Sp12to4
    port map (
            O => \N__8022\,
            I => \N__8019\
        );

    \I__1595\ : Span12Mux_h
    port map (
            O => \N__8019\,
            I => \N__8016\
        );

    \I__1594\ : Odrv12
    port map (
            O => \N__8016\,
            I => \N_182_i\
        );

    \I__1593\ : InMux
    port map (
            O => \N__8013\,
            I => \N__8010\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__8010\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1591\ : InMux
    port map (
            O => \N__8007\,
            I => \N__8004\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__8004\,
            I => \U712_REG_SM.N_434\
        );

    \I__1589\ : IoInMux
    port map (
            O => \N__8001\,
            I => \N__7998\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__7998\,
            I => \N__7995\
        );

    \I__1587\ : Span12Mux_s7_v
    port map (
            O => \N__7995\,
            I => \N__7992\
        );

    \I__1586\ : Odrv12
    port map (
            O => \N__7992\,
            I => \N_198_i\
        );

    \I__1585\ : IoInMux
    port map (
            O => \N__7989\,
            I => \N__7986\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__7986\,
            I => \N__7983\
        );

    \I__1583\ : IoSpan4Mux
    port map (
            O => \N__7983\,
            I => \N__7980\
        );

    \I__1582\ : IoSpan4Mux
    port map (
            O => \N__7980\,
            I => \N__7977\
        );

    \I__1581\ : Span4Mux_s2_v
    port map (
            O => \N__7977\,
            I => \N__7974\
        );

    \I__1580\ : Span4Mux_v
    port map (
            O => \N__7974\,
            I => \N__7971\
        );

    \I__1579\ : Odrv4
    port map (
            O => \N__7971\,
            I => \N_343_i\
        );

    \I__1578\ : InMux
    port map (
            O => \N__7968\,
            I => \N__7965\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__7965\,
            I => \N__7962\
        );

    \I__1576\ : Odrv4
    port map (
            O => \N__7962\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__7959\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_\
        );

    \I__1574\ : IoInMux
    port map (
            O => \N__7956\,
            I => \N__7953\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__7953\,
            I => \N__7950\
        );

    \I__1572\ : Span12Mux_s5_v
    port map (
            O => \N__7950\,
            I => \N__7947\
        );

    \I__1571\ : Odrv12
    port map (
            O => \N__7947\,
            I => \CMA_c_2\
        );

    \I__1570\ : InMux
    port map (
            O => \N__7944\,
            I => \N__7941\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__7941\,
            I => \N__7938\
        );

    \I__1568\ : Span4Mux_v
    port map (
            O => \N__7938\,
            I => \N__7935\
        );

    \I__1567\ : Span4Mux_v
    port map (
            O => \N__7935\,
            I => \N__7932\
        );

    \I__1566\ : Sp12to4
    port map (
            O => \N__7932\,
            I => \N__7929\
        );

    \I__1565\ : Span12Mux_h
    port map (
            O => \N__7929\,
            I => \N__7926\
        );

    \I__1564\ : Odrv12
    port map (
            O => \N__7926\,
            I => \A_c_16\
        );

    \I__1563\ : InMux
    port map (
            O => \N__7923\,
            I => \N__7920\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__7920\,
            I => \N__7917\
        );

    \I__1561\ : Odrv12
    port map (
            O => \N__7917\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\
        );

    \I__1560\ : CascadeMux
    port map (
            O => \N__7914\,
            I => \N__7911\
        );

    \I__1559\ : InMux
    port map (
            O => \N__7911\,
            I => \N__7908\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__7908\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_i_i_0\
        );

    \I__1557\ : InMux
    port map (
            O => \N__7905\,
            I => \N__7902\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__7902\,
            I => \U712_CHIP_RAM.N_408\
        );

    \I__1555\ : InMux
    port map (
            O => \N__7899\,
            I => \N__7894\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7898\,
            I => \N__7889\
        );

    \I__1553\ : InMux
    port map (
            O => \N__7897\,
            I => \N__7889\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__7894\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__7889\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7884\,
            I => \N__7881\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__7881\,
            I => \U712_CHIP_RAM.N_151\
        );

    \I__1548\ : IoInMux
    port map (
            O => \N__7878\,
            I => \N__7875\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__7875\,
            I => \N__7872\
        );

    \I__1546\ : Span4Mux_s0_v
    port map (
            O => \N__7872\,
            I => \N__7869\
        );

    \I__1545\ : Span4Mux_v
    port map (
            O => \N__7869\,
            I => \N__7865\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7868\,
            I => \N__7862\
        );

    \I__1543\ : Span4Mux_v
    port map (
            O => \N__7865\,
            I => \N__7859\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__7862\,
            I => \N__7856\
        );

    \I__1541\ : Sp12to4
    port map (
            O => \N__7859\,
            I => \N__7853\
        );

    \I__1540\ : Span4Mux_v
    port map (
            O => \N__7856\,
            I => \N__7850\
        );

    \I__1539\ : Span12Mux_h
    port map (
            O => \N__7853\,
            I => \N__7847\
        );

    \I__1538\ : Sp12to4
    port map (
            O => \N__7850\,
            I => \N__7844\
        );

    \I__1537\ : Span12Mux_v
    port map (
            O => \N__7847\,
            I => \N__7839\
        );

    \I__1536\ : Span12Mux_h
    port map (
            O => \N__7844\,
            I => \N__7839\
        );

    \I__1535\ : Odrv12
    port map (
            O => \N__7839\,
            I => \A_c_10\
        );

    \I__1534\ : InMux
    port map (
            O => \N__7836\,
            I => \N__7833\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__7833\,
            I => \N__7830\
        );

    \I__1532\ : Span4Mux_v
    port map (
            O => \N__7830\,
            I => \N__7827\
        );

    \I__1531\ : Odrv4
    port map (
            O => \N__7827\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\
        );

    \I__1530\ : CascadeMux
    port map (
            O => \N__7824\,
            I => \N__7821\
        );

    \I__1529\ : InMux
    port map (
            O => \N__7821\,
            I => \N__7818\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__7818\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\
        );

    \I__1527\ : InMux
    port map (
            O => \N__7815\,
            I => \N__7812\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__7812\,
            I => \N__7809\
        );

    \I__1525\ : Sp12to4
    port map (
            O => \N__7809\,
            I => \N__7806\
        );

    \I__1524\ : Span12Mux_v
    port map (
            O => \N__7806\,
            I => \N__7803\
        );

    \I__1523\ : Span12Mux_h
    port map (
            O => \N__7803\,
            I => \N__7800\
        );

    \I__1522\ : Odrv12
    port map (
            O => \N__7800\,
            I => \A_c_17\
        );

    \I__1521\ : InMux
    port map (
            O => \N__7797\,
            I => \N__7793\
        );

    \I__1520\ : InMux
    port map (
            O => \N__7796\,
            I => \N__7790\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__7793\,
            I => \N__7787\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__7790\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__1517\ : Odrv4
    port map (
            O => \N__7787\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__1516\ : InMux
    port map (
            O => \N__7782\,
            I => \N__7779\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__7779\,
            I => \N__7776\
        );

    \I__1514\ : Odrv4
    port map (
            O => \N__7776\,
            I => \U712_CHIP_RAM.N_471\
        );

    \I__1513\ : InMux
    port map (
            O => \N__7773\,
            I => \N__7770\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__7770\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_5\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7767\,
            I => \N__7762\
        );

    \I__1510\ : InMux
    port map (
            O => \N__7766\,
            I => \N__7759\
        );

    \I__1509\ : CascadeMux
    port map (
            O => \N__7765\,
            I => \N__7756\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7762\,
            I => \N__7752\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__7759\,
            I => \N__7749\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7756\,
            I => \N__7746\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7755\,
            I => \N__7743\
        );

    \I__1504\ : Span4Mux_v
    port map (
            O => \N__7752\,
            I => \N__7734\
        );

    \I__1503\ : Span4Mux_h
    port map (
            O => \N__7749\,
            I => \N__7734\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__7746\,
            I => \N__7734\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__7743\,
            I => \N__7734\
        );

    \I__1500\ : Span4Mux_v
    port map (
            O => \N__7734\,
            I => \N__7731\
        );

    \I__1499\ : Span4Mux_h
    port map (
            O => \N__7731\,
            I => \N__7728\
        );

    \I__1498\ : Span4Mux_v
    port map (
            O => \N__7728\,
            I => \N__7725\
        );

    \I__1497\ : Span4Mux_v
    port map (
            O => \N__7725\,
            I => \N__7722\
        );

    \I__1496\ : Odrv4
    port map (
            O => \N__7722\,
            I => \CLK40_PLL_i\
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__7719\,
            I => \N__7716\
        );

    \I__1494\ : InMux
    port map (
            O => \N__7716\,
            I => \N__7711\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7715\,
            I => \N__7708\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7714\,
            I => \N__7704\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__7711\,
            I => \N__7699\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__7708\,
            I => \N__7699\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7707\,
            I => \N__7696\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__7704\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1487\ : Odrv4
    port map (
            O => \N__7699\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__7696\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1485\ : InMux
    port map (
            O => \N__7689\,
            I => \N__7683\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7688\,
            I => \N__7683\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7683\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7680\,
            I => \N__7675\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7679\,
            I => \N__7670\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7678\,
            I => \N__7670\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7675\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__7670\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7665\,
            I => \N__7661\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7664\,
            I => \N__7658\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__7661\,
            I => \N__7655\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7658\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\
        );

    \I__1473\ : Odrv4
    port map (
            O => \N__7655\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7650\,
            I => \N__7646\
        );

    \I__1471\ : InMux
    port map (
            O => \N__7649\,
            I => \N__7643\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__7646\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_1\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__7643\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_1\
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__7638\,
            I => \N__7635\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7635\,
            I => \N__7631\
        );

    \I__1466\ : InMux
    port map (
            O => \N__7634\,
            I => \N__7628\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__7631\,
            I => \N__7625\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__7628\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\
        );

    \I__1463\ : Odrv4
    port map (
            O => \N__7625\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\
        );

    \I__1462\ : CascadeMux
    port map (
            O => \N__7620\,
            I => \N__7615\
        );

    \I__1461\ : CascadeMux
    port map (
            O => \N__7619\,
            I => \N__7610\
        );

    \I__1460\ : CascadeMux
    port map (
            O => \N__7618\,
            I => \N__7607\
        );

    \I__1459\ : InMux
    port map (
            O => \N__7615\,
            I => \N__7604\
        );

    \I__1458\ : InMux
    port map (
            O => \N__7614\,
            I => \N__7597\
        );

    \I__1457\ : InMux
    port map (
            O => \N__7613\,
            I => \N__7597\
        );

    \I__1456\ : InMux
    port map (
            O => \N__7610\,
            I => \N__7597\
        );

    \I__1455\ : InMux
    port map (
            O => \N__7607\,
            I => \N__7592\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__7604\,
            I => \N__7589\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__7597\,
            I => \N__7586\
        );

    \I__1452\ : InMux
    port map (
            O => \N__7596\,
            I => \N__7583\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7595\,
            I => \N__7580\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__7592\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1449\ : Odrv4
    port map (
            O => \N__7589\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1448\ : Odrv4
    port map (
            O => \N__7586\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__7583\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__7580\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1445\ : InMux
    port map (
            O => \N__7569\,
            I => \N__7566\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__7566\,
            I => \N__7562\
        );

    \I__1443\ : InMux
    port map (
            O => \N__7565\,
            I => \N__7559\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__7562\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ0Z_0\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__7559\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ0Z_0\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__7554\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3_cascade_\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7551\,
            I => \N__7545\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7550\,
            I => \N__7542\
        );

    \I__1437\ : InMux
    port map (
            O => \N__7549\,
            I => \N__7539\
        );

    \I__1436\ : CascadeMux
    port map (
            O => \N__7548\,
            I => \N__7535\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__7545\,
            I => \N__7527\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__7542\,
            I => \N__7527\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__7539\,
            I => \N__7527\
        );

    \I__1432\ : InMux
    port map (
            O => \N__7538\,
            I => \N__7521\
        );

    \I__1431\ : InMux
    port map (
            O => \N__7535\,
            I => \N__7516\
        );

    \I__1430\ : InMux
    port map (
            O => \N__7534\,
            I => \N__7516\
        );

    \I__1429\ : Span4Mux_v
    port map (
            O => \N__7527\,
            I => \N__7513\
        );

    \I__1428\ : InMux
    port map (
            O => \N__7526\,
            I => \N__7506\
        );

    \I__1427\ : InMux
    port map (
            O => \N__7525\,
            I => \N__7506\
        );

    \I__1426\ : InMux
    port map (
            O => \N__7524\,
            I => \N__7506\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__7521\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__7516\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1423\ : Odrv4
    port map (
            O => \N__7513\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__7506\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1421\ : InMux
    port map (
            O => \N__7497\,
            I => \N__7494\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__7494\,
            I => \N__7491\
        );

    \I__1419\ : Span4Mux_h
    port map (
            O => \N__7491\,
            I => \N__7488\
        );

    \I__1418\ : Odrv4
    port map (
            O => \N__7488\,
            I => \U712_CHIP_RAM.N_433\
        );

    \I__1417\ : IoInMux
    port map (
            O => \N__7485\,
            I => \N__7482\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__7482\,
            I => \N__7479\
        );

    \I__1415\ : IoSpan4Mux
    port map (
            O => \N__7479\,
            I => \N__7476\
        );

    \I__1414\ : Span4Mux_s0_v
    port map (
            O => \N__7476\,
            I => \N__7473\
        );

    \I__1413\ : Span4Mux_v
    port map (
            O => \N__7473\,
            I => \N__7470\
        );

    \I__1412\ : Sp12to4
    port map (
            O => \N__7470\,
            I => \N__7467\
        );

    \I__1411\ : Span12Mux_h
    port map (
            O => \N__7467\,
            I => \N__7463\
        );

    \I__1410\ : InMux
    port map (
            O => \N__7466\,
            I => \N__7460\
        );

    \I__1409\ : Odrv12
    port map (
            O => \N__7463\,
            I => \LDSn_c\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__7460\,
            I => \LDSn_c\
        );

    \I__1407\ : IoInMux
    port map (
            O => \N__7455\,
            I => \N__7451\
        );

    \I__1406\ : InMux
    port map (
            O => \N__7454\,
            I => \N__7448\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__7451\,
            I => \N__7445\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__7448\,
            I => \N__7442\
        );

    \I__1403\ : Span12Mux_s4_v
    port map (
            O => \N__7445\,
            I => \N__7439\
        );

    \I__1402\ : Sp12to4
    port map (
            O => \N__7442\,
            I => \N__7436\
        );

    \I__1401\ : Span12Mux_v
    port map (
            O => \N__7439\,
            I => \N__7431\
        );

    \I__1400\ : Span12Mux_v
    port map (
            O => \N__7436\,
            I => \N__7431\
        );

    \I__1399\ : Span12Mux_h
    port map (
            O => \N__7431\,
            I => \N__7428\
        );

    \I__1398\ : Odrv12
    port map (
            O => \N__7428\,
            I => \A_c_9\
        );

    \I__1397\ : InMux
    port map (
            O => \N__7425\,
            I => \N__7422\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__7422\,
            I => \N__7419\
        );

    \I__1395\ : Span4Mux_h
    port map (
            O => \N__7419\,
            I => \N__7416\
        );

    \I__1394\ : Odrv4
    port map (
            O => \N__7416\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\
        );

    \I__1393\ : CascadeMux
    port map (
            O => \N__7413\,
            I => \N__7409\
        );

    \I__1392\ : CascadeMux
    port map (
            O => \N__7412\,
            I => \N__7406\
        );

    \I__1391\ : InMux
    port map (
            O => \N__7409\,
            I => \N__7399\
        );

    \I__1390\ : InMux
    port map (
            O => \N__7406\,
            I => \N__7399\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__7405\,
            I => \N__7392\
        );

    \I__1388\ : CascadeMux
    port map (
            O => \N__7404\,
            I => \N__7389\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__7399\,
            I => \N__7381\
        );

    \I__1386\ : CascadeMux
    port map (
            O => \N__7398\,
            I => \N__7374\
        );

    \I__1385\ : InMux
    port map (
            O => \N__7397\,
            I => \N__7366\
        );

    \I__1384\ : InMux
    port map (
            O => \N__7396\,
            I => \N__7366\
        );

    \I__1383\ : InMux
    port map (
            O => \N__7395\,
            I => \N__7366\
        );

    \I__1382\ : InMux
    port map (
            O => \N__7392\,
            I => \N__7363\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7389\,
            I => \N__7360\
        );

    \I__1380\ : InMux
    port map (
            O => \N__7388\,
            I => \N__7355\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7387\,
            I => \N__7355\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7348\
        );

    \I__1377\ : InMux
    port map (
            O => \N__7385\,
            I => \N__7348\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7384\,
            I => \N__7348\
        );

    \I__1375\ : Span4Mux_h
    port map (
            O => \N__7381\,
            I => \N__7345\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7380\,
            I => \N__7336\
        );

    \I__1373\ : InMux
    port map (
            O => \N__7379\,
            I => \N__7336\
        );

    \I__1372\ : InMux
    port map (
            O => \N__7378\,
            I => \N__7336\
        );

    \I__1371\ : InMux
    port map (
            O => \N__7377\,
            I => \N__7336\
        );

    \I__1370\ : InMux
    port map (
            O => \N__7374\,
            I => \N__7331\
        );

    \I__1369\ : InMux
    port map (
            O => \N__7373\,
            I => \N__7331\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__7366\,
            I => \U712_CHIP_RAM.N_476\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__7363\,
            I => \U712_CHIP_RAM.N_476\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__7360\,
            I => \U712_CHIP_RAM.N_476\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__7355\,
            I => \U712_CHIP_RAM.N_476\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__7348\,
            I => \U712_CHIP_RAM.N_476\
        );

    \I__1363\ : Odrv4
    port map (
            O => \N__7345\,
            I => \U712_CHIP_RAM.N_476\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__7336\,
            I => \U712_CHIP_RAM.N_476\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__7331\,
            I => \U712_CHIP_RAM.N_476\
        );

    \I__1360\ : InMux
    port map (
            O => \N__7314\,
            I => \N__7311\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__7311\,
            I => \U712_CHIP_RAM.N_446\
        );

    \I__1358\ : InMux
    port map (
            O => \N__7308\,
            I => \N__7302\
        );

    \I__1357\ : InMux
    port map (
            O => \N__7307\,
            I => \N__7298\
        );

    \I__1356\ : InMux
    port map (
            O => \N__7306\,
            I => \N__7295\
        );

    \I__1355\ : InMux
    port map (
            O => \N__7305\,
            I => \N__7290\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__7302\,
            I => \N__7285\
        );

    \I__1353\ : InMux
    port map (
            O => \N__7301\,
            I => \N__7282\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__7298\,
            I => \N__7277\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__7295\,
            I => \N__7277\
        );

    \I__1350\ : InMux
    port map (
            O => \N__7294\,
            I => \N__7274\
        );

    \I__1349\ : InMux
    port map (
            O => \N__7293\,
            I => \N__7271\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__7290\,
            I => \N__7268\
        );

    \I__1347\ : CascadeMux
    port map (
            O => \N__7289\,
            I => \N__7259\
        );

    \I__1346\ : InMux
    port map (
            O => \N__7288\,
            I => \N__7255\
        );

    \I__1345\ : Span4Mux_v
    port map (
            O => \N__7285\,
            I => \N__7248\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__7282\,
            I => \N__7248\
        );

    \I__1343\ : Span4Mux_v
    port map (
            O => \N__7277\,
            I => \N__7248\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__7274\,
            I => \N__7241\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__7271\,
            I => \N__7241\
        );

    \I__1340\ : Span4Mux_h
    port map (
            O => \N__7268\,
            I => \N__7241\
        );

    \I__1339\ : InMux
    port map (
            O => \N__7267\,
            I => \N__7236\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7266\,
            I => \N__7236\
        );

    \I__1337\ : InMux
    port map (
            O => \N__7265\,
            I => \N__7231\
        );

    \I__1336\ : InMux
    port map (
            O => \N__7264\,
            I => \N__7231\
        );

    \I__1335\ : InMux
    port map (
            O => \N__7263\,
            I => \N__7224\
        );

    \I__1334\ : InMux
    port map (
            O => \N__7262\,
            I => \N__7224\
        );

    \I__1333\ : InMux
    port map (
            O => \N__7259\,
            I => \N__7224\
        );

    \I__1332\ : InMux
    port map (
            O => \N__7258\,
            I => \N__7221\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__7255\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1330\ : Odrv4
    port map (
            O => \N__7248\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1329\ : Odrv4
    port map (
            O => \N__7241\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__7236\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__7231\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__7224\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__7221\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1324\ : InMux
    port map (
            O => \N__7206\,
            I => \N__7198\
        );

    \I__1323\ : InMux
    port map (
            O => \N__7205\,
            I => \N__7195\
        );

    \I__1322\ : InMux
    port map (
            O => \N__7204\,
            I => \N__7192\
        );

    \I__1321\ : CascadeMux
    port map (
            O => \N__7203\,
            I => \N__7187\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__7202\,
            I => \N__7184\
        );

    \I__1319\ : InMux
    port map (
            O => \N__7201\,
            I => \N__7180\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__7198\,
            I => \N__7177\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__7195\,
            I => \N__7174\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__7192\,
            I => \N__7167\
        );

    \I__1315\ : InMux
    port map (
            O => \N__7191\,
            I => \N__7164\
        );

    \I__1314\ : InMux
    port map (
            O => \N__7190\,
            I => \N__7160\
        );

    \I__1313\ : InMux
    port map (
            O => \N__7187\,
            I => \N__7157\
        );

    \I__1312\ : InMux
    port map (
            O => \N__7184\,
            I => \N__7154\
        );

    \I__1311\ : InMux
    port map (
            O => \N__7183\,
            I => \N__7151\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__7180\,
            I => \N__7148\
        );

    \I__1309\ : Span4Mux_v
    port map (
            O => \N__7177\,
            I => \N__7143\
        );

    \I__1308\ : Span4Mux_v
    port map (
            O => \N__7174\,
            I => \N__7143\
        );

    \I__1307\ : InMux
    port map (
            O => \N__7173\,
            I => \N__7138\
        );

    \I__1306\ : InMux
    port map (
            O => \N__7172\,
            I => \N__7138\
        );

    \I__1305\ : InMux
    port map (
            O => \N__7171\,
            I => \N__7133\
        );

    \I__1304\ : InMux
    port map (
            O => \N__7170\,
            I => \N__7133\
        );

    \I__1303\ : Span4Mux_v
    port map (
            O => \N__7167\,
            I => \N__7128\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__7164\,
            I => \N__7128\
        );

    \I__1301\ : InMux
    port map (
            O => \N__7163\,
            I => \N__7125\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__7160\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__7157\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__7154\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__7151\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1296\ : Odrv4
    port map (
            O => \N__7148\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1295\ : Odrv4
    port map (
            O => \N__7143\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__7138\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__7133\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1292\ : Odrv4
    port map (
            O => \N__7128\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__7125\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__7104\,
            I => \N__7099\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__7103\,
            I => \N__7094\
        );

    \I__1288\ : CascadeMux
    port map (
            O => \N__7102\,
            I => \N__7091\
        );

    \I__1287\ : InMux
    port map (
            O => \N__7099\,
            I => \N__7087\
        );

    \I__1286\ : InMux
    port map (
            O => \N__7098\,
            I => \N__7084\
        );

    \I__1285\ : InMux
    port map (
            O => \N__7097\,
            I => \N__7081\
        );

    \I__1284\ : InMux
    port map (
            O => \N__7094\,
            I => \N__7072\
        );

    \I__1283\ : InMux
    port map (
            O => \N__7091\,
            I => \N__7067\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__7090\,
            I => \N__7064\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__7087\,
            I => \N__7061\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__7084\,
            I => \N__7056\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__7081\,
            I => \N__7056\
        );

    \I__1278\ : InMux
    port map (
            O => \N__7080\,
            I => \N__7051\
        );

    \I__1277\ : InMux
    port map (
            O => \N__7079\,
            I => \N__7051\
        );

    \I__1276\ : InMux
    port map (
            O => \N__7078\,
            I => \N__7048\
        );

    \I__1275\ : InMux
    port map (
            O => \N__7077\,
            I => \N__7044\
        );

    \I__1274\ : InMux
    port map (
            O => \N__7076\,
            I => \N__7041\
        );

    \I__1273\ : InMux
    port map (
            O => \N__7075\,
            I => \N__7038\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__7072\,
            I => \N__7035\
        );

    \I__1271\ : InMux
    port map (
            O => \N__7071\,
            I => \N__7030\
        );

    \I__1270\ : InMux
    port map (
            O => \N__7070\,
            I => \N__7030\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__7067\,
            I => \N__7027\
        );

    \I__1268\ : InMux
    port map (
            O => \N__7064\,
            I => \N__7024\
        );

    \I__1267\ : Span4Mux_v
    port map (
            O => \N__7061\,
            I => \N__7017\
        );

    \I__1266\ : Span4Mux_v
    port map (
            O => \N__7056\,
            I => \N__7017\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__7051\,
            I => \N__7017\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__7048\,
            I => \N__7014\
        );

    \I__1263\ : InMux
    port map (
            O => \N__7047\,
            I => \N__7011\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__7044\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__7041\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__7038\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1259\ : Odrv4
    port map (
            O => \N__7035\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__7030\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1257\ : Odrv12
    port map (
            O => \N__7027\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__7024\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1255\ : Odrv4
    port map (
            O => \N__7017\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1254\ : Odrv4
    port map (
            O => \N__7014\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__7011\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1252\ : InMux
    port map (
            O => \N__6990\,
            I => \N__6984\
        );

    \I__1251\ : InMux
    port map (
            O => \N__6989\,
            I => \N__6981\
        );

    \I__1250\ : InMux
    port map (
            O => \N__6988\,
            I => \N__6976\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6987\,
            I => \N__6976\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__6984\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__6981\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__6976\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1245\ : InMux
    port map (
            O => \N__6969\,
            I => \N__6966\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__6966\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_i_i_a2_1_0\
        );

    \I__1243\ : CascadeMux
    port map (
            O => \N__6963\,
            I => \N__6958\
        );

    \I__1242\ : CascadeMux
    port map (
            O => \N__6962\,
            I => \N__6955\
        );

    \I__1241\ : InMux
    port map (
            O => \N__6961\,
            I => \N__6951\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6958\,
            I => \N__6948\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6955\,
            I => \N__6943\
        );

    \I__1238\ : InMux
    port map (
            O => \N__6954\,
            I => \N__6943\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__6951\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__6948\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6943\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1234\ : InMux
    port map (
            O => \N__6936\,
            I => \N__6933\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__6933\,
            I => \U712_CHIP_RAM.N_431\
        );

    \I__1232\ : InMux
    port map (
            O => \N__6930\,
            I => \N__6927\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__6927\,
            I => \N__6924\
        );

    \I__1230\ : Span4Mux_h
    port map (
            O => \N__6924\,
            I => \N__6921\
        );

    \I__1229\ : Sp12to4
    port map (
            O => \N__6921\,
            I => \N__6918\
        );

    \I__1228\ : Span12Mux_v
    port map (
            O => \N__6918\,
            I => \N__6915\
        );

    \I__1227\ : Odrv12
    port map (
            O => \N__6915\,
            I => \A_c_15\
        );

    \I__1226\ : InMux
    port map (
            O => \N__6912\,
            I => \N__6909\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__6909\,
            I => \N__6906\
        );

    \I__1224\ : Odrv12
    port map (
            O => \N__6906\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\
        );

    \I__1223\ : InMux
    port map (
            O => \N__6903\,
            I => \N__6894\
        );

    \I__1222\ : InMux
    port map (
            O => \N__6902\,
            I => \N__6894\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6901\,
            I => \N__6894\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6894\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\
        );

    \I__1219\ : IoInMux
    port map (
            O => \N__6891\,
            I => \N__6888\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__6888\,
            I => \N__6885\
        );

    \I__1217\ : IoSpan4Mux
    port map (
            O => \N__6885\,
            I => \N__6882\
        );

    \I__1216\ : Span4Mux_s2_v
    port map (
            O => \N__6882\,
            I => \N__6878\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6875\
        );

    \I__1214\ : Sp12to4
    port map (
            O => \N__6878\,
            I => \N__6872\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__6875\,
            I => \N__6869\
        );

    \I__1212\ : Span12Mux_s8_v
    port map (
            O => \N__6872\,
            I => \N__6866\
        );

    \I__1211\ : Span4Mux_v
    port map (
            O => \N__6869\,
            I => \N__6863\
        );

    \I__1210\ : Span12Mux_v
    port map (
            O => \N__6866\,
            I => \N__6860\
        );

    \I__1209\ : Sp12to4
    port map (
            O => \N__6863\,
            I => \N__6857\
        );

    \I__1208\ : Span12Mux_h
    port map (
            O => \N__6860\,
            I => \N__6854\
        );

    \I__1207\ : Span12Mux_h
    port map (
            O => \N__6857\,
            I => \N__6851\
        );

    \I__1206\ : Odrv12
    port map (
            O => \N__6854\,
            I => \A_c_11\
        );

    \I__1205\ : Odrv12
    port map (
            O => \N__6851\,
            I => \A_c_11\
        );

    \I__1204\ : InMux
    port map (
            O => \N__6846\,
            I => \N__6843\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__6843\,
            I => \N__6840\
        );

    \I__1202\ : Odrv4
    port map (
            O => \N__6840\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\
        );

    \I__1201\ : InMux
    port map (
            O => \N__6837\,
            I => \N__6831\
        );

    \I__1200\ : InMux
    port map (
            O => \N__6836\,
            I => \N__6831\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__6831\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1198\ : InMux
    port map (
            O => \N__6828\,
            I => \N__6825\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6825\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\
        );

    \I__1196\ : CascadeMux
    port map (
            O => \N__6822\,
            I => \N__6815\
        );

    \I__1195\ : InMux
    port map (
            O => \N__6821\,
            I => \N__6810\
        );

    \I__1194\ : InMux
    port map (
            O => \N__6820\,
            I => \N__6803\
        );

    \I__1193\ : InMux
    port map (
            O => \N__6819\,
            I => \N__6803\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6818\,
            I => \N__6803\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6815\,
            I => \N__6800\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6814\,
            I => \N__6797\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6813\,
            I => \N__6794\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__6810\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__6803\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__6800\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__6797\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6794\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1183\ : InMux
    port map (
            O => \N__6783\,
            I => \N__6780\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__6780\,
            I => \N__6776\
        );

    \I__1181\ : InMux
    port map (
            O => \N__6779\,
            I => \N__6773\
        );

    \I__1180\ : Odrv12
    port map (
            O => \N__6776\,
            I => \U712_CHIP_RAM.N_326\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__6773\,
            I => \U712_CHIP_RAM.N_326\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__6768\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_i_a2_0_1_cascade_\
        );

    \I__1177\ : InMux
    port map (
            O => \N__6765\,
            I => \N__6762\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__6762\,
            I => \N__6758\
        );

    \I__1175\ : InMux
    port map (
            O => \N__6761\,
            I => \N__6755\
        );

    \I__1174\ : Odrv4
    port map (
            O => \N__6758\,
            I => \U712_CHIP_RAM.N_572\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__6755\,
            I => \U712_CHIP_RAM.N_572\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6750\,
            I => \N__6747\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__6747\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER19\
        );

    \I__1170\ : InMux
    port map (
            O => \N__6744\,
            I => \N__6741\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__6741\,
            I => \U712_CHIP_RAM.N_574\
        );

    \I__1168\ : CascadeMux
    port map (
            O => \N__6738\,
            I => \N__6735\
        );

    \I__1167\ : InMux
    port map (
            O => \N__6735\,
            I => \N__6732\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6732\,
            I => \U712_CHIP_RAM.N_571\
        );

    \I__1165\ : CascadeMux
    port map (
            O => \N__6729\,
            I => \N__6726\
        );

    \I__1164\ : InMux
    port map (
            O => \N__6726\,
            I => \N__6721\
        );

    \I__1163\ : InMux
    port map (
            O => \N__6725\,
            I => \N__6718\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6724\,
            I => \N__6715\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__6721\,
            I => \U712_CHIP_RAM.N_566\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__6718\,
            I => \U712_CHIP_RAM.N_566\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__6715\,
            I => \U712_CHIP_RAM.N_566\
        );

    \I__1158\ : InMux
    port map (
            O => \N__6708\,
            I => \N__6705\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__6705\,
            I => \N__6701\
        );

    \I__1156\ : InMux
    port map (
            O => \N__6704\,
            I => \N__6698\
        );

    \I__1155\ : Span4Mux_h
    port map (
            O => \N__6701\,
            I => \N__6694\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__6698\,
            I => \N__6691\
        );

    \I__1153\ : InMux
    port map (
            O => \N__6697\,
            I => \N__6688\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__6694\,
            I => \U712_CHIP_RAM.N_477\
        );

    \I__1151\ : Odrv4
    port map (
            O => \N__6691\,
            I => \U712_CHIP_RAM.N_477\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__6688\,
            I => \U712_CHIP_RAM.N_477\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6681\,
            I => \N__6668\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6680\,
            I => \N__6665\
        );

    \I__1147\ : InMux
    port map (
            O => \N__6679\,
            I => \N__6662\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6678\,
            I => \N__6659\
        );

    \I__1145\ : InMux
    port map (
            O => \N__6677\,
            I => \N__6652\
        );

    \I__1144\ : InMux
    port map (
            O => \N__6676\,
            I => \N__6652\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6652\
        );

    \I__1142\ : CascadeMux
    port map (
            O => \N__6674\,
            I => \N__6641\
        );

    \I__1141\ : CascadeMux
    port map (
            O => \N__6673\,
            I => \N__6637\
        );

    \I__1140\ : CascadeMux
    port map (
            O => \N__6672\,
            I => \N__6633\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6671\,
            I => \N__6629\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__6668\,
            I => \N__6626\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__6665\,
            I => \N__6623\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6662\,
            I => \N__6616\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__6659\,
            I => \N__6616\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__6652\,
            I => \N__6616\
        );

    \I__1133\ : InMux
    port map (
            O => \N__6651\,
            I => \N__6609\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6650\,
            I => \N__6606\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6649\,
            I => \N__6599\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6648\,
            I => \N__6599\
        );

    \I__1129\ : InMux
    port map (
            O => \N__6647\,
            I => \N__6599\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6646\,
            I => \N__6594\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6645\,
            I => \N__6594\
        );

    \I__1126\ : InMux
    port map (
            O => \N__6644\,
            I => \N__6583\
        );

    \I__1125\ : InMux
    port map (
            O => \N__6641\,
            I => \N__6583\
        );

    \I__1124\ : InMux
    port map (
            O => \N__6640\,
            I => \N__6583\
        );

    \I__1123\ : InMux
    port map (
            O => \N__6637\,
            I => \N__6583\
        );

    \I__1122\ : InMux
    port map (
            O => \N__6636\,
            I => \N__6583\
        );

    \I__1121\ : InMux
    port map (
            O => \N__6633\,
            I => \N__6578\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6632\,
            I => \N__6578\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__6629\,
            I => \N__6569\
        );

    \I__1118\ : Span4Mux_h
    port map (
            O => \N__6626\,
            I => \N__6569\
        );

    \I__1117\ : Span4Mux_v
    port map (
            O => \N__6623\,
            I => \N__6569\
        );

    \I__1116\ : Span4Mux_v
    port map (
            O => \N__6616\,
            I => \N__6569\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6615\,
            I => \N__6560\
        );

    \I__1114\ : InMux
    port map (
            O => \N__6614\,
            I => \N__6560\
        );

    \I__1113\ : InMux
    port map (
            O => \N__6613\,
            I => \N__6560\
        );

    \I__1112\ : InMux
    port map (
            O => \N__6612\,
            I => \N__6560\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__6609\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6606\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__6599\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6594\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__6583\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__6578\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1105\ : Odrv4
    port map (
            O => \N__6569\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__6560\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1103\ : InMux
    port map (
            O => \N__6543\,
            I => \N__6535\
        );

    \I__1102\ : InMux
    port map (
            O => \N__6542\,
            I => \N__6535\
        );

    \I__1101\ : InMux
    port map (
            O => \N__6541\,
            I => \N__6530\
        );

    \I__1100\ : InMux
    port map (
            O => \N__6540\,
            I => \N__6530\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__6535\,
            I => \U712_CHIP_RAM.N_555\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__6530\,
            I => \U712_CHIP_RAM.N_555\
        );

    \I__1097\ : InMux
    port map (
            O => \N__6525\,
            I => \N__6522\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__6522\,
            I => \U712_CHIP_RAM.N_349\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6519\,
            I => \N__6516\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6516\,
            I => \U712_CHIP_RAM.N_447\
        );

    \I__1093\ : CascadeMux
    port map (
            O => \N__6513\,
            I => \U712_CHIP_RAM.N_444_cascade_\
        );

    \I__1092\ : InMux
    port map (
            O => \N__6510\,
            I => \N__6507\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__6507\,
            I => \N__6503\
        );

    \I__1090\ : InMux
    port map (
            O => \N__6506\,
            I => \N__6500\
        );

    \I__1089\ : Odrv4
    port map (
            O => \N__6503\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__6500\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6495\,
            I => \N__6489\
        );

    \I__1086\ : InMux
    port map (
            O => \N__6494\,
            I => \N__6489\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__6489\,
            I => \U712_CHIP_RAM.N_410\
        );

    \I__1084\ : InMux
    port map (
            O => \N__6486\,
            I => \N__6483\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__6483\,
            I => \U712_CHIP_RAM.N_411\
        );

    \I__1082\ : CascadeMux
    port map (
            O => \N__6480\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\
        );

    \I__1081\ : InMux
    port map (
            O => \N__6477\,
            I => \N__6473\
        );

    \I__1080\ : InMux
    port map (
            O => \N__6476\,
            I => \N__6470\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__6473\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__6470\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__1077\ : CascadeMux
    port map (
            O => \N__6465\,
            I => \N__6460\
        );

    \I__1076\ : InMux
    port map (
            O => \N__6464\,
            I => \N__6449\
        );

    \I__1075\ : InMux
    port map (
            O => \N__6463\,
            I => \N__6449\
        );

    \I__1074\ : InMux
    port map (
            O => \N__6460\,
            I => \N__6449\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6459\,
            I => \N__6446\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6458\,
            I => \N__6441\
        );

    \I__1071\ : InMux
    port map (
            O => \N__6457\,
            I => \N__6441\
        );

    \I__1070\ : InMux
    port map (
            O => \N__6456\,
            I => \N__6438\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__6449\,
            I => \N__6435\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__6446\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__6441\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__6438\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__1065\ : Odrv4
    port map (
            O => \N__6435\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6426\,
            I => \N__6423\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__6423\,
            I => \N__6420\
        );

    \I__1062\ : Odrv4
    port map (
            O => \N__6420\,
            I => \U712_REG_SM.STATE_COUNTsr_0\
        );

    \I__1061\ : InMux
    port map (
            O => \N__6417\,
            I => \N__6412\
        );

    \I__1060\ : InMux
    port map (
            O => \N__6416\,
            I => \N__6407\
        );

    \I__1059\ : InMux
    port map (
            O => \N__6415\,
            I => \N__6407\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__6412\,
            I => \U712_REG_SM.N_338\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__6407\,
            I => \U712_REG_SM.N_338\
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__6402\,
            I => \N__6397\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6401\,
            I => \N__6393\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6400\,
            I => \N__6390\
        );

    \I__1053\ : InMux
    port map (
            O => \N__6397\,
            I => \N__6385\
        );

    \I__1052\ : InMux
    port map (
            O => \N__6396\,
            I => \N__6385\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__6393\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__6390\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__6385\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1048\ : IoInMux
    port map (
            O => \N__6378\,
            I => \N__6375\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__6375\,
            I => \N__6372\
        );

    \I__1046\ : Span4Mux_s3_v
    port map (
            O => \N__6372\,
            I => \N__6369\
        );

    \I__1045\ : Span4Mux_v
    port map (
            O => \N__6369\,
            I => \N__6366\
        );

    \I__1044\ : Sp12to4
    port map (
            O => \N__6366\,
            I => \N__6362\
        );

    \I__1043\ : CascadeMux
    port map (
            O => \N__6365\,
            I => \N__6359\
        );

    \I__1042\ : Span12Mux_h
    port map (
            O => \N__6362\,
            I => \N__6356\
        );

    \I__1041\ : InMux
    port map (
            O => \N__6359\,
            I => \N__6353\
        );

    \I__1040\ : Odrv12
    port map (
            O => \N__6356\,
            I => \UDSn_c\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__6353\,
            I => \UDSn_c\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6348\,
            I => \N__6345\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__6345\,
            I => \U712_REG_SM.N_435\
        );

    \I__1036\ : IoInMux
    port map (
            O => \N__6342\,
            I => \N__6339\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__6339\,
            I => \N__6336\
        );

    \I__1034\ : Span12Mux_s8_v
    port map (
            O => \N__6336\,
            I => \N__6332\
        );

    \I__1033\ : InMux
    port map (
            O => \N__6335\,
            I => \N__6329\
        );

    \I__1032\ : Odrv12
    port map (
            O => \N__6332\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__6329\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6324\,
            I => \N__6321\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6321\,
            I => \N__6318\
        );

    \I__1028\ : Odrv4
    port map (
            O => \N__6318\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__1027\ : InMux
    port map (
            O => \N__6315\,
            I => \N__6312\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__6312\,
            I => \U712_CHIP_RAM.N_320\
        );

    \I__1025\ : InMux
    port map (
            O => \N__6309\,
            I => \N__6302\
        );

    \I__1024\ : CascadeMux
    port map (
            O => \N__6308\,
            I => \N__6297\
        );

    \I__1023\ : InMux
    port map (
            O => \N__6307\,
            I => \N__6289\
        );

    \I__1022\ : InMux
    port map (
            O => \N__6306\,
            I => \N__6289\
        );

    \I__1021\ : InMux
    port map (
            O => \N__6305\,
            I => \N__6289\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__6302\,
            I => \N__6286\
        );

    \I__1019\ : InMux
    port map (
            O => \N__6301\,
            I => \N__6283\
        );

    \I__1018\ : InMux
    port map (
            O => \N__6300\,
            I => \N__6280\
        );

    \I__1017\ : InMux
    port map (
            O => \N__6297\,
            I => \N__6273\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6296\,
            I => \N__6273\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__6289\,
            I => \N__6270\
        );

    \I__1014\ : Span4Mux_h
    port map (
            O => \N__6286\,
            I => \N__6267\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__6283\,
            I => \N__6262\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__6280\,
            I => \N__6262\
        );

    \I__1011\ : InMux
    port map (
            O => \N__6279\,
            I => \N__6257\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6278\,
            I => \N__6257\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__6273\,
            I => \N__6254\
        );

    \I__1008\ : Span4Mux_v
    port map (
            O => \N__6270\,
            I => \N__6251\
        );

    \I__1007\ : Odrv4
    port map (
            O => \N__6267\,
            I => \U712_CHIP_RAM.N_480\
        );

    \I__1006\ : Odrv4
    port map (
            O => \N__6262\,
            I => \U712_CHIP_RAM.N_480\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__6257\,
            I => \U712_CHIP_RAM.N_480\
        );

    \I__1004\ : Odrv12
    port map (
            O => \N__6254\,
            I => \U712_CHIP_RAM.N_480\
        );

    \I__1003\ : Odrv4
    port map (
            O => \N__6251\,
            I => \U712_CHIP_RAM.N_480\
        );

    \I__1002\ : CascadeMux
    port map (
            O => \N__6240\,
            I => \U712_CHIP_RAM.N_571_cascade_\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6237\,
            I => \N__6228\
        );

    \I__1000\ : InMux
    port map (
            O => \N__6236\,
            I => \N__6228\
        );

    \I__999\ : InMux
    port map (
            O => \N__6235\,
            I => \N__6228\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__6228\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__997\ : InMux
    port map (
            O => \N__6225\,
            I => \N__6222\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__6222\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\
        );

    \I__995\ : CascadeMux
    port map (
            O => \N__6219\,
            I => \N__6214\
        );

    \I__994\ : InMux
    port map (
            O => \N__6218\,
            I => \N__6210\
        );

    \I__993\ : CascadeMux
    port map (
            O => \N__6217\,
            I => \N__6207\
        );

    \I__992\ : InMux
    port map (
            O => \N__6214\,
            I => \N__6202\
        );

    \I__991\ : InMux
    port map (
            O => \N__6213\,
            I => \N__6202\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__6210\,
            I => \N__6199\
        );

    \I__989\ : InMux
    port map (
            O => \N__6207\,
            I => \N__6196\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__6202\,
            I => \N__6193\
        );

    \I__987\ : Span4Mux_h
    port map (
            O => \N__6199\,
            I => \N__6190\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__6196\,
            I => \REG_TACK\
        );

    \I__985\ : Odrv4
    port map (
            O => \N__6193\,
            I => \REG_TACK\
        );

    \I__984\ : Odrv4
    port map (
            O => \N__6190\,
            I => \REG_TACK\
        );

    \I__983\ : InMux
    port map (
            O => \N__6183\,
            I => \N__6178\
        );

    \I__982\ : InMux
    port map (
            O => \N__6182\,
            I => \N__6173\
        );

    \I__981\ : InMux
    port map (
            O => \N__6181\,
            I => \N__6173\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__6178\,
            I => \N__6170\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__6173\,
            I => \N__6166\
        );

    \I__978\ : Span4Mux_h
    port map (
            O => \N__6170\,
            I => \N__6163\
        );

    \I__977\ : InMux
    port map (
            O => \N__6169\,
            I => \N__6160\
        );

    \I__976\ : Span4Mux_v
    port map (
            O => \N__6166\,
            I => \N__6157\
        );

    \I__975\ : Span4Mux_v
    port map (
            O => \N__6163\,
            I => \N__6154\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__6160\,
            I => \CPU_TACKm\
        );

    \I__973\ : Odrv4
    port map (
            O => \N__6157\,
            I => \CPU_TACKm\
        );

    \I__972\ : Odrv4
    port map (
            O => \N__6154\,
            I => \CPU_TACKm\
        );

    \I__971\ : InMux
    port map (
            O => \N__6147\,
            I => \N__6144\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__6144\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__969\ : IoInMux
    port map (
            O => \N__6141\,
            I => \N__6138\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__6138\,
            I => \N__6134\
        );

    \I__967\ : IoInMux
    port map (
            O => \N__6137\,
            I => \N__6131\
        );

    \I__966\ : IoSpan4Mux
    port map (
            O => \N__6134\,
            I => \N__6126\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__6131\,
            I => \N__6126\
        );

    \I__964\ : IoSpan4Mux
    port map (
            O => \N__6126\,
            I => \N__6122\
        );

    \I__963\ : IoInMux
    port map (
            O => \N__6125\,
            I => \N__6119\
        );

    \I__962\ : Span4Mux_s1_v
    port map (
            O => \N__6122\,
            I => \N__6116\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__6119\,
            I => \N__6113\
        );

    \I__960\ : Span4Mux_v
    port map (
            O => \N__6116\,
            I => \N__6110\
        );

    \I__959\ : IoSpan4Mux
    port map (
            O => \N__6113\,
            I => \N__6107\
        );

    \I__958\ : Sp12to4
    port map (
            O => \N__6110\,
            I => \N__6104\
        );

    \I__957\ : Sp12to4
    port map (
            O => \N__6107\,
            I => \N__6101\
        );

    \I__956\ : Span12Mux_h
    port map (
            O => \N__6104\,
            I => \N__6096\
        );

    \I__955\ : Span12Mux_h
    port map (
            O => \N__6101\,
            I => \N__6096\
        );

    \I__954\ : Odrv12
    port map (
            O => \N__6096\,
            I => \CLK40_PLL_i_i\
        );

    \I__953\ : InMux
    port map (
            O => \N__6093\,
            I => \N__6084\
        );

    \I__952\ : InMux
    port map (
            O => \N__6092\,
            I => \N__6079\
        );

    \I__951\ : InMux
    port map (
            O => \N__6091\,
            I => \N__6079\
        );

    \I__950\ : CascadeMux
    port map (
            O => \N__6090\,
            I => \N__6074\
        );

    \I__949\ : InMux
    port map (
            O => \N__6089\,
            I => \N__6069\
        );

    \I__948\ : InMux
    port map (
            O => \N__6088\,
            I => \N__6064\
        );

    \I__947\ : InMux
    port map (
            O => \N__6087\,
            I => \N__6064\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__6084\,
            I => \N__6059\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__6079\,
            I => \N__6059\
        );

    \I__944\ : InMux
    port map (
            O => \N__6078\,
            I => \N__6054\
        );

    \I__943\ : InMux
    port map (
            O => \N__6077\,
            I => \N__6054\
        );

    \I__942\ : InMux
    port map (
            O => \N__6074\,
            I => \N__6047\
        );

    \I__941\ : InMux
    port map (
            O => \N__6073\,
            I => \N__6047\
        );

    \I__940\ : InMux
    port map (
            O => \N__6072\,
            I => \N__6047\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__6069\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__6064\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__937\ : Odrv4
    port map (
            O => \N__6059\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__6054\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__6047\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__934\ : InMux
    port map (
            O => \N__6036\,
            I => \N__6033\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__6033\,
            I => \N__6030\
        );

    \I__932\ : Span4Mux_v
    port map (
            O => \N__6030\,
            I => \N__6027\
        );

    \I__931\ : Odrv4
    port map (
            O => \N__6027\,
            I => \U712_REG_SM.N_416\
        );

    \I__930\ : InMux
    port map (
            O => \N__6024\,
            I => \N__6018\
        );

    \I__929\ : InMux
    port map (
            O => \N__6023\,
            I => \N__6011\
        );

    \I__928\ : InMux
    port map (
            O => \N__6022\,
            I => \N__6011\
        );

    \I__927\ : InMux
    port map (
            O => \N__6021\,
            I => \N__6011\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__6018\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__6011\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__924\ : CascadeMux
    port map (
            O => \N__6006\,
            I => \N__6001\
        );

    \I__923\ : InMux
    port map (
            O => \N__6005\,
            I => \N__5998\
        );

    \I__922\ : InMux
    port map (
            O => \N__6004\,
            I => \N__5995\
        );

    \I__921\ : InMux
    port map (
            O => \N__6001\,
            I => \N__5992\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__5998\,
            I => \N__5989\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__5995\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5992\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__917\ : Odrv12
    port map (
            O => \N__5989\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__916\ : InMux
    port map (
            O => \N__5982\,
            I => \N__5977\
        );

    \I__915\ : InMux
    port map (
            O => \N__5981\,
            I => \N__5972\
        );

    \I__914\ : InMux
    port map (
            O => \N__5980\,
            I => \N__5972\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__5977\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__5972\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__911\ : CascadeMux
    port map (
            O => \N__5967\,
            I => \N__5964\
        );

    \I__910\ : InMux
    port map (
            O => \N__5964\,
            I => \N__5959\
        );

    \I__909\ : InMux
    port map (
            O => \N__5963\,
            I => \N__5954\
        );

    \I__908\ : InMux
    port map (
            O => \N__5962\,
            I => \N__5951\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__5959\,
            I => \N__5948\
        );

    \I__906\ : InMux
    port map (
            O => \N__5958\,
            I => \N__5943\
        );

    \I__905\ : InMux
    port map (
            O => \N__5957\,
            I => \N__5943\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__5954\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5951\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__902\ : Odrv4
    port map (
            O => \N__5948\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__5943\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__900\ : InMux
    port map (
            O => \N__5934\,
            I => \N__5931\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__5931\,
            I => \N__5927\
        );

    \I__898\ : InMux
    port map (
            O => \N__5930\,
            I => \N__5924\
        );

    \I__897\ : Span4Mux_h
    port map (
            O => \N__5927\,
            I => \N__5921\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__5924\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__895\ : Odrv4
    port map (
            O => \N__5921\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__894\ : CascadeMux
    port map (
            O => \N__5916\,
            I => \N__5913\
        );

    \I__893\ : InMux
    port map (
            O => \N__5913\,
            I => \N__5910\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__5910\,
            I => \N__5907\
        );

    \I__891\ : Odrv4
    port map (
            O => \N__5907\,
            I => \U712_CHIP_RAM.REFRESH5lto7_0\
        );

    \I__890\ : InMux
    port map (
            O => \N__5904\,
            I => \N__5901\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__5901\,
            I => \N__5898\
        );

    \I__888\ : Span4Mux_h
    port map (
            O => \N__5898\,
            I => \N__5895\
        );

    \I__887\ : Odrv4
    port map (
            O => \N__5895\,
            I => \U712_CHIP_RAM.REFRESH5lt7\
        );

    \I__886\ : InMux
    port map (
            O => \N__5892\,
            I => \N__5889\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5889\,
            I => \N__5886\
        );

    \I__884\ : Odrv4
    port map (
            O => \N__5886\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3\
        );

    \I__883\ : InMux
    port map (
            O => \N__5883\,
            I => \N__5880\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__5880\,
            I => \U712_CHIP_RAM.N_327\
        );

    \I__881\ : InMux
    port map (
            O => \N__5877\,
            I => \N__5874\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__5874\,
            I => \N__5871\
        );

    \I__879\ : Span4Mux_h
    port map (
            O => \N__5871\,
            I => \N__5867\
        );

    \I__878\ : InMux
    port map (
            O => \N__5870\,
            I => \N__5864\
        );

    \I__877\ : Span4Mux_h
    port map (
            O => \N__5867\,
            I => \N__5861\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__5864\,
            I => \N__5858\
        );

    \I__875\ : Sp12to4
    port map (
            O => \N__5861\,
            I => \N__5853\
        );

    \I__874\ : Span12Mux_h
    port map (
            O => \N__5858\,
            I => \N__5853\
        );

    \I__873\ : Span12Mux_v
    port map (
            O => \N__5853\,
            I => \N__5850\
        );

    \I__872\ : Odrv12
    port map (
            O => \N__5850\,
            I => \TSn_c\
        );

    \I__871\ : InMux
    port map (
            O => \N__5847\,
            I => \N__5844\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__5844\,
            I => \N__5841\
        );

    \I__869\ : Span4Mux_h
    port map (
            O => \N__5841\,
            I => \N__5838\
        );

    \I__868\ : Sp12to4
    port map (
            O => \N__5838\,
            I => \N__5835\
        );

    \I__867\ : Span12Mux_v
    port map (
            O => \N__5835\,
            I => \N__5832\
        );

    \I__866\ : Odrv12
    port map (
            O => \N__5832\,
            I => \RAMSPACEn_c\
        );

    \I__865\ : InMux
    port map (
            O => \N__5829\,
            I => \N__5826\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__5826\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__863\ : CEMux
    port map (
            O => \N__5823\,
            I => \N__5820\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__5820\,
            I => \N__5817\
        );

    \I__861\ : Odrv4
    port map (
            O => \N__5817\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0\
        );

    \I__860\ : InMux
    port map (
            O => \N__5814\,
            I => \N__5809\
        );

    \I__859\ : CascadeMux
    port map (
            O => \N__5813\,
            I => \N__5804\
        );

    \I__858\ : InMux
    port map (
            O => \N__5812\,
            I => \N__5799\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__5809\,
            I => \N__5796\
        );

    \I__856\ : InMux
    port map (
            O => \N__5808\,
            I => \N__5793\
        );

    \I__855\ : InMux
    port map (
            O => \N__5807\,
            I => \N__5790\
        );

    \I__854\ : InMux
    port map (
            O => \N__5804\,
            I => \N__5783\
        );

    \I__853\ : InMux
    port map (
            O => \N__5803\,
            I => \N__5783\
        );

    \I__852\ : InMux
    port map (
            O => \N__5802\,
            I => \N__5783\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__5799\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__850\ : Odrv4
    port map (
            O => \N__5796\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__5793\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__5790\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__5783\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__846\ : InMux
    port map (
            O => \N__5772\,
            I => \N__5768\
        );

    \I__845\ : InMux
    port map (
            O => \N__5771\,
            I => \N__5764\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__5768\,
            I => \N__5761\
        );

    \I__843\ : InMux
    port map (
            O => \N__5767\,
            I => \N__5758\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__5764\,
            I => \N__5755\
        );

    \I__841\ : Span4Mux_h
    port map (
            O => \N__5761\,
            I => \N__5750\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__5758\,
            I => \N__5750\
        );

    \I__839\ : Span4Mux_v
    port map (
            O => \N__5755\,
            I => \N__5747\
        );

    \I__838\ : Span4Mux_v
    port map (
            O => \N__5750\,
            I => \N__5744\
        );

    \I__837\ : Sp12to4
    port map (
            O => \N__5747\,
            I => \N__5741\
        );

    \I__836\ : Span4Mux_h
    port map (
            O => \N__5744\,
            I => \N__5738\
        );

    \I__835\ : Span12Mux_h
    port map (
            O => \N__5741\,
            I => \N__5733\
        );

    \I__834\ : Sp12to4
    port map (
            O => \N__5738\,
            I => \N__5733\
        );

    \I__833\ : Span12Mux_v
    port map (
            O => \N__5733\,
            I => \N__5730\
        );

    \I__832\ : Odrv12
    port map (
            O => \N__5730\,
            I => \AWEn_c\
        );

    \I__831\ : CascadeMux
    port map (
            O => \N__5727\,
            I => \N__5723\
        );

    \I__830\ : InMux
    port map (
            O => \N__5726\,
            I => \N__5720\
        );

    \I__829\ : InMux
    port map (
            O => \N__5723\,
            I => \N__5716\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__5720\,
            I => \N__5713\
        );

    \I__827\ : InMux
    port map (
            O => \N__5719\,
            I => \N__5710\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__5716\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__825\ : Odrv4
    port map (
            O => \N__5713\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__5710\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__823\ : IoInMux
    port map (
            O => \N__5703\,
            I => \N__5700\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5700\,
            I => \N__5697\
        );

    \I__821\ : IoSpan4Mux
    port map (
            O => \N__5697\,
            I => \N__5694\
        );

    \I__820\ : Sp12to4
    port map (
            O => \N__5694\,
            I => \N__5691\
        );

    \I__819\ : Span12Mux_s9_v
    port map (
            O => \N__5691\,
            I => \N__5687\
        );

    \I__818\ : InMux
    port map (
            O => \N__5690\,
            I => \N__5684\
        );

    \I__817\ : Odrv12
    port map (
            O => \N__5687\,
            I => \DBDIR_c\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__5684\,
            I => \DBDIR_c\
        );

    \I__815\ : IoInMux
    port map (
            O => \N__5679\,
            I => \N__5675\
        );

    \I__814\ : IoInMux
    port map (
            O => \N__5678\,
            I => \N__5672\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5675\,
            I => \N__5668\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5672\,
            I => \N__5665\
        );

    \I__811\ : IoInMux
    port map (
            O => \N__5671\,
            I => \N__5662\
        );

    \I__810\ : Span4Mux_s2_v
    port map (
            O => \N__5668\,
            I => \N__5659\
        );

    \I__809\ : Span12Mux_s2_v
    port map (
            O => \N__5665\,
            I => \N__5656\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__5662\,
            I => \N__5653\
        );

    \I__807\ : Sp12to4
    port map (
            O => \N__5659\,
            I => \N__5650\
        );

    \I__806\ : Span12Mux_h
    port map (
            O => \N__5656\,
            I => \N__5647\
        );

    \I__805\ : Span12Mux_s4_h
    port map (
            O => \N__5653\,
            I => \N__5644\
        );

    \I__804\ : Span12Mux_h
    port map (
            O => \N__5650\,
            I => \N__5641\
        );

    \I__803\ : Span12Mux_v
    port map (
            O => \N__5647\,
            I => \N__5635\
        );

    \I__802\ : Span12Mux_v
    port map (
            O => \N__5644\,
            I => \N__5635\
        );

    \I__801\ : Span12Mux_v
    port map (
            O => \N__5641\,
            I => \N__5632\
        );

    \I__800\ : InMux
    port map (
            O => \N__5640\,
            I => \N__5629\
        );

    \I__799\ : Odrv12
    port map (
            O => \N__5635\,
            I => \TACK_OUTn\
        );

    \I__798\ : Odrv12
    port map (
            O => \N__5632\,
            I => \TACK_OUTn\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5629\,
            I => \TACK_OUTn\
        );

    \I__796\ : InMux
    port map (
            O => \N__5622\,
            I => \N__5619\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__5619\,
            I => \U712_CYCLE_TERM.N_340\
        );

    \I__794\ : IoInMux
    port map (
            O => \N__5616\,
            I => \N__5613\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__5613\,
            I => \N__5609\
        );

    \I__792\ : IoInMux
    port map (
            O => \N__5612\,
            I => \N__5606\
        );

    \I__791\ : Span4Mux_s3_v
    port map (
            O => \N__5609\,
            I => \N__5603\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__5606\,
            I => \N__5599\
        );

    \I__789\ : Span4Mux_v
    port map (
            O => \N__5603\,
            I => \N__5596\
        );

    \I__788\ : IoInMux
    port map (
            O => \N__5602\,
            I => \N__5593\
        );

    \I__787\ : Span4Mux_s2_v
    port map (
            O => \N__5599\,
            I => \N__5590\
        );

    \I__786\ : Span4Mux_h
    port map (
            O => \N__5596\,
            I => \N__5587\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__5593\,
            I => \N__5584\
        );

    \I__784\ : Sp12to4
    port map (
            O => \N__5590\,
            I => \N__5581\
        );

    \I__783\ : Sp12to4
    port map (
            O => \N__5587\,
            I => \N__5578\
        );

    \I__782\ : Span12Mux_s11_h
    port map (
            O => \N__5584\,
            I => \N__5575\
        );

    \I__781\ : Span12Mux_s11_h
    port map (
            O => \N__5581\,
            I => \N__5572\
        );

    \I__780\ : Span12Mux_h
    port map (
            O => \N__5578\,
            I => \N__5568\
        );

    \I__779\ : Span12Mux_v
    port map (
            O => \N__5575\,
            I => \N__5563\
        );

    \I__778\ : Span12Mux_v
    port map (
            O => \N__5572\,
            I => \N__5563\
        );

    \I__777\ : InMux
    port map (
            O => \N__5571\,
            I => \N__5560\
        );

    \I__776\ : Odrv12
    port map (
            O => \N__5568\,
            I => \TACK_EN\
        );

    \I__775\ : Odrv12
    port map (
            O => \N__5563\,
            I => \TACK_EN\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__5560\,
            I => \TACK_EN\
        );

    \I__773\ : CascadeMux
    port map (
            O => \N__5553\,
            I => \U712_CHIP_RAM.N_574_cascade_\
        );

    \I__772\ : InMux
    port map (
            O => \N__5550\,
            I => \N__5543\
        );

    \I__771\ : InMux
    port map (
            O => \N__5549\,
            I => \N__5540\
        );

    \I__770\ : InMux
    port map (
            O => \N__5548\,
            I => \N__5535\
        );

    \I__769\ : InMux
    port map (
            O => \N__5547\,
            I => \N__5535\
        );

    \I__768\ : InMux
    port map (
            O => \N__5546\,
            I => \N__5532\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__5543\,
            I => \N__5529\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__5540\,
            I => \U712_CHIP_RAM.N_475\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__5535\,
            I => \U712_CHIP_RAM.N_475\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5532\,
            I => \U712_CHIP_RAM.N_475\
        );

    \I__763\ : Odrv4
    port map (
            O => \N__5529\,
            I => \U712_CHIP_RAM.N_475\
        );

    \I__762\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5516\
        );

    \I__761\ : InMux
    port map (
            O => \N__5519\,
            I => \N__5513\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__5516\,
            I => \U712_CHIP_RAM.N_328\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__5513\,
            I => \U712_CHIP_RAM.N_328\
        );

    \I__758\ : InMux
    port map (
            O => \N__5508\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__757\ : InMux
    port map (
            O => \N__5505\,
            I => \N__5502\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__5502\,
            I => \N__5499\
        );

    \I__755\ : Odrv4
    port map (
            O => \N__5499\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa\
        );

    \I__754\ : InMux
    port map (
            O => \N__5496\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__753\ : InMux
    port map (
            O => \N__5493\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__752\ : InMux
    port map (
            O => \N__5490\,
            I => \N__5486\
        );

    \I__751\ : InMux
    port map (
            O => \N__5489\,
            I => \N__5483\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__5486\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__5483\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__748\ : InMux
    port map (
            O => \N__5478\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__5475\,
            I => \N__5471\
        );

    \I__746\ : InMux
    port map (
            O => \N__5474\,
            I => \N__5468\
        );

    \I__745\ : InMux
    port map (
            O => \N__5471\,
            I => \N__5465\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__5468\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__5465\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__742\ : InMux
    port map (
            O => \N__5460\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__741\ : InMux
    port map (
            O => \N__5457\,
            I => \N__5453\
        );

    \I__740\ : InMux
    port map (
            O => \N__5456\,
            I => \N__5450\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__5453\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__5450\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__737\ : InMux
    port map (
            O => \N__5445\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__736\ : CascadeMux
    port map (
            O => \N__5442\,
            I => \N__5437\
        );

    \I__735\ : InMux
    port map (
            O => \N__5441\,
            I => \N__5425\
        );

    \I__734\ : InMux
    port map (
            O => \N__5440\,
            I => \N__5425\
        );

    \I__733\ : InMux
    port map (
            O => \N__5437\,
            I => \N__5425\
        );

    \I__732\ : InMux
    port map (
            O => \N__5436\,
            I => \N__5422\
        );

    \I__731\ : InMux
    port map (
            O => \N__5435\,
            I => \N__5413\
        );

    \I__730\ : InMux
    port map (
            O => \N__5434\,
            I => \N__5413\
        );

    \I__729\ : InMux
    port map (
            O => \N__5433\,
            I => \N__5413\
        );

    \I__728\ : InMux
    port map (
            O => \N__5432\,
            I => \N__5413\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__5425\,
            I => \N__5410\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5422\,
            I => \U712_CHIP_RAM.N_47\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__5413\,
            I => \U712_CHIP_RAM.N_47\
        );

    \I__724\ : Odrv4
    port map (
            O => \N__5410\,
            I => \U712_CHIP_RAM.N_47\
        );

    \I__723\ : InMux
    port map (
            O => \N__5403\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__722\ : InMux
    port map (
            O => \N__5400\,
            I => \N__5396\
        );

    \I__721\ : InMux
    port map (
            O => \N__5399\,
            I => \N__5393\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__5396\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__5393\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__718\ : CEMux
    port map (
            O => \N__5388\,
            I => \N__5384\
        );

    \I__717\ : CEMux
    port map (
            O => \N__5387\,
            I => \N__5381\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__5384\,
            I => \N__5378\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__5381\,
            I => \N__5375\
        );

    \I__714\ : Odrv12
    port map (
            O => \N__5378\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__713\ : Odrv12
    port map (
            O => \N__5375\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__712\ : InMux
    port map (
            O => \N__5370\,
            I => \N__5367\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__5367\,
            I => \U712_REG_SM.REGENn_e_1\
        );

    \I__710\ : IoInMux
    port map (
            O => \N__5364\,
            I => \N__5361\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__5361\,
            I => \N__5358\
        );

    \I__708\ : Span4Mux_s1_v
    port map (
            O => \N__5358\,
            I => \N__5355\
        );

    \I__707\ : Sp12to4
    port map (
            O => \N__5355\,
            I => \N__5352\
        );

    \I__706\ : Span12Mux_s7_h
    port map (
            O => \N__5352\,
            I => \N__5349\
        );

    \I__705\ : Span12Mux_v
    port map (
            O => \N__5349\,
            I => \N__5344\
        );

    \I__704\ : InMux
    port map (
            O => \N__5348\,
            I => \N__5341\
        );

    \I__703\ : InMux
    port map (
            O => \N__5347\,
            I => \N__5338\
        );

    \I__702\ : Odrv12
    port map (
            O => \N__5344\,
            I => \REGENn_c\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__5341\,
            I => \REGENn_c\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__5338\,
            I => \REGENn_c\
        );

    \I__699\ : InMux
    port map (
            O => \N__5331\,
            I => \N__5328\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__5328\,
            I => \N__5325\
        );

    \I__697\ : Odrv4
    port map (
            O => \N__5325\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__696\ : InMux
    port map (
            O => \N__5322\,
            I => \N__5318\
        );

    \I__695\ : IoInMux
    port map (
            O => \N__5321\,
            I => \N__5315\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__5318\,
            I => \N__5312\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__5315\,
            I => \N__5309\
        );

    \I__692\ : Span4Mux_v
    port map (
            O => \N__5312\,
            I => \N__5306\
        );

    \I__691\ : IoSpan4Mux
    port map (
            O => \N__5309\,
            I => \N__5303\
        );

    \I__690\ : Sp12to4
    port map (
            O => \N__5306\,
            I => \N__5300\
        );

    \I__689\ : IoSpan4Mux
    port map (
            O => \N__5303\,
            I => \N__5297\
        );

    \I__688\ : Span12Mux_h
    port map (
            O => \N__5300\,
            I => \N__5294\
        );

    \I__687\ : IoSpan4Mux
    port map (
            O => \N__5297\,
            I => \N__5291\
        );

    \I__686\ : Odrv12
    port map (
            O => \N__5294\,
            I => \C1_c\
        );

    \I__685\ : Odrv4
    port map (
            O => \N__5291\,
            I => \C1_c\
        );

    \I__684\ : InMux
    port map (
            O => \N__5286\,
            I => \N__5283\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__5283\,
            I => \N__5280\
        );

    \I__682\ : Odrv4
    port map (
            O => \N__5280\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__681\ : InMux
    port map (
            O => \N__5277\,
            I => \N__5274\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__5274\,
            I => \U712_CHIP_RAM.N_463\
        );

    \I__679\ : CascadeMux
    port map (
            O => \N__5271\,
            I => \N__5268\
        );

    \I__678\ : InMux
    port map (
            O => \N__5268\,
            I => \N__5265\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__5265\,
            I => \U712_CHIP_RAM.N_461\
        );

    \I__676\ : IoInMux
    port map (
            O => \N__5262\,
            I => \N__5259\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__5259\,
            I => \N__5256\
        );

    \I__674\ : Span4Mux_s1_v
    port map (
            O => \N__5256\,
            I => \N__5253\
        );

    \I__673\ : Span4Mux_v
    port map (
            O => \N__5253\,
            I => \N__5250\
        );

    \I__672\ : Span4Mux_v
    port map (
            O => \N__5250\,
            I => \N__5247\
        );

    \I__671\ : Odrv4
    port map (
            O => \N__5247\,
            I => \VBENn_c\
        );

    \I__670\ : InMux
    port map (
            O => \N__5244\,
            I => \N__5241\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__5241\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3\
        );

    \I__668\ : CascadeMux
    port map (
            O => \N__5238\,
            I => \U712_REG_SM.N_337_cascade_\
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__5235\,
            I => \U712_REG_SM.REG_CYCLE_5_iv_0_0_cascade_\
        );

    \I__666\ : InMux
    port map (
            O => \N__5232\,
            I => \N__5229\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__5229\,
            I => \U712_REG_SM.N_424\
        );

    \I__664\ : CascadeMux
    port map (
            O => \N__5226\,
            I => \U712_REG_SM.N_338_cascade_\
        );

    \I__663\ : InMux
    port map (
            O => \N__5223\,
            I => \N__5219\
        );

    \I__662\ : InMux
    port map (
            O => \N__5222\,
            I => \N__5216\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__5219\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_5\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__5216\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_5\
        );

    \I__659\ : InMux
    port map (
            O => \N__5211\,
            I => \N__5208\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__5208\,
            I => \U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1\
        );

    \I__657\ : InMux
    port map (
            O => \N__5205\,
            I => \N__5202\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__5202\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_6\
        );

    \I__655\ : CascadeMux
    port map (
            O => \N__5199\,
            I => \N__5196\
        );

    \I__654\ : InMux
    port map (
            O => \N__5196\,
            I => \N__5193\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__5193\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_7\
        );

    \I__652\ : InMux
    port map (
            O => \N__5190\,
            I => \N__5187\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__5187\,
            I => \N__5183\
        );

    \I__650\ : InMux
    port map (
            O => \N__5186\,
            I => \N__5180\
        );

    \I__649\ : Span4Mux_h
    port map (
            O => \N__5183\,
            I => \N__5177\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__5180\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__647\ : Odrv4
    port map (
            O => \N__5177\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__646\ : InMux
    port map (
            O => \N__5172\,
            I => \N__5169\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__5169\,
            I => \N__5165\
        );

    \I__644\ : InMux
    port map (
            O => \N__5168\,
            I => \N__5162\
        );

    \I__643\ : Span4Mux_h
    port map (
            O => \N__5165\,
            I => \N__5159\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__5162\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__641\ : Odrv4
    port map (
            O => \N__5159\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__640\ : InMux
    port map (
            O => \N__5154\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\
        );

    \I__639\ : InMux
    port map (
            O => \N__5151\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\
        );

    \I__638\ : InMux
    port map (
            O => \N__5148\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\
        );

    \I__637\ : InMux
    port map (
            O => \N__5145\,
            I => \N__5142\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__5142\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\
        );

    \I__635\ : InMux
    port map (
            O => \N__5139\,
            I => \N__5136\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__5136\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\
        );

    \I__633\ : CascadeMux
    port map (
            O => \N__5133\,
            I => \N__5129\
        );

    \I__632\ : InMux
    port map (
            O => \N__5132\,
            I => \N__5126\
        );

    \I__631\ : InMux
    port map (
            O => \N__5129\,
            I => \N__5123\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__5126\,
            I => \DBR_SYNC_i_1\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__5123\,
            I => \DBR_SYNC_i_1\
        );

    \I__628\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5115\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__5115\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a7_0_a2_0\
        );

    \I__626\ : CascadeMux
    port map (
            O => \N__5112\,
            I => \U712_CHIP_RAM.N_475_cascade_\
        );

    \I__625\ : InMux
    port map (
            O => \N__5109\,
            I => \N__5106\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__5106\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0\
        );

    \I__623\ : CascadeMux
    port map (
            O => \N__5103\,
            I => \U712_CHIP_RAM.DBENn_8_0_0_cascade_\
        );

    \I__622\ : InMux
    port map (
            O => \N__5100\,
            I => \N__5096\
        );

    \I__621\ : InMux
    port map (
            O => \N__5099\,
            I => \N__5093\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__5096\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__5093\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__618\ : InMux
    port map (
            O => \N__5088\,
            I => \N__5085\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__5085\,
            I => \N__5082\
        );

    \I__616\ : Span4Mux_v
    port map (
            O => \N__5082\,
            I => \N__5079\
        );

    \I__615\ : Sp12to4
    port map (
            O => \N__5079\,
            I => \N__5076\
        );

    \I__614\ : Span12Mux_h
    port map (
            O => \N__5076\,
            I => \N__5073\
        );

    \I__613\ : Span12Mux_v
    port map (
            O => \N__5073\,
            I => \N__5070\
        );

    \I__612\ : Odrv12
    port map (
            O => \N__5070\,
            I => \A_c_20\
        );

    \I__611\ : InMux
    port map (
            O => \N__5067\,
            I => \N__5060\
        );

    \I__610\ : CascadeMux
    port map (
            O => \N__5066\,
            I => \N__5057\
        );

    \I__609\ : InMux
    port map (
            O => \N__5065\,
            I => \N__5051\
        );

    \I__608\ : InMux
    port map (
            O => \N__5064\,
            I => \N__5051\
        );

    \I__607\ : InMux
    port map (
            O => \N__5063\,
            I => \N__5048\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__5060\,
            I => \N__5045\
        );

    \I__605\ : InMux
    port map (
            O => \N__5057\,
            I => \N__5040\
        );

    \I__604\ : InMux
    port map (
            O => \N__5056\,
            I => \N__5040\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__5051\,
            I => \N__5035\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__5048\,
            I => \N__5035\
        );

    \I__601\ : Odrv4
    port map (
            O => \N__5045\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__5040\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__599\ : Odrv4
    port map (
            O => \N__5035\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__598\ : CascadeMux
    port map (
            O => \N__5028\,
            I => \U712_CYCLE_TERM.N_466_cascade_\
        );

    \I__597\ : CascadeMux
    port map (
            O => \N__5025\,
            I => \U712_CHIP_RAM.N_485_cascade_\
        );

    \I__596\ : InMux
    port map (
            O => \N__5022\,
            I => \N__5019\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__5019\,
            I => \U712_CHIP_RAM.N_325\
        );

    \I__594\ : CascadeMux
    port map (
            O => \N__5016\,
            I => \U712_CHIP_RAM.N_329_cascade_\
        );

    \I__593\ : InMux
    port map (
            O => \N__5013\,
            I => \N__5009\
        );

    \I__592\ : InMux
    port map (
            O => \N__5012\,
            I => \N__5006\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__5009\,
            I => \U712_CHIP_RAM.N_389\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__5006\,
            I => \U712_CHIP_RAM.N_389\
        );

    \I__589\ : InMux
    port map (
            O => \N__5001\,
            I => \N__4995\
        );

    \I__588\ : InMux
    port map (
            O => \N__5000\,
            I => \N__4995\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__4995\,
            I => \N__4991\
        );

    \I__586\ : InMux
    port map (
            O => \N__4994\,
            I => \N__4988\
        );

    \I__585\ : Odrv4
    port map (
            O => \N__4991\,
            I => \U712_CHIP_RAM.N_489\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__4988\,
            I => \U712_CHIP_RAM.N_489\
        );

    \I__583\ : InMux
    port map (
            O => \N__4983\,
            I => \N__4979\
        );

    \I__582\ : InMux
    port map (
            O => \N__4982\,
            I => \N__4976\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__4979\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_a2_1\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__4976\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_a2_1\
        );

    \I__579\ : CascadeMux
    port map (
            O => \N__4971\,
            I => \U712_CHIP_RAM.N_441_cascade_\
        );

    \I__578\ : CascadeMux
    port map (
            O => \N__4968\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_cascade_\
        );

    \I__577\ : CEMux
    port map (
            O => \N__4965\,
            I => \N__4962\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__4962\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0\
        );

    \I__575\ : CascadeMux
    port map (
            O => \N__4959\,
            I => \U712_REG_SM.N_573_cascade_\
        );

    \I__574\ : InMux
    port map (
            O => \N__4956\,
            I => \N__4953\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__4953\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_4\
        );

    \I__572\ : InMux
    port map (
            O => \N__4950\,
            I => \N__4947\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__4947\,
            I => \U712_REG_SM.N_426\
        );

    \I__570\ : InMux
    port map (
            O => \N__4944\,
            I => \N__4939\
        );

    \I__569\ : InMux
    port map (
            O => \N__4943\,
            I => \N__4934\
        );

    \I__568\ : InMux
    port map (
            O => \N__4942\,
            I => \N__4934\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__4939\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_3\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__4934\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_3\
        );

    \I__565\ : CascadeMux
    port map (
            O => \N__4929\,
            I => \U712_CHIP_RAM.N_463_cascade_\
        );

    \I__564\ : CascadeMux
    port map (
            O => \N__4926\,
            I => \N__4923\
        );

    \I__563\ : InMux
    port map (
            O => \N__4923\,
            I => \N__4920\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__4920\,
            I => \U712_REG_SM.N_383\
        );

    \I__561\ : InMux
    port map (
            O => \N__4917\,
            I => \N__4914\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__4914\,
            I => \U712_REG_SM.N_339\
        );

    \I__559\ : CascadeMux
    port map (
            O => \N__4911\,
            I => \U712_REG_SM.N_339_cascade_\
        );

    \I__558\ : InMux
    port map (
            O => \N__4908\,
            I => \N__4905\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__4905\,
            I => \U712_REG_SM.N_350\
        );

    \I__556\ : InMux
    port map (
            O => \N__4902\,
            I => \N__4893\
        );

    \I__555\ : InMux
    port map (
            O => \N__4901\,
            I => \N__4893\
        );

    \I__554\ : InMux
    port map (
            O => \N__4900\,
            I => \N__4893\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__4893\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__552\ : InMux
    port map (
            O => \N__4890\,
            I => \N__4887\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__4887\,
            I => \N__4884\
        );

    \I__550\ : Odrv4
    port map (
            O => \N__4884\,
            I => \U712_REG_SM.N_573\
        );

    \I__549\ : CascadeMux
    port map (
            O => \N__4881\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\
        );

    \I__548\ : InMux
    port map (
            O => \N__4878\,
            I => \N__4875\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4875\,
            I => \N__4872\
        );

    \I__546\ : Sp12to4
    port map (
            O => \N__4872\,
            I => \N__4869\
        );

    \I__545\ : Span12Mux_v
    port map (
            O => \N__4869\,
            I => \N__4866\
        );

    \I__544\ : Odrv12
    port map (
            O => \N__4866\,
            I => \A_c_2\
        );

    \I__543\ : InMux
    port map (
            O => \N__4863\,
            I => \N__4860\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__4860\,
            I => \N__4857\
        );

    \I__541\ : Span4Mux_v
    port map (
            O => \N__4857\,
            I => \N__4854\
        );

    \I__540\ : Span4Mux_v
    port map (
            O => \N__4854\,
            I => \N__4851\
        );

    \I__539\ : Span4Mux_v
    port map (
            O => \N__4851\,
            I => \N__4848\
        );

    \I__538\ : Sp12to4
    port map (
            O => \N__4848\,
            I => \N__4845\
        );

    \I__537\ : Odrv12
    port map (
            O => \N__4845\,
            I => \A_c_3\
        );

    \I__536\ : InMux
    port map (
            O => \N__4842\,
            I => \N__4839\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4839\,
            I => \N__4836\
        );

    \I__534\ : Span4Mux_v
    port map (
            O => \N__4836\,
            I => \N__4833\
        );

    \I__533\ : Span4Mux_v
    port map (
            O => \N__4833\,
            I => \N__4830\
        );

    \I__532\ : Sp12to4
    port map (
            O => \N__4830\,
            I => \N__4827\
        );

    \I__531\ : Odrv12
    port map (
            O => \N__4827\,
            I => \A_c_4\
        );

    \I__530\ : InMux
    port map (
            O => \N__4824\,
            I => \N__4821\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__4821\,
            I => \N__4818\
        );

    \I__528\ : Span4Mux_h
    port map (
            O => \N__4818\,
            I => \N__4815\
        );

    \I__527\ : Span4Mux_v
    port map (
            O => \N__4815\,
            I => \N__4812\
        );

    \I__526\ : Span4Mux_h
    port map (
            O => \N__4812\,
            I => \N__4809\
        );

    \I__525\ : Odrv4
    port map (
            O => \N__4809\,
            I => \A_c_7\
        );

    \I__524\ : InMux
    port map (
            O => \N__4806\,
            I => \N__4803\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4803\,
            I => \N__4800\
        );

    \I__522\ : Sp12to4
    port map (
            O => \N__4800\,
            I => \N__4797\
        );

    \I__521\ : Span12Mux_v
    port map (
            O => \N__4797\,
            I => \N__4794\
        );

    \I__520\ : Odrv12
    port map (
            O => \N__4794\,
            I => \A_c_5\
        );

    \I__519\ : InMux
    port map (
            O => \N__4791\,
            I => \N__4788\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__4788\,
            I => \N__4785\
        );

    \I__517\ : Span4Mux_h
    port map (
            O => \N__4785\,
            I => \N__4782\
        );

    \I__516\ : Span4Mux_v
    port map (
            O => \N__4782\,
            I => \N__4779\
        );

    \I__515\ : Span4Mux_h
    port map (
            O => \N__4779\,
            I => \N__4776\
        );

    \I__514\ : Odrv4
    port map (
            O => \N__4776\,
            I => \A_c_6\
        );

    \I__513\ : InMux
    port map (
            O => \N__4773\,
            I => \N__4770\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__4770\,
            I => \N__4767\
        );

    \I__511\ : Span4Mux_v
    port map (
            O => \N__4767\,
            I => \N__4764\
        );

    \I__510\ : Sp12to4
    port map (
            O => \N__4764\,
            I => \N__4761\
        );

    \I__509\ : Odrv12
    port map (
            O => \N__4761\,
            I => \A_c_8\
        );

    \I__508\ : CEMux
    port map (
            O => \N__4758\,
            I => \N__4754\
        );

    \I__507\ : CEMux
    port map (
            O => \N__4757\,
            I => \N__4751\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__4754\,
            I => \N__4746\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4751\,
            I => \N__4746\
        );

    \I__504\ : Odrv4
    port map (
            O => \N__4746\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\
        );

    \I__503\ : InMux
    port map (
            O => \N__4743\,
            I => \N__4740\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__4740\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__501\ : CascadeMux
    port map (
            O => \N__4737\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_cascade_\
        );

    \I__500\ : IoInMux
    port map (
            O => \N__4734\,
            I => \N__4731\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4731\,
            I => \N__4728\
        );

    \I__498\ : Span4Mux_s3_v
    port map (
            O => \N__4728\,
            I => \N__4725\
        );

    \I__497\ : Span4Mux_h
    port map (
            O => \N__4725\,
            I => \N__4722\
        );

    \I__496\ : Sp12to4
    port map (
            O => \N__4722\,
            I => \N__4719\
        );

    \I__495\ : Span12Mux_v
    port map (
            O => \N__4719\,
            I => \N__4715\
        );

    \I__494\ : InMux
    port map (
            O => \N__4718\,
            I => \N__4712\
        );

    \I__493\ : Odrv12
    port map (
            O => \N__4715\,
            I => \LATCH_CLK_c\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__4712\,
            I => \LATCH_CLK_c\
        );

    \I__491\ : InMux
    port map (
            O => \N__4707\,
            I => \N__4704\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__4704\,
            I => \N__4701\
        );

    \I__489\ : Span4Mux_v
    port map (
            O => \N__4701\,
            I => \N__4698\
        );

    \I__488\ : Span4Mux_v
    port map (
            O => \N__4698\,
            I => \N__4695\
        );

    \I__487\ : Sp12to4
    port map (
            O => \N__4695\,
            I => \N__4692\
        );

    \I__486\ : Odrv12
    port map (
            O => \N__4692\,
            I => \A_c_18\
        );

    \I__485\ : InMux
    port map (
            O => \N__4689\,
            I => \N__4686\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4686\,
            I => \U712_CHIP_RAM.N_462\
        );

    \I__483\ : InMux
    port map (
            O => \N__4683\,
            I => \N__4680\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__4680\,
            I => \U712_CHIP_RAM.N_443\
        );

    \I__481\ : CascadeMux
    port map (
            O => \N__4677\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_1_1_cascade_\
        );

    \I__480\ : InMux
    port map (
            O => \N__4674\,
            I => \N__4671\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4671\,
            I => \N__4668\
        );

    \I__478\ : Odrv4
    port map (
            O => \N__4668\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_1_2\
        );

    \I__477\ : CascadeMux
    port map (
            O => \N__4665\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_1_2_cascade_\
        );

    \I__476\ : CascadeMux
    port map (
            O => \N__4662\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_cascade_\
        );

    \I__475\ : CEMux
    port map (
            O => \N__4659\,
            I => \N__4656\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4656\,
            I => \N__4653\
        );

    \I__473\ : Odrv4
    port map (
            O => \N__4653\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0\
        );

    \I__472\ : InMux
    port map (
            O => \N__4650\,
            I => \N__4647\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__4647\,
            I => \N__4643\
        );

    \I__470\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4640\
        );

    \I__469\ : Span4Mux_h
    port map (
            O => \N__4643\,
            I => \N__4635\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__4640\,
            I => \N__4635\
        );

    \I__467\ : Span4Mux_h
    port map (
            O => \N__4635\,
            I => \N__4632\
        );

    \I__466\ : Sp12to4
    port map (
            O => \N__4632\,
            I => \N__4629\
        );

    \I__465\ : Span12Mux_v
    port map (
            O => \N__4629\,
            I => \N__4626\
        );

    \I__464\ : Odrv12
    port map (
            O => \N__4626\,
            I => \DBRn_c\
        );

    \I__463\ : IoInMux
    port map (
            O => \N__4623\,
            I => \N__4620\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__4620\,
            I => \N__4617\
        );

    \I__461\ : IoSpan4Mux
    port map (
            O => \N__4617\,
            I => \N__4614\
        );

    \I__460\ : Span4Mux_s3_h
    port map (
            O => \N__4614\,
            I => \N__4611\
        );

    \I__459\ : Span4Mux_v
    port map (
            O => \N__4611\,
            I => \N__4607\
        );

    \I__458\ : InMux
    port map (
            O => \N__4610\,
            I => \N__4604\
        );

    \I__457\ : Span4Mux_h
    port map (
            O => \N__4607\,
            I => \N__4601\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__4604\,
            I => \N__4598\
        );

    \I__455\ : Sp12to4
    port map (
            O => \N__4601\,
            I => \N__4595\
        );

    \I__454\ : Span4Mux_v
    port map (
            O => \N__4598\,
            I => \N__4592\
        );

    \I__453\ : Span12Mux_h
    port map (
            O => \N__4595\,
            I => \N__4587\
        );

    \I__452\ : Sp12to4
    port map (
            O => \N__4592\,
            I => \N__4587\
        );

    \I__451\ : Span12Mux_h
    port map (
            O => \N__4587\,
            I => \N__4584\
        );

    \I__450\ : Odrv12
    port map (
            O => \N__4584\,
            I => \C3_c\
        );

    \I__449\ : CascadeMux
    port map (
            O => \N__4581\,
            I => \U712_CHIP_RAM.N_489_cascade_\
        );

    \I__448\ : InMux
    port map (
            O => \N__4578\,
            I => \N__4575\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__4575\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_1\
        );

    \I__446\ : CascadeMux
    port map (
            O => \N__4572\,
            I => \U712_CHIP_RAM.N_413_cascade_\
        );

    \I__445\ : CascadeMux
    port map (
            O => \N__4569\,
            I => \U712_CHIP_RAM.N_159_cascade_\
        );

    \I__444\ : InMux
    port map (
            O => \N__4566\,
            I => \N__4563\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__4563\,
            I => \U712_CHIP_RAM.N_413\
        );

    \I__442\ : InMux
    port map (
            O => \N__4560\,
            I => \N__4556\
        );

    \I__441\ : InMux
    port map (
            O => \N__4559\,
            I => \N__4553\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__4556\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__4553\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__438\ : InMux
    port map (
            O => \N__4548\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__437\ : InMux
    port map (
            O => \N__4545\,
            I => \N__4541\
        );

    \I__436\ : InMux
    port map (
            O => \N__4544\,
            I => \N__4538\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__4541\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__4538\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__433\ : InMux
    port map (
            O => \N__4533\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__432\ : InMux
    port map (
            O => \N__4530\,
            I => \N__4526\
        );

    \I__431\ : InMux
    port map (
            O => \N__4529\,
            I => \N__4523\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__4526\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__4523\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__428\ : InMux
    port map (
            O => \N__4518\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__427\ : CascadeMux
    port map (
            O => \N__4515\,
            I => \N__4511\
        );

    \I__426\ : InMux
    port map (
            O => \N__4514\,
            I => \N__4508\
        );

    \I__425\ : InMux
    port map (
            O => \N__4511\,
            I => \N__4505\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__4508\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__4505\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__422\ : InMux
    port map (
            O => \N__4500\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__421\ : InMux
    port map (
            O => \N__4497\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__420\ : InMux
    port map (
            O => \N__4494\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__419\ : InMux
    port map (
            O => \N__4491\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__418\ : ClkMux
    port map (
            O => \N__4488\,
            I => \N__4467\
        );

    \I__417\ : ClkMux
    port map (
            O => \N__4487\,
            I => \N__4467\
        );

    \I__416\ : ClkMux
    port map (
            O => \N__4486\,
            I => \N__4467\
        );

    \I__415\ : ClkMux
    port map (
            O => \N__4485\,
            I => \N__4467\
        );

    \I__414\ : ClkMux
    port map (
            O => \N__4484\,
            I => \N__4467\
        );

    \I__413\ : ClkMux
    port map (
            O => \N__4483\,
            I => \N__4467\
        );

    \I__412\ : ClkMux
    port map (
            O => \N__4482\,
            I => \N__4467\
        );

    \I__411\ : GlobalMux
    port map (
            O => \N__4467\,
            I => \N__4464\
        );

    \I__410\ : gio2CtrlBuf
    port map (
            O => \N__4464\,
            I => \C1_c_g\
        );

    \I__409\ : IoInMux
    port map (
            O => \N__4461\,
            I => \N__4458\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__4458\,
            I => \N__4455\
        );

    \I__407\ : IoSpan4Mux
    port map (
            O => \N__4455\,
            I => \N__4452\
        );

    \I__406\ : IoSpan4Mux
    port map (
            O => \N__4452\,
            I => \N__4449\
        );

    \I__405\ : Span4Mux_s3_h
    port map (
            O => \N__4449\,
            I => \N__4446\
        );

    \I__404\ : Sp12to4
    port map (
            O => \N__4446\,
            I => \N__4443\
        );

    \I__403\ : Span12Mux_h
    port map (
            O => \N__4443\,
            I => \N__4440\
        );

    \I__402\ : Odrv12
    port map (
            O => \N__4440\,
            I => \CLK_EN_c\
        );

    \I__401\ : InMux
    port map (
            O => \N__4437\,
            I => \N__4434\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__4434\,
            I => \N__4431\
        );

    \I__399\ : Span4Mux_h
    port map (
            O => \N__4431\,
            I => \N__4428\
        );

    \I__398\ : Sp12to4
    port map (
            O => \N__4428\,
            I => \N__4425\
        );

    \I__397\ : Span12Mux_v
    port map (
            O => \N__4425\,
            I => \N__4422\
        );

    \I__396\ : Odrv12
    port map (
            O => \N__4422\,
            I => \REGSPACEn_c\
        );

    \I__395\ : IoInMux
    port map (
            O => \N__4419\,
            I => \N__4416\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__4416\,
            I => \N__4413\
        );

    \I__393\ : Span12Mux_s1_h
    port map (
            O => \N__4413\,
            I => \N__4410\
        );

    \I__392\ : Odrv12
    port map (
            O => \N__4410\,
            I => \DBRn_c_i_0\
        );

    \I__391\ : IoInMux
    port map (
            O => \N__4407\,
            I => \N__4404\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__4404\,
            I => \N__4401\
        );

    \I__389\ : Span4Mux_s2_v
    port map (
            O => \N__4401\,
            I => \N__4398\
        );

    \I__388\ : Span4Mux_v
    port map (
            O => \N__4398\,
            I => \N__4395\
        );

    \I__387\ : Span4Mux_h
    port map (
            O => \N__4395\,
            I => \N__4392\
        );

    \I__386\ : Odrv4
    port map (
            O => \N__4392\,
            I => \CLK80_PLL_i_i\
        );

    \I__385\ : InMux
    port map (
            O => \N__4389\,
            I => \N__4386\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__4386\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__383\ : InMux
    port map (
            O => \N__4383\,
            I => \bfn_6_6_0_\
        );

    \I__382\ : IoInMux
    port map (
            O => \N__4380\,
            I => \N__4377\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__4377\,
            I => \N__4374\
        );

    \I__380\ : IoSpan4Mux
    port map (
            O => \N__4374\,
            I => \N__4371\
        );

    \I__379\ : Span4Mux_s2_v
    port map (
            O => \N__4371\,
            I => \N__4368\
        );

    \I__378\ : Sp12to4
    port map (
            O => \N__4368\,
            I => \N__4365\
        );

    \I__377\ : Span12Mux_v
    port map (
            O => \N__4365\,
            I => \N__4362\
        );

    \I__376\ : Odrv12
    port map (
            O => \N__4362\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            I => \N__4486\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__4487\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__4485\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            I => \N__4482\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            I => \N__4483\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            I => \N__4484\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_6_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_6_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_10_0_\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5321\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__9192\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4419\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4623\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11175\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9878\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10692\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBRn_ibuf_RNIBAB_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4646\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__4529\,
            in1 => \N__4559\,
            in2 => \N__4515\,
            in3 => \N__4544\,
            lcout => \U712_CHIP_RAM.REFRESH5lt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4389\,
            in2 => \_gnd_net_\,
            in3 => \N__4383\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_6_6_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__4488\,
            ce => 'H',
            sr => \N__8130\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4560\,
            in2 => \_gnd_net_\,
            in3 => \N__4548\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__4488\,
            ce => 'H',
            sr => \N__8130\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4545\,
            in2 => \_gnd_net_\,
            in3 => \N__4533\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__4488\,
            ce => 'H',
            sr => \N__8130\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4530\,
            in2 => \_gnd_net_\,
            in3 => \N__4518\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__4488\,
            ce => 'H',
            sr => \N__8130\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4514\,
            in2 => \_gnd_net_\,
            in3 => \N__4500\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__4488\,
            ce => 'H',
            sr => \N__8130\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5168\,
            in2 => \_gnd_net_\,
            in3 => \N__4497\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__4488\,
            ce => 'H',
            sr => \N__8130\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5186\,
            in2 => \_gnd_net_\,
            in3 => \N__4494\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__4488\,
            ce => 'H',
            sr => \N__8130\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5930\,
            in2 => \_gnd_net_\,
            in3 => \N__4491\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4488\,
            ce => 'H',
            sr => \N__8130\
        );

    \U712_CHIP_RAM.CLK_EN_ess_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__7204\,
            in1 => \N__7098\,
            in2 => \_gnd_net_\,
            in3 => \N__7308\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10669\,
            ce => \N__4659\,
            sr => \N__11144\
        );

    \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4437\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5870\,
            lcout => \U712_REG_SM.N_416\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_0_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4650\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10682\,
            ce => 'H',
            sr => \N__11114\
        );

    \U712_REG_SM.C3_SYNC_0_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4610\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10686\,
            ce => 'H',
            sr => \N__11099\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6680\,
            in1 => \N__7206\,
            in2 => \N__7104\,
            in3 => \N__6779\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__7079\,
            in1 => \N__7191\,
            in2 => \_gnd_net_\,
            in3 => \N__7266\,
            lcout => \U712_CHIP_RAM.N_489\,
            ltout => \U712_CHIP_RAM.N_489_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1NGC4_0_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5065\,
            in1 => \N__6681\,
            in2 => \N__4581\,
            in3 => \N__7395\,
            lcout => \U712_CHIP_RAM.N_413\,
            ltout => \U712_CHIP_RAM.N_413_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__7396\,
            in1 => \N__4578\,
            in2 => \N__4572\,
            in3 => \N__4674\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_159_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011111010"
        )
    port map (
            in0 => \N__6169\,
            in1 => \N__4689\,
            in2 => \N__4569\,
            in3 => \N__7080\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10655\,
            ce => 'H',
            sr => \N__11147\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIVFJO_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5064\,
            in2 => \_gnd_net_\,
            in3 => \N__7267\,
            lcout => \U712_CHIP_RAM.N_326\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__7397\,
            in1 => \N__4983\,
            in2 => \_gnd_net_\,
            in3 => \N__4566\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__4718\,
            in1 => \N__7294\,
            in2 => \N__4737\,
            in3 => \N__8404\,
            lcout => \LATCH_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10655\,
            ce => 'H',
            sr => \N__11147\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4707\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10659\,
            ce => \N__4757\,
            sr => \N__11145\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6708\,
            in1 => \N__9599\,
            in2 => \_gnd_net_\,
            in3 => \N__6765\,
            lcout => \U712_CHIP_RAM.N_462\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__9565\,
            in1 => \N__4683\,
            in2 => \_gnd_net_\,
            in3 => \N__5099\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10663\,
            ce => 'H',
            sr => \N__11131\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__7388\,
            in1 => \N__5001\,
            in2 => \N__5066\,
            in3 => \N__6678\,
            lcout => \U712_CHIP_RAM.N_443\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIN93S_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__9564\,
            in1 => \N__5056\,
            in2 => \_gnd_net_\,
            in3 => \N__6675\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIIFS82_3_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__7205\,
            in1 => \N__7097\,
            in2 => \N__4677\,
            in3 => \N__7293\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_1_2\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__5000\,
            in1 => \N__6676\,
            in2 => \N__4665\,
            in3 => \N__7387\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_RNO_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4662\,
            in3 => \N__11172\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIU7TF5_2_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6300\,
            in1 => \N__5892\,
            in2 => \N__7404\,
            in3 => \N__6677\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_1_2_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4881\,
            in3 => \N__11173\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4878\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10670\,
            ce => \N__4758\,
            sr => \N__11127\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4863\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10670\,
            ce => \N__4758\,
            sr => \N__11127\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4842\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10670\,
            ce => \N__4758\,
            sr => \N__11127\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4824\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10670\,
            ce => \N__4758\,
            sr => \N__11127\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4806\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10670\,
            ce => \N__4758\,
            sr => \N__11127\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4791\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10670\,
            ce => \N__4758\,
            sr => \N__11127\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4773\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10670\,
            ce => \N__4758\,
            sr => \N__11127\
        );

    \DBR_SYNC_1_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4743\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10679\,
            ce => 'H',
            sr => \N__11109\
        );

    \U712_REG_SM.REG_TACK_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__4890\,
            in1 => \N__4908\,
            in2 => \N__6217\,
            in3 => \N__5211\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10679\,
            ce => 'H',
            sr => \N__11109\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001010"
        )
    port map (
            in0 => \N__10972\,
            in1 => \N__4917\,
            in2 => \N__4926\,
            in3 => \N__11256\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000110011"
        )
    port map (
            in0 => \N__11254\,
            in1 => \N__4902\,
            in2 => \N__6090\,
            in3 => \N__5958\,
            lcout => \U712_REG_SM.N_383\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIH4AH_1_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6073\,
            in2 => \_gnd_net_\,
            in3 => \N__7534\,
            lcout => \U712_REG_SM.N_339\,
            ltout => \U712_REG_SM.N_339_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_0_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__11255\,
            in1 => \N__4901\,
            in2 => \N__4911\,
            in3 => \N__6464\,
            lcout => \U712_REG_SM.N_424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI3HF31_1_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__5957\,
            in1 => \N__11253\,
            in2 => \N__6465\,
            in3 => \N__6072\,
            lcout => \U712_REG_SM.N_171\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6463\,
            in1 => \N__6005\,
            in2 => \_gnd_net_\,
            in3 => \N__4942\,
            lcout => \U712_REG_SM.N_350\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__4943\,
            in1 => \N__4900\,
            in2 => \N__7548\,
            in3 => \N__6089\,
            lcout => \U712_REG_SM.N_426\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIJUGT_3_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__4944\,
            in1 => \N__11265\,
            in2 => \_gnd_net_\,
            in3 => \N__6077\,
            lcout => \U712_REG_SM.N_573\,
            ltout => \U712_REG_SM.N_573_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4959\,
            in3 => \N__10974\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10975\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4956\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10976\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5223\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011000100"
        )
    port map (
            in0 => \N__6078\,
            in1 => \N__10973\,
            in2 => \N__11285\,
            in3 => \N__4950\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000101110"
        )
    port map (
            in0 => \N__6324\,
            in1 => \N__5436\,
            in2 => \N__5271\,
            in3 => \N__5013\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10648\,
            ce => \N__5387\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_3_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__7163\,
            in1 => \N__7047\,
            in2 => \_gnd_net_\,
            in3 => \N__7258\,
            lcout => \U712_CHIP_RAM.N_480\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI4VIE1_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7171\,
            in1 => \N__8400\,
            in2 => \N__7102\,
            in3 => \N__7263\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6279\,
            in1 => \N__5814\,
            in2 => \N__7398\,
            in3 => \N__6615\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10653\,
            ce => \N__4965\,
            sr => \N__11146\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000000"
        )
    port map (
            in0 => \N__6614\,
            in1 => \N__5546\,
            in2 => \N__6822\,
            in3 => \N__6278\,
            lcout => \U712_CHIP_RAM.N_463\,
            ltout => \U712_CHIP_RAM.N_463_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI0416C_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4929\,
            in3 => \N__5012\,
            lcout => \U712_CHIP_RAM.N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI324S_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6612\,
            in1 => \N__8399\,
            in2 => \_gnd_net_\,
            in3 => \N__6814\,
            lcout => \U712_CHIP_RAM.N_325\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI37LE3_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__7373\,
            in1 => \N__6613\,
            in2 => \N__7289\,
            in3 => \N__5063\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_485_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIDDEL6_0_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__5550\,
            in1 => \N__7262\,
            in2 => \N__5025\,
            in3 => \N__5022\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_329_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI17638_3_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011111111"
        )
    port map (
            in0 => \N__7078\,
            in1 => \N__7170\,
            in2 => \N__5016\,
            in3 => \N__10986\,
            lcout => \U712_CHIP_RAM.N_389\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1NGC4_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5067\,
            in1 => \N__4994\,
            in2 => \N__7405\,
            in3 => \N__6649\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_441_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIMAOKC_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__7386\,
            in1 => \N__4982\,
            in2 => \N__4971\,
            in3 => \N__5719\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__11174\,
            in1 => \_gnd_net_\,
            in2 => \N__4968\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7385\,
            in1 => \N__10985\,
            in2 => \_gnd_net_\,
            in3 => \N__5118\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5808\,
            in1 => \N__6647\,
            in2 => \N__6308\,
            in3 => \N__7384\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6648\,
            in1 => \N__5519\,
            in2 => \_gnd_net_\,
            in3 => \N__6296\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a7_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5456\,
            in1 => \N__5489\,
            in2 => \N__5475\,
            in3 => \N__5399\,
            lcout => \U712_CHIP_RAM.N_475\,
            ltout => \U712_CHIP_RAM.N_475_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5112\,
            in3 => \N__6813\,
            lcout => \U712_CHIP_RAM.N_476\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6301\,
            in1 => \N__6679\,
            in2 => \_gnd_net_\,
            in3 => \N__5549\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.DBENn_8_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010111011101110"
        )
    port map (
            in0 => \N__8449\,
            in1 => \N__5109\,
            in2 => \N__5103\,
            in3 => \N__10386\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10660\,
            ce => 'H',
            sr => \N__11128\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__5100\,
            in1 => \N__5088\,
            in2 => \N__11574\,
            in3 => \N__7796\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10660\,
            ce => 'H',
            sr => \N__11128\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__10533\,
            in1 => \N__5767\,
            in2 => \_gnd_net_\,
            in3 => \N__5812\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10664\,
            ce => \N__5823\,
            sr => \N__11119\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010011"
        )
    port map (
            in0 => \N__6236\,
            in1 => \N__7707\,
            in2 => \N__6219\,
            in3 => \N__6182\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_466_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__7755\,
            in1 => \N__10966\,
            in2 => \N__5028\,
            in3 => \N__6237\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10671\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5190\,
            in2 => \_gnd_net_\,
            in3 => \N__5172\,
            lcout => \U712_CHIP_RAM.REFRESH5lto7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__6181\,
            in1 => \N__6235\,
            in2 => \_gnd_net_\,
            in3 => \N__6213\,
            lcout => \U712_CYCLE_TERM.N_340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7565\,
            in2 => \N__5133\,
            in3 => \N__5132\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7650\,
            in2 => \_gnd_net_\,
            in3 => \N__5154\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7634\,
            in2 => \_gnd_net_\,
            in3 => \N__5151\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7664\,
            in2 => \_gnd_net_\,
            in3 => \N__5148\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_0_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__7538\,
            in1 => \N__5145\,
            in2 => \N__7619\,
            in3 => \N__10959\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10673\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_2_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__7525\,
            in1 => \N__7613\,
            in2 => \N__10987\,
            in3 => \N__5139\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10673\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_RNITKK4_1_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7524\,
            lcout => \DBR_SYNC_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_3_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__7526\,
            in1 => \N__7614\,
            in2 => \N__10988\,
            in3 => \N__5244\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10673\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11284\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6093\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_337_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__10807\,
            in1 => \N__5982\,
            in2 => \N__5238\,
            in3 => \N__5963\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_1_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__6457\,
            in1 => \N__8050\,
            in2 => \N__6006\,
            in3 => \N__6415\,
            lcout => OPEN,
            ltout => \U712_REG_SM.REG_CYCLE_5_iv_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__8051\,
            in1 => \N__10967\,
            in2 => \N__5235\,
            in3 => \N__5232\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11269\,
            in2 => \_gnd_net_\,
            in3 => \N__6087\,
            lcout => \U712_REG_SM.N_338\,
            ltout => \U712_REG_SM.N_338_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__6456\,
            in1 => \N__6400\,
            in2 => \N__5226\,
            in3 => \N__5222\,
            lcout => \U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_8_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__6416\,
            in1 => \N__10969\,
            in2 => \N__5199\,
            in3 => \N__6458\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_7_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10968\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5205\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_RNO_0_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001100010"
        )
    port map (
            in0 => \N__6088\,
            in1 => \N__5347\,
            in2 => \N__5967\,
            in3 => \N__6024\,
            lcout => \U712_REG_SM.REGENn_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010011010100010"
        )
    port map (
            in0 => \N__5348\,
            in1 => \N__5370\,
            in2 => \N__11292\,
            in3 => \N__6401\,
            lcout => \REGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10684\,
            ce => 'H',
            sr => \N__11094\
        );

    \U712_REG_SM.C1_SYNC_1_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5286\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10684\,
            ce => 'H',
            sr => \N__11094\
        );

    \U712_REG_SM.C3_SYNC_1_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5331\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10684\,
            ce => 'H',
            sr => \N__11094\
        );

    \U712_REG_SM.C1_SYNC_0_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5322\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10687\,
            ce => 'H',
            sr => \N__11092\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__5277\,
            in1 => \_gnd_net_\,
            in2 => \N__6672\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_461\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000011000"
        )
    port map (
            in0 => \N__7264\,
            in1 => \N__6632\,
            in2 => \N__7090\,
            in3 => \N__7172\,
            lcout => \U712_CHIP_RAM.N_320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_0_a2_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__8070\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9664\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_0_2_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6510\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7265\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7173\,
            lcout => \U712_CHIP_RAM.N_477\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7288\,
            in2 => \_gnd_net_\,
            in3 => \N__6724\,
            lcout => \U712_CHIP_RAM.N_411\,
            ltout => OPEN,
            carryin => \bfn_9_5_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5432\,
            in1 => \N__7077\,
            in2 => \_gnd_net_\,
            in3 => \N__5508\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__10649\,
            ce => \N__5388\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__5505\,
            in1 => \N__6671\,
            in2 => \N__5442\,
            in3 => \N__5496\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \N__10649\,
            ce => \N__5388\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5433\,
            in1 => \N__7190\,
            in2 => \_gnd_net_\,
            in3 => \N__5493\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__10649\,
            ce => \N__5388\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5440\,
            in1 => \N__5490\,
            in2 => \_gnd_net_\,
            in3 => \N__5478\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__10649\,
            ce => \N__5388\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5434\,
            in1 => \N__5474\,
            in2 => \_gnd_net_\,
            in3 => \N__5460\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__10649\,
            ce => \N__5388\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5441\,
            in1 => \N__5457\,
            in2 => \_gnd_net_\,
            in3 => \N__5445\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__10649\,
            ce => \N__5388\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5435\,
            in1 => \N__5400\,
            in2 => \_gnd_net_\,
            in3 => \N__5403\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10649\,
            ce => \N__5388\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_1_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6306\,
            in1 => \N__5520\,
            in2 => \N__6673\,
            in3 => \N__7378\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__10979\,
            in1 => \N__6750\,
            in2 => \_gnd_net_\,
            in3 => \N__6821\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10654\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_2_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6307\,
            in1 => \N__10981\,
            in2 => \N__6674\,
            in3 => \N__7380\,
            lcout => \U712_CHIP_RAM.N_447\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_2_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5548\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6640\,
            lcout => \U712_CHIP_RAM.N_572\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNI81M63_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__5807\,
            in1 => \N__10978\,
            in2 => \_gnd_net_\,
            in3 => \N__7377\,
            lcout => \U712_CHIP_RAM.N_574\,
            ltout => \U712_CHIP_RAM.N_574_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_2_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5883\,
            in1 => \N__6305\,
            in2 => \N__5553\,
            in3 => \N__6636\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10980\,
            in2 => \_gnd_net_\,
            in3 => \N__5547\,
            lcout => \U712_CHIP_RAM.N_555\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_1_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7379\,
            in1 => \N__7075\,
            in2 => \N__10989\,
            in3 => \N__6644\,
            lcout => \U712_CHIP_RAM.N_566\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__6901\,
            in1 => \N__6988\,
            in2 => \N__6963\,
            in3 => \N__5802\,
            lcout => \U712_CHIP_RAM.N_328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101000100000"
        )
    port map (
            in0 => \N__10939\,
            in1 => \N__5772\,
            in2 => \N__5727\,
            in3 => \N__11806\,
            lcout => \DMA_WRITE_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10656\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001100"
        )
    port map (
            in0 => \N__5934\,
            in1 => \N__10940\,
            in2 => \N__5916\,
            in3 => \N__5904\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10656\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_0_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5803\,
            in1 => \N__6989\,
            in2 => \N__6962\,
            in3 => \N__6903\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__6902\,
            in1 => \N__6954\,
            in2 => \_gnd_net_\,
            in3 => \N__6987\,
            lcout => \U712_CHIP_RAM.N_327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000010000"
        )
    port map (
            in0 => \N__5877\,
            in1 => \N__5847\,
            in2 => \N__10977\,
            in3 => \N__6936\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10656\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11171\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5829\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010101000"
        )
    port map (
            in0 => \N__10938\,
            in1 => \N__7782\,
            in2 => \N__5813\,
            in3 => \N__8412\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10656\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBDIR_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__5771\,
            in1 => \N__5726\,
            in2 => \_gnd_net_\,
            in3 => \N__5690\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10661\,
            ce => 'H',
            sr => \N__11115\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110100010"
        )
    port map (
            in0 => \N__5640\,
            in1 => \N__7714\,
            in2 => \N__7765\,
            in3 => \N__7680\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10665\,
            ce => 'H',
            sr => \N__11110\
        );

    \U712_CYCLE_TERM.TACK_EN_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011111111"
        )
    port map (
            in0 => \N__6836\,
            in1 => \N__5571\,
            in2 => \_gnd_net_\,
            in3 => \N__5622\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10665\,
            ce => 'H',
            sr => \N__11110\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000111000001100"
        )
    port map (
            in0 => \N__6828\,
            in1 => \N__6837\,
            in2 => \N__7719\,
            in3 => \N__6147\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10665\,
            ce => 'H',
            sr => \N__11110\
        );

    \U712_CHIP_RAM.CAS_COUNTER_1_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__7550\,
            in1 => \N__10958\,
            in2 => \N__7618\,
            in3 => \N__6225\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6218\,
            in2 => \_gnd_net_\,
            in3 => \N__6183\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6021\,
            in1 => \N__6092\,
            in2 => \N__6402\,
            in3 => \N__11283\,
            lcout => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_RNI8MQ3_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7767\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011001100"
        )
    port map (
            in0 => \N__6091\,
            in1 => \N__6396\,
            in2 => \N__11293\,
            in3 => \N__6022\,
            lcout => \U712_REG_SM.STATE_COUNTsr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011100000"
        )
    port map (
            in0 => \N__6023\,
            in1 => \N__6036\,
            in2 => \N__10846\,
            in3 => \N__6477\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10674\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.WRITE_CYCLE_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__10528\,
            in1 => \N__5980\,
            in2 => \_gnd_net_\,
            in3 => \N__6004\,
            lcout => \U712_REG_SM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10677\,
            ce => 'H',
            sr => \N__11095\
        );

    \U712_REG_SM.START_RST_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__6476\,
            in1 => \N__5981\,
            in2 => \_gnd_net_\,
            in3 => \N__5962\,
            lcout => \U712_REG_SM.START_RSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10677\,
            ce => 'H',
            sr => \N__11095\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__6459\,
            in1 => \N__6426\,
            in2 => \_gnd_net_\,
            in3 => \N__6417\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10677\,
            ce => 'H',
            sr => \N__11095\
        );

    \U712_REG_SM.UDSn_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__6348\,
            in1 => \N__11693\,
            in2 => \N__6365\,
            in3 => \N__11279\,
            lcout => \UDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10677\,
            ce => 'H',
            sr => \N__11095\
        );

    \U712_REG_SM.UDSn_RNO_0_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__8944\,
            in1 => \N__9144\,
            in2 => \N__8877\,
            in3 => \N__10508\,
            lcout => \U712_REG_SM.N_435\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_10_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__6335\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7301\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOV791_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7070\,
            in1 => \N__6645\,
            in2 => \_gnd_net_\,
            in3 => \N__6818\,
            lcout => \U712_CHIP_RAM.N_349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6819\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6315\,
            lcout => \U712_CHIP_RAM.N_571\,
            ltout => \U712_CHIP_RAM.N_571_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIF4EE6_2_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101000"
        )
    port map (
            in0 => \N__6543\,
            in1 => \N__6309\,
            in2 => \N__6240\,
            in3 => \N__6646\,
            lcout => \U712_CHIP_RAM.N_410\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__6650\,
            in1 => \N__6820\,
            in2 => \_gnd_net_\,
            in3 => \N__6697\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_i_a2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__6783\,
            in1 => \N__6542\,
            in2 => \N__6768\,
            in3 => \N__6725\,
            lcout => \U712_CHIP_RAM.N_151\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7071\,
            in1 => \N__7307\,
            in2 => \N__7203\,
            in3 => \N__6761\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__6969\,
            in1 => \N__6744\,
            in2 => \N__6738\,
            in3 => \N__6541\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_i_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110100000001"
        )
    port map (
            in0 => \N__6495\,
            in1 => \N__7899\,
            in2 => \N__6729\,
            in3 => \N__8763\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6704\,
            in1 => \N__10970\,
            in2 => \N__7413\,
            in3 => \N__6651\,
            lcout => \U712_CHIP_RAM.N_408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_3_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6540\,
            in1 => \N__7306\,
            in2 => \N__7202\,
            in3 => \N__6525\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_444_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNINN3QI_2_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6519\,
            in1 => \N__7314\,
            in2 => \N__6513\,
            in3 => \N__6506\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000001"
        )
    port map (
            in0 => \N__6494\,
            in1 => \N__6486\,
            in2 => \N__6480\,
            in3 => \N__9833\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIPORK3_3_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7183\,
            in1 => \N__10971\,
            in2 => \N__7412\,
            in3 => \N__7076\,
            lcout => \U712_CHIP_RAM.N_446\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__7305\,
            in1 => \N__7201\,
            in2 => \N__7103\,
            in3 => \N__6990\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_i_i_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6961\,
            in2 => \_gnd_net_\,
            in3 => \N__9606\,
            lcout => \U712_CHIP_RAM.N_431\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6930\,
            in1 => \N__6912\,
            in2 => \_gnd_net_\,
            in3 => \N__8652\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000100010"
        )
    port map (
            in0 => \N__10917\,
            in1 => \N__7497\,
            in2 => \N__7620\,
            in3 => \N__7551\,
            lcout => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8653\,
            in1 => \N__6881\,
            in2 => \_gnd_net_\,
            in3 => \N__6846\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10916\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7679\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10662\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7678\,
            in2 => \_gnd_net_\,
            in3 => \N__7688\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__7773\,
            in1 => \N__8096\,
            in2 => \_gnd_net_\,
            in3 => \N__7596\,
            lcout => \U712_CHIP_RAM.N_471\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_5_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__8097\,
            in1 => \N__10913\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10662\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__10914\,
            in1 => \N__7766\,
            in2 => \_gnd_net_\,
            in3 => \N__7715\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10662\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__7689\,
            in1 => \N__10915\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10662\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10911\,
            in2 => \_gnd_net_\,
            in3 => \N__8013\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__7665\,
            in1 => \N__7649\,
            in2 => \N__7638\,
            in3 => \N__7595\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7569\,
            in2 => \N__7554\,
            in3 => \N__7549\,
            lcout => \U712_CHIP_RAM.N_433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__7466\,
            in1 => \N__11694\,
            in2 => \N__11298\,
            in3 => \N__8007\,
            lcout => \LDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10675\,
            ce => 'H',
            sr => \N__11093\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7454\,
            in1 => \N__7425\,
            in2 => \_gnd_net_\,
            in3 => \N__8619\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9635\,
            in1 => \N__7968\,
            in2 => \N__8664\,
            in3 => \N__9912\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__9333\,
            in1 => \N__9387\,
            in2 => \N__7959\,
            in3 => \N__9783\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10640\,
            ce => \N__9262\,
            sr => \N__11120\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9824\,
            in1 => \N__11666\,
            in2 => \N__8769\,
            in3 => \N__8608\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8609\,
            in1 => \N__7944\,
            in2 => \_gnd_net_\,
            in3 => \N__7923\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001101"
        )
    port map (
            in0 => \N__7898\,
            in1 => \N__8610\,
            in2 => \N__7914\,
            in3 => \N__7905\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10643\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__7897\,
            in1 => \N__7884\,
            in2 => \_gnd_net_\,
            in3 => \N__11667\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10643\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7868\,
            in1 => \N__7836\,
            in2 => \_gnd_net_\,
            in3 => \N__8616\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8618\,
            in1 => \N__9651\,
            in2 => \N__7824\,
            in3 => \N__9234\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7815\,
            in1 => \N__7797\,
            in2 => \_gnd_net_\,
            in3 => \N__8617\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8106\,
            in1 => \N__9633\,
            in2 => \_gnd_net_\,
            in3 => \N__9900\,
            lcout => \U712_CHIP_RAM.N_374\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_4_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10912\,
            in2 => \_gnd_net_\,
            in3 => \N__9210\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10658\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_217_i_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000101"
        )
    port map (
            in0 => \N__8355\,
            in1 => \N__11788\,
            in2 => \N__8430\,
            in3 => \N__8476\,
            lcout => \N_217_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.N_182_i_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100000"
        )
    port map (
            in0 => \N__10459\,
            in1 => \N__8063\,
            in2 => \N__11789\,
            in3 => \N__9634\,
            lcout => \N_182_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_i_x2_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__8876\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9149\,
            lcout => \U712_BYTE_ENABLE.N_315_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__11772\,
            in1 => \N__10790\,
            in2 => \_gnd_net_\,
            in3 => \N__10424\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10667\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_RNO_0_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__10515\,
            in1 => \N__8969\,
            in2 => \N__9148\,
            in3 => \N__8853\,
            lcout => \U712_REG_SM.N_434\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.N_198_i_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__11771\,
            in1 => \N__10442\,
            in2 => \_gnd_net_\,
            in3 => \N__11831\,
            lcout => \N_198_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_343_i_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010110000"
        )
    port map (
            in0 => \N__9052\,
            in1 => \N__8976\,
            in2 => \N__8871\,
            in3 => \N__9135\,
            lcout => \N_343_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CASn_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8663\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10637\,
            ce => 'H',
            sr => \N__11126\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9671\,
            in1 => \N__8220\,
            in2 => \N__8667\,
            in3 => \N__10233\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__9374\,
            in1 => \N__8295\,
            in2 => \N__8665\,
            in3 => \N__8214\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10638\,
            ce => \N__9260\,
            sr => \N__11113\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__9373\,
            in1 => \N__8777\,
            in2 => \_gnd_net_\,
            in3 => \N__8651\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10638\,
            ce => \N__9260\,
            sr => \N__11113\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8112\,
            in2 => \N__8139\,
            in3 => \N__8286\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10638\,
            ce => \N__9260\,
            sr => \N__11113\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8642\,
            in1 => \N__9669\,
            in2 => \N__8148\,
            in3 => \N__10221\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__9838\,
            in1 => \N__8770\,
            in2 => \N__8659\,
            in3 => \N__8129\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_CMA25_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__11170\,
            in1 => \_gnd_net_\,
            in2 => \N__8115\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_CMA25_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011111111"
        )
    port map (
            in0 => \N__11706\,
            in1 => \N__9372\,
            in2 => \N__9680\,
            in3 => \N__8644\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8316\,
            in1 => \N__9665\,
            in2 => \_gnd_net_\,
            in3 => \N__10245\,
            lcout => \U712_CHIP_RAM.N_368\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9837\,
            in2 => \_gnd_net_\,
            in3 => \N__11668\,
            lcout => \U712_CHIP_RAM.N_330\,
            ltout => \U712_CHIP_RAM.N_330_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100000101"
        )
    port map (
            in0 => \N__8643\,
            in1 => \N__9670\,
            in2 => \N__8289\,
            in3 => \N__11705\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__9839\,
            in1 => \N__8641\,
            in2 => \_gnd_net_\,
            in3 => \N__11669\,
            lcout => \U712_CHIP_RAM.CMA_5_i_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9630\,
            in1 => \N__8280\,
            in2 => \N__8666\,
            in3 => \N__9720\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__8630\,
            in1 => \N__8274\,
            in2 => \N__9861\,
            in3 => \N__9631\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8268\,
            in1 => \N__8253\,
            in2 => \_gnd_net_\,
            in3 => \N__8629\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8631\,
            in1 => \N__9632\,
            in2 => \N__8238\,
            in3 => \N__9216\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNI8NM9_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9629\,
            in2 => \_gnd_net_\,
            in3 => \N__8628\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8694\,
            in1 => \N__8685\,
            in2 => \_gnd_net_\,
            in3 => \N__8654\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8655\,
            in1 => \N__9675\,
            in2 => \N__8526\,
            in3 => \N__9222\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_a2_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000000"
        )
    port map (
            in0 => \N__8348\,
            in1 => \N__9051\,
            in2 => \N__8980\,
            in3 => \N__9676\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_454_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_215_i_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001101"
        )
    port map (
            in0 => \N__8425\,
            in1 => \N__10461\,
            in2 => \N__8523\,
            in3 => \N__8475\,
            lcout => \N_215_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_213_i_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__8474\,
            in1 => \N__8322\,
            in2 => \N__11790\,
            in3 => \N__8424\,
            lcout => \N_213_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011100000000"
        )
    port map (
            in0 => \N__8347\,
            in1 => \N__8982\,
            in2 => \N__9054\,
            in3 => \N__9679\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_450_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_211_i_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__8477\,
            in1 => \N__10460\,
            in2 => \N__8433\,
            in3 => \N__8429\,
            lcout => \N_211_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100000000"
        )
    port map (
            in0 => \N__9044\,
            in1 => \N__9203\,
            in2 => \N__8349\,
            in3 => \N__9677\,
            lcout => \U712_BYTE_ENABLE.N_456\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000000"
        )
    port map (
            in0 => \N__8346\,
            in1 => \N__9204\,
            in2 => \N__9053\,
            in3 => \N__9678\,
            lcout => \U712_BYTE_ENABLE.N_452\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_3_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10873\,
            in2 => \_gnd_net_\,
            in3 => \N__11310\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_6_i_o2_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9153\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8981\,
            lcout => \N_322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10890\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_342_i_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100100010"
        )
    port map (
            in0 => \N__9152\,
            in1 => \N__9020\,
            in2 => \N__8973\,
            in3 => \N__8872\,
            lcout => \N_342_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_345_i_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010010101000"
        )
    port map (
            in0 => \N__9151\,
            in1 => \N__9043\,
            in2 => \N__8975\,
            in3 => \N__8861\,
            lcout => \N_345_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_344_i_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000110100010"
        )
    port map (
            in0 => \N__9150\,
            in1 => \N__9042\,
            in2 => \N__8974\,
            in3 => \N__8860\,
            lcout => \N_344_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CRCSn_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8781\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10639\,
            ce => 'H',
            sr => \N__11129\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__9332\,
            in1 => \N__10344\,
            in2 => \N__9388\,
            in3 => \N__8718\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10641\,
            ce => \N__9263\,
            sr => \N__11121\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__9708\,
            in1 => \N__9702\,
            in2 => \N__9681\,
            in3 => \N__11388\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10644\,
            ce => \N__9261\,
            sr => \N__11116\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__9321\,
            in1 => \N__10041\,
            in2 => \N__9389\,
            in3 => \N__9507\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10651\,
            ce => \N__9264\,
            sr => \N__11111\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010010000000"
        )
    port map (
            in0 => \N__9323\,
            in1 => \N__9385\,
            in2 => \N__10332\,
            in3 => \N__9480\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10651\,
            ce => \N__9264\,
            sr => \N__11111\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__9322\,
            in1 => \N__9771\,
            in2 => \N__9390\,
            in3 => \N__9453\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10651\,
            ce => \N__9264\,
            sr => \N__11111\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__9324\,
            in1 => \N__9386\,
            in2 => \N__9420\,
            in3 => \N__9726\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10651\,
            ce => \N__9264\,
            sr => \N__11111\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__9384\,
            in1 => \N__9325\,
            in2 => \N__9294\,
            in3 => \N__10167\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10651\,
            ce => \N__9264\,
            sr => \N__11111\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__9763\,
            in1 => \_gnd_net_\,
            in2 => \N__11565\,
            in3 => \N__10209\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__11341\,
            sr => \N__11100\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11546\,
            in1 => \N__10277\,
            in2 => \_gnd_net_\,
            in3 => \N__10107\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__11341\,
            sr => \N__11100\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__10317\,
            in1 => \_gnd_net_\,
            in2 => \N__10281\,
            in3 => \N__11547\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__11341\,
            sr => \N__11100\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10105\,
            in1 => \N__11544\,
            in2 => \_gnd_net_\,
            in3 => \N__10150\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__11339\,
            sr => \N__11097\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11545\,
            in1 => \N__9762\,
            in2 => \_gnd_net_\,
            in3 => \N__10316\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__11339\,
            sr => \N__11097\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__11617\,
            in1 => \N__11504\,
            in2 => \N__9888\,
            in3 => \N__9857\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            ce => 'H',
            sr => \N__11096\
        );

    \U712_CHIP_RAM.RASn_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9843\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10642\,
            ce => 'H',
            sr => \N__11132\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10021\,
            in1 => \N__11551\,
            in2 => \_gnd_net_\,
            in3 => \N__10143\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11373\,
            ce => \N__11344\,
            sr => \N__11117\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9764\,
            in1 => \N__11552\,
            in2 => \_gnd_net_\,
            in3 => \N__10315\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11373\,
            ce => \N__11344\,
            sr => \N__11117\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__10208\,
            in1 => \_gnd_net_\,
            in2 => \N__11566\,
            in3 => \N__9765\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11373\,
            ce => \N__11344\,
            sr => \N__11117\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11543\,
            in1 => \N__11625\,
            in2 => \_gnd_net_\,
            in3 => \N__10207\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__11343\,
            sr => \N__11112\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9964\,
            in1 => \N__11542\,
            in2 => \_gnd_net_\,
            in3 => \N__10371\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__11343\,
            sr => \N__11112\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10370\,
            in1 => \N__11477\,
            in2 => \_gnd_net_\,
            in3 => \N__9948\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11370\,
            ce => \N__11342\,
            sr => \N__11101\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11541\,
            in1 => \N__10271\,
            in2 => \_gnd_net_\,
            in3 => \N__10106\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11370\,
            ce => \N__11342\,
            sr => \N__11101\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10308\,
            in1 => \N__11476\,
            in2 => \_gnd_net_\,
            in3 => \N__10270\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11369\,
            ce => \N__11340\,
            sr => \N__11098\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10029\,
            in1 => \N__11567\,
            in2 => \_gnd_net_\,
            in3 => \N__9966\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__11347\,
            sr => \N__11130\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10155\,
            in1 => \N__11557\,
            in2 => \_gnd_net_\,
            in3 => \N__10020\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__11346\,
            sr => \N__11122\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__10206\,
            in1 => \_gnd_net_\,
            in2 => \N__11564\,
            in3 => \N__11624\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11371\,
            ce => \N__11345\,
            sr => \N__11118\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10151\,
            in1 => \N__10095\,
            in2 => \_gnd_net_\,
            in3 => \N__11537\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11371\,
            ce => \N__11345\,
            sr => \N__11118\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11556\,
            in1 => \N__10028\,
            in2 => \_gnd_net_\,
            in3 => \N__9965\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11372\,
            ce => \N__11348\,
            sr => \N__11133\
        );

    \U712_REG_SM.ASn_ess_RNO_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11169\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11692\,
            lcout => \U712_REG_SM.N_171_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WEn_LC_18_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11673\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10668\,
            ce => 'H',
            sr => \N__11148\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__11603\,
            in1 => \N__10712\,
            in2 => \_gnd_net_\,
            in3 => \N__11527\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11368\,
            ce => \N__11349\,
            sr => \N__11134\
        );

    \U712_CHIP_RAM.RAS_SYNC_2_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10810\,
            in2 => \_gnd_net_\,
            in3 => \N__10995\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11294\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10688\,
            ce => \N__11181\,
            sr => \N__11102\
        );

    \U712_CHIP_RAM.RAS_SYNC_1_LC_19_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10809\,
            in2 => \_gnd_net_\,
            in3 => \N__10698\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10681\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_0_LC_19_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__10808\,
            in1 => \N__10731\,
            in2 => \_gnd_net_\,
            in3 => \N__10719\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10681\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011100001111"
        )
    port map (
            in0 => \N__10532\,
            in1 => \N__10420\,
            in2 => \N__11832\,
            in3 => \N__11746\,
            lcout => \N_385\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 12 2025 19:38:10

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U111_TOP" view "INTERFACE"

module U111_TOP (
    D_UU_AMIGA,
    D_LL_AMIGA,
    D_UM_AMIGA,
    D_LM_AMIGA,
    D_UU_040,
    D_LM_040,
    D_UM_040,
    D_LL_040,
    A_AMIGA,
    A_040,
    SIZ,
    TEAn,
    TSn,
    RESETn,
    CLKRAMA,
    PORTSIZE,
    TEA_CPUn,
    LBENn,
    CLK40B,
    TBI_CPUn,
    TAn,
    CPUBGn,
    BUFENn,
    RnW,
    CLK80_CPU,
    BUFDIR,
    TCI_CPUn,
    TS_CPUn,
    CLKRAMB,
    CLK40A,
    TCIn,
    TBIn,
    DMAn,
    CLK40C,
    CLK40_IN,
    TACKn,
    BGn);

    inout [7:0] D_UU_AMIGA;
    inout [7:0] D_LL_AMIGA;
    inout [7:0] D_UM_AMIGA;
    inout [7:0] D_LM_AMIGA;
    inout [7:0] D_UU_040;
    inout [7:0] D_LM_040;
    inout [7:0] D_UM_040;
    inout [7:0] D_LL_040;
    output [1:0] A_AMIGA;
    input [1:0] A_040;
    input [1:0] SIZ;
    input TEAn;
    output TSn;
    input RESETn;
    output CLKRAMA;
    input PORTSIZE;
    output TEA_CPUn;
    input LBENn;
    output CLK40B;
    output TBI_CPUn;
    inout TAn;
    output CPUBGn;
    output BUFENn;
    input RnW;
    output CLK80_CPU;
    output BUFDIR;
    output TCI_CPUn;
    input TS_CPUn;
    output CLKRAMB;
    output CLK40A;
    input TCIn;
    input TBIn;
    output DMAn;
    output CLK40C;
    input CLK40_IN;
    inout TACKn;
    input BGn;

    wire N__12664;
    wire N__12648;
    wire N__12647;
    wire N__12646;
    wire N__12639;
    wire N__12638;
    wire N__12637;
    wire N__12630;
    wire N__12629;
    wire N__12628;
    wire N__12621;
    wire N__12620;
    wire N__12619;
    wire N__12612;
    wire N__12611;
    wire N__12610;
    wire N__12603;
    wire N__12602;
    wire N__12601;
    wire N__12594;
    wire N__12593;
    wire N__12592;
    wire N__12585;
    wire N__12584;
    wire N__12583;
    wire N__12576;
    wire N__12575;
    wire N__12574;
    wire N__12567;
    wire N__12566;
    wire N__12565;
    wire N__12558;
    wire N__12557;
    wire N__12556;
    wire N__12549;
    wire N__12548;
    wire N__12547;
    wire N__12540;
    wire N__12539;
    wire N__12538;
    wire N__12531;
    wire N__12530;
    wire N__12529;
    wire N__12522;
    wire N__12521;
    wire N__12520;
    wire N__12513;
    wire N__12512;
    wire N__12511;
    wire N__12504;
    wire N__12503;
    wire N__12502;
    wire N__12495;
    wire N__12494;
    wire N__12493;
    wire N__12486;
    wire N__12485;
    wire N__12484;
    wire N__12477;
    wire N__12476;
    wire N__12475;
    wire N__12468;
    wire N__12467;
    wire N__12466;
    wire N__12459;
    wire N__12458;
    wire N__12457;
    wire N__12450;
    wire N__12449;
    wire N__12448;
    wire N__12441;
    wire N__12440;
    wire N__12439;
    wire N__12432;
    wire N__12431;
    wire N__12430;
    wire N__12423;
    wire N__12422;
    wire N__12421;
    wire N__12414;
    wire N__12413;
    wire N__12412;
    wire N__12405;
    wire N__12404;
    wire N__12403;
    wire N__12396;
    wire N__12395;
    wire N__12394;
    wire N__12387;
    wire N__12386;
    wire N__12385;
    wire N__12378;
    wire N__12377;
    wire N__12376;
    wire N__12369;
    wire N__12368;
    wire N__12367;
    wire N__12360;
    wire N__12359;
    wire N__12358;
    wire N__12351;
    wire N__12350;
    wire N__12349;
    wire N__12342;
    wire N__12341;
    wire N__12340;
    wire N__12333;
    wire N__12332;
    wire N__12331;
    wire N__12324;
    wire N__12323;
    wire N__12322;
    wire N__12315;
    wire N__12314;
    wire N__12313;
    wire N__12306;
    wire N__12305;
    wire N__12304;
    wire N__12297;
    wire N__12296;
    wire N__12295;
    wire N__12288;
    wire N__12287;
    wire N__12286;
    wire N__12279;
    wire N__12278;
    wire N__12277;
    wire N__12270;
    wire N__12269;
    wire N__12268;
    wire N__12261;
    wire N__12260;
    wire N__12259;
    wire N__12252;
    wire N__12251;
    wire N__12250;
    wire N__12243;
    wire N__12242;
    wire N__12241;
    wire N__12234;
    wire N__12233;
    wire N__12232;
    wire N__12225;
    wire N__12224;
    wire N__12223;
    wire N__12216;
    wire N__12215;
    wire N__12214;
    wire N__12207;
    wire N__12206;
    wire N__12205;
    wire N__12198;
    wire N__12197;
    wire N__12196;
    wire N__12189;
    wire N__12188;
    wire N__12187;
    wire N__12180;
    wire N__12179;
    wire N__12178;
    wire N__12171;
    wire N__12170;
    wire N__12169;
    wire N__12162;
    wire N__12161;
    wire N__12160;
    wire N__12153;
    wire N__12152;
    wire N__12151;
    wire N__12144;
    wire N__12143;
    wire N__12142;
    wire N__12135;
    wire N__12134;
    wire N__12133;
    wire N__12126;
    wire N__12125;
    wire N__12124;
    wire N__12117;
    wire N__12116;
    wire N__12115;
    wire N__12108;
    wire N__12107;
    wire N__12106;
    wire N__12099;
    wire N__12098;
    wire N__12097;
    wire N__12090;
    wire N__12089;
    wire N__12088;
    wire N__12081;
    wire N__12080;
    wire N__12079;
    wire N__12072;
    wire N__12071;
    wire N__12070;
    wire N__12063;
    wire N__12062;
    wire N__12061;
    wire N__12054;
    wire N__12053;
    wire N__12052;
    wire N__12045;
    wire N__12044;
    wire N__12043;
    wire N__12036;
    wire N__12035;
    wire N__12034;
    wire N__12027;
    wire N__12026;
    wire N__12025;
    wire N__12018;
    wire N__12017;
    wire N__12016;
    wire N__12009;
    wire N__12008;
    wire N__12007;
    wire N__12000;
    wire N__11999;
    wire N__11998;
    wire N__11991;
    wire N__11990;
    wire N__11989;
    wire N__11982;
    wire N__11981;
    wire N__11980;
    wire N__11973;
    wire N__11972;
    wire N__11971;
    wire N__11964;
    wire N__11963;
    wire N__11962;
    wire N__11955;
    wire N__11954;
    wire N__11953;
    wire N__11946;
    wire N__11945;
    wire N__11944;
    wire N__11937;
    wire N__11936;
    wire N__11935;
    wire N__11928;
    wire N__11927;
    wire N__11926;
    wire N__11919;
    wire N__11918;
    wire N__11917;
    wire N__11910;
    wire N__11909;
    wire N__11908;
    wire N__11901;
    wire N__11900;
    wire N__11899;
    wire N__11892;
    wire N__11891;
    wire N__11890;
    wire N__11883;
    wire N__11882;
    wire N__11881;
    wire N__11874;
    wire N__11873;
    wire N__11872;
    wire N__11865;
    wire N__11864;
    wire N__11863;
    wire N__11856;
    wire N__11855;
    wire N__11854;
    wire N__11847;
    wire N__11846;
    wire N__11845;
    wire N__11838;
    wire N__11837;
    wire N__11836;
    wire N__11829;
    wire N__11828;
    wire N__11827;
    wire N__11820;
    wire N__11819;
    wire N__11818;
    wire N__11811;
    wire N__11810;
    wire N__11809;
    wire N__11802;
    wire N__11801;
    wire N__11800;
    wire N__11783;
    wire N__11780;
    wire N__11777;
    wire N__11774;
    wire N__11771;
    wire N__11768;
    wire N__11765;
    wire N__11762;
    wire N__11759;
    wire N__11756;
    wire N__11753;
    wire N__11750;
    wire N__11747;
    wire N__11744;
    wire N__11741;
    wire N__11738;
    wire N__11735;
    wire N__11732;
    wire N__11729;
    wire N__11726;
    wire N__11723;
    wire N__11720;
    wire N__11717;
    wire N__11714;
    wire N__11711;
    wire N__11708;
    wire N__11705;
    wire N__11702;
    wire N__11699;
    wire N__11696;
    wire N__11693;
    wire N__11690;
    wire N__11687;
    wire N__11684;
    wire N__11681;
    wire N__11678;
    wire N__11675;
    wire N__11672;
    wire N__11669;
    wire N__11666;
    wire N__11663;
    wire N__11660;
    wire N__11657;
    wire N__11654;
    wire N__11651;
    wire N__11648;
    wire N__11645;
    wire N__11642;
    wire N__11639;
    wire N__11636;
    wire N__11633;
    wire N__11630;
    wire N__11627;
    wire N__11624;
    wire N__11621;
    wire N__11618;
    wire N__11615;
    wire N__11612;
    wire N__11609;
    wire N__11606;
    wire N__11603;
    wire N__11600;
    wire N__11597;
    wire N__11594;
    wire N__11591;
    wire N__11588;
    wire N__11585;
    wire N__11582;
    wire N__11579;
    wire N__11576;
    wire N__11573;
    wire N__11570;
    wire N__11567;
    wire N__11564;
    wire N__11561;
    wire N__11558;
    wire N__11555;
    wire N__11552;
    wire N__11549;
    wire N__11546;
    wire N__11543;
    wire N__11540;
    wire N__11537;
    wire N__11534;
    wire N__11531;
    wire N__11528;
    wire N__11525;
    wire N__11522;
    wire N__11519;
    wire N__11516;
    wire N__11513;
    wire N__11510;
    wire N__11507;
    wire N__11504;
    wire N__11501;
    wire N__11498;
    wire N__11495;
    wire N__11492;
    wire N__11489;
    wire N__11486;
    wire N__11483;
    wire N__11482;
    wire N__11479;
    wire N__11476;
    wire N__11473;
    wire N__11470;
    wire N__11467;
    wire N__11464;
    wire N__11461;
    wire N__11458;
    wire N__11455;
    wire N__11452;
    wire N__11449;
    wire N__11446;
    wire N__11443;
    wire N__11440;
    wire N__11435;
    wire N__11432;
    wire N__11429;
    wire N__11426;
    wire N__11423;
    wire N__11420;
    wire N__11417;
    wire N__11414;
    wire N__11411;
    wire N__11408;
    wire N__11405;
    wire N__11402;
    wire N__11399;
    wire N__11396;
    wire N__11393;
    wire N__11390;
    wire N__11387;
    wire N__11384;
    wire N__11381;
    wire N__11378;
    wire N__11375;
    wire N__11372;
    wire N__11369;
    wire N__11366;
    wire N__11363;
    wire N__11360;
    wire N__11357;
    wire N__11354;
    wire N__11351;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11333;
    wire N__11330;
    wire N__11327;
    wire N__11324;
    wire N__11321;
    wire N__11318;
    wire N__11315;
    wire N__11312;
    wire N__11309;
    wire N__11306;
    wire N__11303;
    wire N__11302;
    wire N__11299;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11284;
    wire N__11281;
    wire N__11278;
    wire N__11275;
    wire N__11272;
    wire N__11269;
    wire N__11266;
    wire N__11263;
    wire N__11260;
    wire N__11255;
    wire N__11252;
    wire N__11249;
    wire N__11246;
    wire N__11243;
    wire N__11240;
    wire N__11237;
    wire N__11234;
    wire N__11231;
    wire N__11228;
    wire N__11225;
    wire N__11224;
    wire N__11221;
    wire N__11218;
    wire N__11215;
    wire N__11212;
    wire N__11209;
    wire N__11206;
    wire N__11203;
    wire N__11200;
    wire N__11197;
    wire N__11194;
    wire N__11189;
    wire N__11186;
    wire N__11183;
    wire N__11180;
    wire N__11177;
    wire N__11174;
    wire N__11171;
    wire N__11170;
    wire N__11169;
    wire N__11168;
    wire N__11167;
    wire N__11166;
    wire N__11165;
    wire N__11164;
    wire N__11163;
    wire N__11162;
    wire N__11161;
    wire N__11158;
    wire N__11155;
    wire N__11152;
    wire N__11151;
    wire N__11148;
    wire N__11145;
    wire N__11144;
    wire N__11143;
    wire N__11140;
    wire N__11139;
    wire N__11134;
    wire N__11131;
    wire N__11130;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11122;
    wire N__11121;
    wire N__11120;
    wire N__11119;
    wire N__11118;
    wire N__11117;
    wire N__11112;
    wire N__11111;
    wire N__11108;
    wire N__11105;
    wire N__11102;
    wire N__11099;
    wire N__11094;
    wire N__11093;
    wire N__11090;
    wire N__11087;
    wire N__11086;
    wire N__11083;
    wire N__11080;
    wire N__11077;
    wire N__11076;
    wire N__11073;
    wire N__11068;
    wire N__11065;
    wire N__11062;
    wire N__11061;
    wire N__11058;
    wire N__11055;
    wire N__11052;
    wire N__11049;
    wire N__11048;
    wire N__11047;
    wire N__11046;
    wire N__11043;
    wire N__11040;
    wire N__11037;
    wire N__11034;
    wire N__11031;
    wire N__11026;
    wire N__11023;
    wire N__11018;
    wire N__11015;
    wire N__11012;
    wire N__11007;
    wire N__11004;
    wire N__11001;
    wire N__10996;
    wire N__10993;
    wire N__10990;
    wire N__10985;
    wire N__10980;
    wire N__10977;
    wire N__10972;
    wire N__10971;
    wire N__10970;
    wire N__10967;
    wire N__10964;
    wire N__10959;
    wire N__10954;
    wire N__10951;
    wire N__10946;
    wire N__10939;
    wire N__10936;
    wire N__10933;
    wire N__10928;
    wire N__10921;
    wire N__10918;
    wire N__10915;
    wire N__10912;
    wire N__10907;
    wire N__10900;
    wire N__10895;
    wire N__10884;
    wire N__10881;
    wire N__10878;
    wire N__10865;
    wire N__10862;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10847;
    wire N__10844;
    wire N__10841;
    wire N__10838;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10826;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10811;
    wire N__10808;
    wire N__10805;
    wire N__10802;
    wire N__10799;
    wire N__10796;
    wire N__10793;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10772;
    wire N__10769;
    wire N__10766;
    wire N__10763;
    wire N__10760;
    wire N__10757;
    wire N__10754;
    wire N__10751;
    wire N__10748;
    wire N__10745;
    wire N__10742;
    wire N__10739;
    wire N__10736;
    wire N__10733;
    wire N__10730;
    wire N__10727;
    wire N__10724;
    wire N__10721;
    wire N__10718;
    wire N__10715;
    wire N__10712;
    wire N__10709;
    wire N__10706;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10691;
    wire N__10688;
    wire N__10685;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10670;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10655;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10639;
    wire N__10636;
    wire N__10633;
    wire N__10630;
    wire N__10627;
    wire N__10624;
    wire N__10621;
    wire N__10618;
    wire N__10615;
    wire N__10610;
    wire N__10607;
    wire N__10604;
    wire N__10601;
    wire N__10598;
    wire N__10595;
    wire N__10592;
    wire N__10589;
    wire N__10586;
    wire N__10583;
    wire N__10580;
    wire N__10577;
    wire N__10574;
    wire N__10571;
    wire N__10568;
    wire N__10565;
    wire N__10562;
    wire N__10559;
    wire N__10556;
    wire N__10553;
    wire N__10550;
    wire N__10547;
    wire N__10544;
    wire N__10541;
    wire N__10538;
    wire N__10535;
    wire N__10532;
    wire N__10529;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10517;
    wire N__10514;
    wire N__10511;
    wire N__10508;
    wire N__10505;
    wire N__10502;
    wire N__10499;
    wire N__10496;
    wire N__10493;
    wire N__10490;
    wire N__10487;
    wire N__10484;
    wire N__10481;
    wire N__10478;
    wire N__10475;
    wire N__10472;
    wire N__10471;
    wire N__10468;
    wire N__10465;
    wire N__10462;
    wire N__10461;
    wire N__10458;
    wire N__10455;
    wire N__10452;
    wire N__10449;
    wire N__10446;
    wire N__10443;
    wire N__10440;
    wire N__10435;
    wire N__10432;
    wire N__10429;
    wire N__10426;
    wire N__10421;
    wire N__10418;
    wire N__10415;
    wire N__10412;
    wire N__10409;
    wire N__10408;
    wire N__10407;
    wire N__10406;
    wire N__10405;
    wire N__10404;
    wire N__10403;
    wire N__10396;
    wire N__10395;
    wire N__10394;
    wire N__10393;
    wire N__10390;
    wire N__10385;
    wire N__10382;
    wire N__10381;
    wire N__10380;
    wire N__10379;
    wire N__10376;
    wire N__10371;
    wire N__10368;
    wire N__10367;
    wire N__10360;
    wire N__10357;
    wire N__10354;
    wire N__10351;
    wire N__10350;
    wire N__10343;
    wire N__10340;
    wire N__10331;
    wire N__10328;
    wire N__10327;
    wire N__10326;
    wire N__10321;
    wire N__10316;
    wire N__10313;
    wire N__10310;
    wire N__10307;
    wire N__10304;
    wire N__10301;
    wire N__10298;
    wire N__10289;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10274;
    wire N__10271;
    wire N__10268;
    wire N__10265;
    wire N__10262;
    wire N__10259;
    wire N__10256;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10244;
    wire N__10241;
    wire N__10238;
    wire N__10235;
    wire N__10232;
    wire N__10229;
    wire N__10226;
    wire N__10223;
    wire N__10220;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10202;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10181;
    wire N__10178;
    wire N__10175;
    wire N__10174;
    wire N__10171;
    wire N__10168;
    wire N__10165;
    wire N__10162;
    wire N__10159;
    wire N__10156;
    wire N__10153;
    wire N__10150;
    wire N__10147;
    wire N__10144;
    wire N__10141;
    wire N__10138;
    wire N__10133;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10118;
    wire N__10115;
    wire N__10112;
    wire N__10109;
    wire N__10106;
    wire N__10103;
    wire N__10100;
    wire N__10097;
    wire N__10094;
    wire N__10091;
    wire N__10090;
    wire N__10087;
    wire N__10086;
    wire N__10085;
    wire N__10084;
    wire N__10083;
    wire N__10082;
    wire N__10081;
    wire N__10078;
    wire N__10077;
    wire N__10074;
    wire N__10073;
    wire N__10066;
    wire N__10059;
    wire N__10058;
    wire N__10057;
    wire N__10052;
    wire N__10051;
    wire N__10050;
    wire N__10049;
    wire N__10048;
    wire N__10047;
    wire N__10044;
    wire N__10043;
    wire N__10042;
    wire N__10041;
    wire N__10040;
    wire N__10039;
    wire N__10038;
    wire N__10035;
    wire N__10032;
    wire N__10029;
    wire N__10026;
    wire N__10023;
    wire N__10020;
    wire N__10015;
    wire N__10014;
    wire N__10013;
    wire N__10012;
    wire N__10011;
    wire N__10010;
    wire N__10009;
    wire N__10008;
    wire N__10007;
    wire N__10006;
    wire N__10005;
    wire N__10004;
    wire N__10003;
    wire N__10002;
    wire N__10001;
    wire N__10000;
    wire N__9999;
    wire N__9996;
    wire N__9993;
    wire N__9992;
    wire N__9989;
    wire N__9988;
    wire N__9985;
    wire N__9980;
    wire N__9975;
    wire N__9972;
    wire N__9969;
    wire N__9966;
    wire N__9957;
    wire N__9952;
    wire N__9949;
    wire N__9946;
    wire N__9943;
    wire N__9940;
    wire N__9939;
    wire N__9938;
    wire N__9931;
    wire N__9914;
    wire N__9901;
    wire N__9900;
    wire N__9899;
    wire N__9898;
    wire N__9897;
    wire N__9896;
    wire N__9895;
    wire N__9884;
    wire N__9881;
    wire N__9874;
    wire N__9865;
    wire N__9864;
    wire N__9861;
    wire N__9860;
    wire N__9857;
    wire N__9852;
    wire N__9851;
    wire N__9850;
    wire N__9847;
    wire N__9846;
    wire N__9843;
    wire N__9842;
    wire N__9841;
    wire N__9840;
    wire N__9839;
    wire N__9838;
    wire N__9837;
    wire N__9836;
    wire N__9835;
    wire N__9834;
    wire N__9831;
    wire N__9830;
    wire N__9827;
    wire N__9824;
    wire N__9823;
    wire N__9820;
    wire N__9819;
    wire N__9814;
    wire N__9809;
    wire N__9802;
    wire N__9797;
    wire N__9784;
    wire N__9767;
    wire N__9752;
    wire N__9747;
    wire N__9744;
    wire N__9733;
    wire N__9730;
    wire N__9727;
    wire N__9724;
    wire N__9719;
    wire N__9718;
    wire N__9717;
    wire N__9710;
    wire N__9709;
    wire N__9708;
    wire N__9707;
    wire N__9706;
    wire N__9705;
    wire N__9704;
    wire N__9703;
    wire N__9702;
    wire N__9701;
    wire N__9700;
    wire N__9699;
    wire N__9698;
    wire N__9697;
    wire N__9696;
    wire N__9695;
    wire N__9694;
    wire N__9693;
    wire N__9692;
    wire N__9691;
    wire N__9690;
    wire N__9687;
    wire N__9684;
    wire N__9683;
    wire N__9682;
    wire N__9681;
    wire N__9680;
    wire N__9679;
    wire N__9676;
    wire N__9675;
    wire N__9674;
    wire N__9671;
    wire N__9664;
    wire N__9655;
    wire N__9652;
    wire N__9649;
    wire N__9648;
    wire N__9647;
    wire N__9646;
    wire N__9645;
    wire N__9644;
    wire N__9643;
    wire N__9642;
    wire N__9639;
    wire N__9632;
    wire N__9627;
    wire N__9622;
    wire N__9621;
    wire N__9620;
    wire N__9619;
    wire N__9618;
    wire N__9617;
    wire N__9616;
    wire N__9615;
    wire N__9614;
    wire N__9613;
    wire N__9612;
    wire N__9611;
    wire N__9610;
    wire N__9609;
    wire N__9608;
    wire N__9603;
    wire N__9598;
    wire N__9591;
    wire N__9588;
    wire N__9583;
    wire N__9582;
    wire N__9581;
    wire N__9580;
    wire N__9579;
    wire N__9578;
    wire N__9577;
    wire N__9576;
    wire N__9575;
    wire N__9574;
    wire N__9573;
    wire N__9572;
    wire N__9571;
    wire N__9570;
    wire N__9569;
    wire N__9568;
    wire N__9567;
    wire N__9564;
    wire N__9559;
    wire N__9554;
    wire N__9539;
    wire N__9534;
    wire N__9531;
    wire N__9528;
    wire N__9515;
    wire N__9498;
    wire N__9487;
    wire N__9470;
    wire N__9457;
    wire N__9454;
    wire N__9451;
    wire N__9422;
    wire N__9419;
    wire N__9418;
    wire N__9417;
    wire N__9416;
    wire N__9413;
    wire N__9412;
    wire N__9411;
    wire N__9410;
    wire N__9409;
    wire N__9408;
    wire N__9407;
    wire N__9406;
    wire N__9405;
    wire N__9404;
    wire N__9403;
    wire N__9402;
    wire N__9401;
    wire N__9400;
    wire N__9399;
    wire N__9398;
    wire N__9397;
    wire N__9396;
    wire N__9395;
    wire N__9394;
    wire N__9393;
    wire N__9392;
    wire N__9391;
    wire N__9390;
    wire N__9389;
    wire N__9388;
    wire N__9387;
    wire N__9386;
    wire N__9385;
    wire N__9384;
    wire N__9317;
    wire N__9314;
    wire N__9313;
    wire N__9312;
    wire N__9311;
    wire N__9310;
    wire N__9309;
    wire N__9308;
    wire N__9307;
    wire N__9306;
    wire N__9305;
    wire N__9304;
    wire N__9303;
    wire N__9302;
    wire N__9301;
    wire N__9300;
    wire N__9299;
    wire N__9298;
    wire N__9297;
    wire N__9296;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9247;
    wire N__9246;
    wire N__9245;
    wire N__9244;
    wire N__9243;
    wire N__9242;
    wire N__9241;
    wire N__9240;
    wire N__9239;
    wire N__9238;
    wire N__9237;
    wire N__9236;
    wire N__9235;
    wire N__9234;
    wire N__9233;
    wire N__9232;
    wire N__9231;
    wire N__9230;
    wire N__9229;
    wire N__9228;
    wire N__9227;
    wire N__9226;
    wire N__9225;
    wire N__9224;
    wire N__9221;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9145;
    wire N__9144;
    wire N__9141;
    wire N__9138;
    wire N__9135;
    wire N__9128;
    wire N__9125;
    wire N__9122;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9107;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9094;
    wire N__9091;
    wire N__9090;
    wire N__9087;
    wire N__9084;
    wire N__9081;
    wire N__9078;
    wire N__9075;
    wire N__9072;
    wire N__9069;
    wire N__9064;
    wire N__9059;
    wire N__9056;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9025;
    wire N__9024;
    wire N__9021;
    wire N__9018;
    wire N__9015;
    wire N__9012;
    wire N__9009;
    wire N__9006;
    wire N__9003;
    wire N__9000;
    wire N__8997;
    wire N__8994;
    wire N__8989;
    wire N__8986;
    wire N__8983;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8960;
    wire N__8957;
    wire N__8954;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8921;
    wire N__8920;
    wire N__8917;
    wire N__8914;
    wire N__8911;
    wire N__8908;
    wire N__8905;
    wire N__8902;
    wire N__8899;
    wire N__8896;
    wire N__8893;
    wire N__8890;
    wire N__8885;
    wire N__8882;
    wire N__8879;
    wire N__8876;
    wire N__8873;
    wire N__8870;
    wire N__8867;
    wire N__8864;
    wire N__8861;
    wire N__8858;
    wire N__8855;
    wire N__8852;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8824;
    wire N__8823;
    wire N__8820;
    wire N__8817;
    wire N__8814;
    wire N__8811;
    wire N__8808;
    wire N__8805;
    wire N__8800;
    wire N__8797;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8777;
    wire N__8774;
    wire N__8771;
    wire N__8768;
    wire N__8765;
    wire N__8762;
    wire N__8761;
    wire N__8760;
    wire N__8757;
    wire N__8754;
    wire N__8751;
    wire N__8748;
    wire N__8745;
    wire N__8742;
    wire N__8739;
    wire N__8736;
    wire N__8733;
    wire N__8728;
    wire N__8725;
    wire N__8722;
    wire N__8719;
    wire N__8714;
    wire N__8711;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8696;
    wire N__8693;
    wire N__8690;
    wire N__8687;
    wire N__8686;
    wire N__8683;
    wire N__8682;
    wire N__8679;
    wire N__8676;
    wire N__8673;
    wire N__8670;
    wire N__8665;
    wire N__8662;
    wire N__8659;
    wire N__8656;
    wire N__8653;
    wire N__8650;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8596;
    wire N__8593;
    wire N__8590;
    wire N__8587;
    wire N__8584;
    wire N__8581;
    wire N__8578;
    wire N__8575;
    wire N__8572;
    wire N__8569;
    wire N__8566;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8527;
    wire N__8524;
    wire N__8521;
    wire N__8518;
    wire N__8517;
    wire N__8514;
    wire N__8511;
    wire N__8508;
    wire N__8505;
    wire N__8500;
    wire N__8497;
    wire N__8494;
    wire N__8491;
    wire N__8488;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8452;
    wire N__8449;
    wire N__8448;
    wire N__8445;
    wire N__8442;
    wire N__8439;
    wire N__8436;
    wire N__8431;
    wire N__8428;
    wire N__8425;
    wire N__8422;
    wire N__8419;
    wire N__8416;
    wire N__8413;
    wire N__8408;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8384;
    wire N__8381;
    wire N__8378;
    wire N__8375;
    wire N__8372;
    wire N__8371;
    wire N__8368;
    wire N__8365;
    wire N__8362;
    wire N__8359;
    wire N__8356;
    wire N__8353;
    wire N__8352;
    wire N__8349;
    wire N__8346;
    wire N__8343;
    wire N__8340;
    wire N__8337;
    wire N__8334;
    wire N__8331;
    wire N__8326;
    wire N__8321;
    wire N__8318;
    wire N__8315;
    wire N__8312;
    wire N__8309;
    wire N__8306;
    wire N__8303;
    wire N__8300;
    wire N__8297;
    wire N__8294;
    wire N__8291;
    wire N__8288;
    wire N__8285;
    wire N__8282;
    wire N__8279;
    wire N__8276;
    wire N__8273;
    wire N__8272;
    wire N__8271;
    wire N__8268;
    wire N__8265;
    wire N__8262;
    wire N__8255;
    wire N__8252;
    wire N__8249;
    wire N__8246;
    wire N__8243;
    wire N__8240;
    wire N__8237;
    wire N__8236;
    wire N__8235;
    wire N__8234;
    wire N__8231;
    wire N__8228;
    wire N__8225;
    wire N__8222;
    wire N__8213;
    wire N__8212;
    wire N__8211;
    wire N__8208;
    wire N__8205;
    wire N__8202;
    wire N__8201;
    wire N__8198;
    wire N__8195;
    wire N__8192;
    wire N__8189;
    wire N__8184;
    wire N__8179;
    wire N__8176;
    wire N__8173;
    wire N__8168;
    wire N__8165;
    wire N__8164;
    wire N__8163;
    wire N__8160;
    wire N__8157;
    wire N__8154;
    wire N__8151;
    wire N__8146;
    wire N__8143;
    wire N__8140;
    wire N__8137;
    wire N__8134;
    wire N__8131;
    wire N__8128;
    wire N__8123;
    wire N__8120;
    wire N__8117;
    wire N__8114;
    wire N__8111;
    wire N__8108;
    wire N__8105;
    wire N__8102;
    wire N__8099;
    wire N__8096;
    wire N__8093;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8069;
    wire N__8068;
    wire N__8065;
    wire N__8062;
    wire N__8059;
    wire N__8056;
    wire N__8051;
    wire N__8050;
    wire N__8049;
    wire N__8046;
    wire N__8043;
    wire N__8040;
    wire N__8037;
    wire N__8034;
    wire N__8033;
    wire N__8030;
    wire N__8025;
    wire N__8022;
    wire N__8019;
    wire N__8016;
    wire N__8015;
    wire N__8012;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__7996;
    wire N__7993;
    wire N__7990;
    wire N__7987;
    wire N__7982;
    wire N__7979;
    wire N__7976;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7957;
    wire N__7954;
    wire N__7951;
    wire N__7948;
    wire N__7945;
    wire N__7942;
    wire N__7939;
    wire N__7934;
    wire N__7931;
    wire N__7928;
    wire N__7925;
    wire N__7922;
    wire N__7919;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7904;
    wire N__7901;
    wire N__7898;
    wire N__7895;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7877;
    wire N__7874;
    wire N__7871;
    wire N__7868;
    wire N__7865;
    wire N__7862;
    wire N__7859;
    wire N__7856;
    wire N__7853;
    wire N__7850;
    wire N__7847;
    wire N__7844;
    wire N__7841;
    wire N__7838;
    wire N__7835;
    wire N__7832;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7814;
    wire N__7813;
    wire N__7810;
    wire N__7807;
    wire N__7804;
    wire N__7801;
    wire N__7798;
    wire N__7795;
    wire N__7792;
    wire N__7789;
    wire N__7786;
    wire N__7783;
    wire N__7780;
    wire N__7777;
    wire N__7772;
    wire N__7769;
    wire N__7766;
    wire N__7763;
    wire N__7760;
    wire N__7757;
    wire N__7754;
    wire N__7751;
    wire N__7748;
    wire N__7745;
    wire N__7742;
    wire N__7739;
    wire N__7736;
    wire N__7733;
    wire N__7730;
    wire N__7727;
    wire N__7724;
    wire N__7721;
    wire N__7718;
    wire N__7715;
    wire N__7712;
    wire N__7709;
    wire N__7706;
    wire N__7703;
    wire N__7700;
    wire N__7699;
    wire N__7696;
    wire N__7693;
    wire N__7690;
    wire N__7687;
    wire N__7684;
    wire N__7681;
    wire N__7678;
    wire N__7675;
    wire N__7672;
    wire N__7669;
    wire N__7664;
    wire N__7661;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7637;
    wire N__7634;
    wire N__7631;
    wire N__7628;
    wire N__7625;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7613;
    wire N__7610;
    wire N__7607;
    wire N__7606;
    wire N__7603;
    wire N__7600;
    wire N__7597;
    wire N__7594;
    wire N__7591;
    wire N__7588;
    wire N__7583;
    wire N__7580;
    wire N__7577;
    wire N__7574;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7550;
    wire N__7547;
    wire N__7546;
    wire N__7545;
    wire N__7542;
    wire N__7539;
    wire N__7536;
    wire N__7531;
    wire N__7528;
    wire N__7525;
    wire N__7522;
    wire N__7519;
    wire N__7514;
    wire N__7511;
    wire N__7508;
    wire N__7505;
    wire N__7502;
    wire N__7499;
    wire N__7496;
    wire N__7493;
    wire N__7490;
    wire N__7487;
    wire N__7486;
    wire N__7485;
    wire N__7482;
    wire N__7479;
    wire N__7476;
    wire N__7471;
    wire N__7468;
    wire N__7465;
    wire N__7462;
    wire N__7459;
    wire N__7456;
    wire N__7453;
    wire N__7450;
    wire N__7447;
    wire N__7442;
    wire N__7439;
    wire N__7436;
    wire N__7433;
    wire N__7430;
    wire N__7427;
    wire N__7424;
    wire N__7421;
    wire N__7418;
    wire N__7415;
    wire N__7412;
    wire N__7409;
    wire N__7408;
    wire N__7405;
    wire N__7402;
    wire N__7401;
    wire N__7398;
    wire N__7395;
    wire N__7392;
    wire N__7389;
    wire N__7384;
    wire N__7381;
    wire N__7378;
    wire N__7375;
    wire N__7372;
    wire N__7367;
    wire N__7364;
    wire N__7361;
    wire N__7358;
    wire N__7355;
    wire N__7352;
    wire N__7349;
    wire N__7346;
    wire N__7343;
    wire N__7340;
    wire N__7337;
    wire N__7334;
    wire N__7331;
    wire N__7328;
    wire N__7325;
    wire N__7322;
    wire N__7319;
    wire N__7318;
    wire N__7317;
    wire N__7314;
    wire N__7311;
    wire N__7308;
    wire N__7305;
    wire N__7302;
    wire N__7299;
    wire N__7296;
    wire N__7291;
    wire N__7286;
    wire N__7283;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7271;
    wire N__7268;
    wire N__7265;
    wire N__7262;
    wire N__7259;
    wire N__7256;
    wire N__7253;
    wire N__7250;
    wire N__7247;
    wire N__7246;
    wire N__7243;
    wire N__7240;
    wire N__7235;
    wire N__7234;
    wire N__7233;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7223;
    wire N__7220;
    wire N__7217;
    wire N__7212;
    wire N__7205;
    wire N__7202;
    wire N__7199;
    wire N__7198;
    wire N__7197;
    wire N__7194;
    wire N__7193;
    wire N__7190;
    wire N__7189;
    wire N__7188;
    wire N__7185;
    wire N__7184;
    wire N__7181;
    wire N__7178;
    wire N__7171;
    wire N__7166;
    wire N__7163;
    wire N__7156;
    wire N__7155;
    wire N__7150;
    wire N__7147;
    wire N__7146;
    wire N__7143;
    wire N__7138;
    wire N__7133;
    wire N__7130;
    wire N__7127;
    wire N__7126;
    wire N__7125;
    wire N__7124;
    wire N__7123;
    wire N__7120;
    wire N__7117;
    wire N__7108;
    wire N__7103;
    wire N__7100;
    wire N__7097;
    wire N__7094;
    wire N__7091;
    wire N__7088;
    wire N__7085;
    wire N__7084;
    wire N__7083;
    wire N__7082;
    wire N__7081;
    wire N__7078;
    wire N__7075;
    wire N__7072;
    wire N__7069;
    wire N__7066;
    wire N__7063;
    wire N__7052;
    wire N__7051;
    wire N__7048;
    wire N__7045;
    wire N__7040;
    wire N__7037;
    wire N__7036;
    wire N__7035;
    wire N__7034;
    wire N__7031;
    wire N__7028;
    wire N__7025;
    wire N__7022;
    wire N__7013;
    wire N__7010;
    wire N__7007;
    wire N__7004;
    wire N__7003;
    wire N__7000;
    wire N__6997;
    wire N__6994;
    wire N__6991;
    wire N__6988;
    wire N__6985;
    wire N__6980;
    wire N__6977;
    wire N__6976;
    wire N__6975;
    wire N__6972;
    wire N__6969;
    wire N__6966;
    wire N__6959;
    wire N__6958;
    wire N__6955;
    wire N__6952;
    wire N__6947;
    wire N__6944;
    wire N__6943;
    wire N__6942;
    wire N__6941;
    wire N__6940;
    wire N__6939;
    wire N__6936;
    wire N__6927;
    wire N__6924;
    wire N__6917;
    wire N__6914;
    wire N__6913;
    wire N__6910;
    wire N__6907;
    wire N__6904;
    wire N__6899;
    wire N__6896;
    wire N__6893;
    wire N__6892;
    wire N__6891;
    wire N__6888;
    wire N__6883;
    wire N__6878;
    wire N__6875;
    wire N__6874;
    wire N__6871;
    wire N__6870;
    wire N__6867;
    wire N__6864;
    wire N__6861;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6847;
    wire N__6844;
    wire N__6843;
    wire N__6842;
    wire N__6841;
    wire N__6838;
    wire N__6837;
    wire N__6836;
    wire N__6835;
    wire N__6832;
    wire N__6825;
    wire N__6820;
    wire N__6815;
    wire N__6812;
    wire N__6807;
    wire N__6804;
    wire N__6801;
    wire N__6798;
    wire N__6795;
    wire N__6792;
    wire N__6789;
    wire N__6786;
    wire N__6779;
    wire N__6776;
    wire N__6773;
    wire N__6772;
    wire N__6771;
    wire N__6770;
    wire N__6769;
    wire N__6764;
    wire N__6761;
    wire N__6756;
    wire N__6749;
    wire N__6748;
    wire N__6747;
    wire N__6746;
    wire N__6745;
    wire N__6744;
    wire N__6743;
    wire N__6742;
    wire N__6737;
    wire N__6730;
    wire N__6725;
    wire N__6722;
    wire N__6719;
    wire N__6716;
    wire N__6713;
    wire N__6710;
    wire N__6709;
    wire N__6704;
    wire N__6701;
    wire N__6698;
    wire N__6695;
    wire N__6688;
    wire N__6685;
    wire N__6680;
    wire N__6677;
    wire N__6674;
    wire N__6671;
    wire N__6668;
    wire N__6665;
    wire N__6662;
    wire N__6659;
    wire N__6656;
    wire N__6653;
    wire N__6650;
    wire N__6647;
    wire N__6644;
    wire N__6641;
    wire N__6638;
    wire N__6635;
    wire N__6632;
    wire N__6629;
    wire N__6626;
    wire N__6623;
    wire N__6620;
    wire N__6617;
    wire N__6614;
    wire N__6611;
    wire N__6608;
    wire N__6605;
    wire N__6602;
    wire N__6599;
    wire N__6596;
    wire N__6593;
    wire N__6590;
    wire N__6587;
    wire N__6584;
    wire N__6581;
    wire N__6578;
    wire N__6575;
    wire N__6572;
    wire N__6569;
    wire N__6566;
    wire N__6563;
    wire N__6560;
    wire N__6557;
    wire N__6554;
    wire N__6551;
    wire N__6548;
    wire N__6545;
    wire N__6542;
    wire N__6539;
    wire N__6536;
    wire N__6533;
    wire N__6530;
    wire N__6527;
    wire N__6524;
    wire N__6521;
    wire N__6518;
    wire N__6515;
    wire N__6512;
    wire N__6509;
    wire N__6506;
    wire N__6503;
    wire N__6500;
    wire N__6499;
    wire N__6498;
    wire N__6495;
    wire N__6492;
    wire N__6489;
    wire N__6482;
    wire N__6481;
    wire N__6478;
    wire N__6475;
    wire N__6472;
    wire N__6469;
    wire N__6466;
    wire N__6465;
    wire N__6462;
    wire N__6459;
    wire N__6456;
    wire N__6449;
    wire N__6446;
    wire N__6443;
    wire N__6440;
    wire N__6437;
    wire N__6436;
    wire N__6435;
    wire N__6434;
    wire N__6433;
    wire N__6432;
    wire N__6429;
    wire N__6424;
    wire N__6419;
    wire N__6416;
    wire N__6407;
    wire N__6404;
    wire N__6401;
    wire N__6398;
    wire N__6395;
    wire N__6392;
    wire N__6389;
    wire N__6386;
    wire N__6383;
    wire N__6380;
    wire N__6377;
    wire N__6374;
    wire N__6371;
    wire N__6368;
    wire N__6365;
    wire N__6362;
    wire N__6359;
    wire N__6358;
    wire N__6357;
    wire N__6356;
    wire N__6355;
    wire N__6352;
    wire N__6349;
    wire N__6342;
    wire N__6335;
    wire N__6334;
    wire N__6329;
    wire N__6326;
    wire N__6323;
    wire N__6320;
    wire N__6317;
    wire N__6314;
    wire N__6311;
    wire N__6310;
    wire N__6307;
    wire N__6304;
    wire N__6301;
    wire N__6298;
    wire N__6293;
    wire N__6290;
    wire N__6287;
    wire N__6284;
    wire N__6281;
    wire N__6278;
    wire N__6275;
    wire N__6272;
    wire N__6269;
    wire N__6266;
    wire N__6263;
    wire N__6260;
    wire N__6257;
    wire N__6254;
    wire N__6251;
    wire N__6248;
    wire N__6245;
    wire N__6242;
    wire N__6239;
    wire N__6236;
    wire N__6233;
    wire N__6230;
    wire N__6227;
    wire N__6224;
    wire N__6221;
    wire N__6218;
    wire N__6215;
    wire N__6212;
    wire N__6209;
    wire N__6206;
    wire N__6203;
    wire N__6200;
    wire N__6197;
    wire N__6194;
    wire N__6191;
    wire N__6188;
    wire N__6185;
    wire N__6184;
    wire N__6181;
    wire N__6178;
    wire N__6173;
    wire N__6170;
    wire N__6167;
    wire N__6164;
    wire N__6161;
    wire N__6158;
    wire N__6155;
    wire N__6152;
    wire N__6149;
    wire N__6146;
    wire N__6143;
    wire N__6140;
    wire N__6137;
    wire N__6134;
    wire N__6133;
    wire N__6130;
    wire N__6127;
    wire N__6124;
    wire N__6123;
    wire N__6122;
    wire N__6119;
    wire N__6116;
    wire N__6113;
    wire N__6110;
    wire N__6107;
    wire N__6104;
    wire N__6101;
    wire N__6098;
    wire N__6095;
    wire N__6090;
    wire N__6087;
    wire N__6084;
    wire N__6081;
    wire N__6078;
    wire N__6075;
    wire N__6072;
    wire N__6069;
    wire N__6066;
    wire N__6061;
    wire N__6056;
    wire N__6053;
    wire N__6050;
    wire N__6047;
    wire N__6044;
    wire N__6043;
    wire N__6038;
    wire N__6035;
    wire N__6034;
    wire N__6031;
    wire N__6028;
    wire N__6023;
    wire N__6020;
    wire N__6017;
    wire N__6014;
    wire N__6011;
    wire N__6008;
    wire N__6007;
    wire N__6004;
    wire N__6001;
    wire N__5996;
    wire N__5993;
    wire N__5990;
    wire N__5987;
    wire N__5986;
    wire N__5983;
    wire N__5980;
    wire N__5977;
    wire N__5974;
    wire N__5971;
    wire N__5968;
    wire N__5965;
    wire N__5962;
    wire N__5959;
    wire N__5956;
    wire N__5951;
    wire N__5948;
    wire N__5945;
    wire N__5942;
    wire N__5939;
    wire N__5936;
    wire N__5933;
    wire N__5930;
    wire N__5927;
    wire N__5924;
    wire N__5921;
    wire N__5918;
    wire N__5915;
    wire N__5912;
    wire N__5909;
    wire N__5906;
    wire N__5903;
    wire N__5902;
    wire N__5899;
    wire N__5896;
    wire N__5893;
    wire N__5890;
    wire N__5887;
    wire N__5884;
    wire N__5881;
    wire N__5878;
    wire N__5873;
    wire N__5870;
    wire N__5867;
    wire N__5864;
    wire N__5861;
    wire N__5858;
    wire N__5855;
    wire N__5852;
    wire N__5849;
    wire N__5846;
    wire N__5843;
    wire N__5840;
    wire N__5837;
    wire N__5834;
    wire N__5831;
    wire N__5828;
    wire N__5825;
    wire N__5822;
    wire N__5819;
    wire N__5816;
    wire N__5813;
    wire N__5810;
    wire N__5807;
    wire N__5804;
    wire N__5801;
    wire N__5798;
    wire N__5795;
    wire N__5792;
    wire N__5789;
    wire N__5786;
    wire N__5783;
    wire N__5780;
    wire N__5777;
    wire N__5774;
    wire N__5771;
    wire N__5768;
    wire N__5765;
    wire N__5762;
    wire N__5759;
    wire N__5756;
    wire N__5753;
    wire N__5750;
    wire N__5747;
    wire N__5744;
    wire N__5741;
    wire N__5738;
    wire N__5735;
    wire N__5732;
    wire N__5729;
    wire N__5726;
    wire N__5723;
    wire N__5720;
    wire N__5717;
    wire N__5714;
    wire N__5711;
    wire N__5708;
    wire N__5705;
    wire N__5702;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5681;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5669;
    wire N__5666;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5654;
    wire N__5651;
    wire N__5648;
    wire N__5645;
    wire N__5642;
    wire N__5639;
    wire N__5636;
    wire N__5633;
    wire N__5630;
    wire N__5627;
    wire N__5624;
    wire N__5621;
    wire N__5618;
    wire N__5615;
    wire N__5612;
    wire N__5609;
    wire N__5606;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5594;
    wire N__5591;
    wire N__5588;
    wire N__5585;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5567;
    wire N__5564;
    wire N__5561;
    wire N__5558;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5546;
    wire N__5543;
    wire N__5540;
    wire N__5537;
    wire N__5534;
    wire N__5531;
    wire N__5528;
    wire N__5525;
    wire N__5522;
    wire N__5519;
    wire N__5516;
    wire N__5513;
    wire N__5510;
    wire N__5507;
    wire N__5504;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5489;
    wire N__5486;
    wire N__5483;
    wire N__5480;
    wire N__5477;
    wire N__5474;
    wire N__5471;
    wire N__5468;
    wire N__5465;
    wire N__5462;
    wire N__5459;
    wire N__5456;
    wire N__5453;
    wire N__5450;
    wire N__5447;
    wire N__5444;
    wire N__5441;
    wire N__5438;
    wire N__5435;
    wire N__5432;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5393;
    wire N__5390;
    wire N__5387;
    wire N__5384;
    wire N__5381;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5330;
    wire N__5327;
    wire N__5324;
    wire N__5321;
    wire N__5318;
    wire N__5315;
    wire N__5312;
    wire N__5309;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5288;
    wire N__5285;
    wire N__5284;
    wire N__5281;
    wire N__5278;
    wire N__5275;
    wire N__5272;
    wire N__5267;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5243;
    wire N__5240;
    wire N__5237;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5222;
    wire N__5219;
    wire N__5216;
    wire N__5213;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5198;
    wire N__5195;
    wire N__5192;
    wire N__5189;
    wire N__5186;
    wire N__5183;
    wire N__5180;
    wire N__5177;
    wire N__5174;
    wire N__5171;
    wire N__5168;
    wire N__5165;
    wire N__5162;
    wire N__5159;
    wire N__5156;
    wire N__5153;
    wire N__5150;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5137;
    wire N__5134;
    wire N__5131;
    wire N__5128;
    wire N__5125;
    wire N__5122;
    wire N__5119;
    wire N__5116;
    wire N__5113;
    wire N__5110;
    wire N__5107;
    wire N__5104;
    wire N__5099;
    wire N__5096;
    wire N__5093;
    wire N__5090;
    wire N__5087;
    wire N__5084;
    wire N__5081;
    wire N__5078;
    wire N__5075;
    wire N__5072;
    wire N__5069;
    wire N__5066;
    wire N__5063;
    wire N__5060;
    wire N__5057;
    wire N__5054;
    wire N__5051;
    wire N__5048;
    wire N__5045;
    wire N__5042;
    wire N__5039;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5027;
    wire N__5024;
    wire N__5021;
    wire N__5018;
    wire N__5015;
    wire N__5012;
    wire N__5009;
    wire N__5006;
    wire N__5003;
    wire N__5000;
    wire N__4997;
    wire N__4994;
    wire N__4991;
    wire N__4988;
    wire N__4985;
    wire N__4982;
    wire N__4979;
    wire N__4976;
    wire N__4973;
    wire N__4970;
    wire N__4967;
    wire N__4964;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4943;
    wire N__4940;
    wire N__4937;
    wire N__4934;
    wire N__4931;
    wire N__4928;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4916;
    wire N__4913;
    wire N__4910;
    wire N__4907;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4895;
    wire N__4892;
    wire N__4889;
    wire N__4886;
    wire N__4883;
    wire N__4880;
    wire N__4877;
    wire N__4874;
    wire N__4871;
    wire N__4868;
    wire N__4865;
    wire N__4862;
    wire N__4859;
    wire N__4856;
    wire N__4853;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4841;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4793;
    wire N__4790;
    wire N__4787;
    wire N__4784;
    wire N__4781;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4745;
    wire N__4742;
    wire N__4739;
    wire N__4736;
    wire N__4733;
    wire N__4730;
    wire N__4727;
    wire N__4724;
    wire N__4721;
    wire N__4718;
    wire N__4715;
    wire N__4712;
    wire N__4709;
    wire N__4706;
    wire N__4703;
    wire N__4700;
    wire N__4697;
    wire N__4694;
    wire N__4691;
    wire N__4688;
    wire N__4685;
    wire N__4682;
    wire N__4679;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4667;
    wire N__4664;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4640;
    wire N__4637;
    wire N__4634;
    wire N__4631;
    wire N__4630;
    wire N__4627;
    wire N__4624;
    wire N__4621;
    wire N__4618;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4586;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4562;
    wire N__4559;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4531;
    wire N__4528;
    wire N__4525;
    wire N__4522;
    wire N__4519;
    wire N__4516;
    wire N__4513;
    wire N__4510;
    wire N__4507;
    wire N__4504;
    wire N__4501;
    wire N__4498;
    wire N__4495;
    wire N__4492;
    wire N__4489;
    wire N__4484;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4463;
    wire N__4460;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4445;
    wire N__4442;
    wire N__4439;
    wire N__4436;
    wire N__4433;
    wire N__4430;
    wire N__4427;
    wire N__4424;
    wire N__4421;
    wire N__4418;
    wire N__4415;
    wire N__4412;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4402;
    wire N__4399;
    wire N__4396;
    wire N__4393;
    wire N__4390;
    wire N__4387;
    wire N__4384;
    wire N__4381;
    wire N__4378;
    wire N__4375;
    wire N__4372;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4343;
    wire N__4340;
    wire N__4337;
    wire N__4334;
    wire N__4331;
    wire N__4328;
    wire N__4325;
    wire N__4322;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4310;
    wire N__4307;
    wire N__4304;
    wire N__4301;
    wire N__4298;
    wire N__4295;
    wire N__4292;
    wire N__4289;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4277;
    wire N__4274;
    wire N__4271;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4238;
    wire N__4235;
    wire N__4232;
    wire N__4229;
    wire N__4226;
    wire N__4223;
    wire N__4220;
    wire N__4217;
    wire N__4214;
    wire N__4211;
    wire N__4208;
    wire N__4205;
    wire N__4202;
    wire N__4199;
    wire N__4196;
    wire N__4193;
    wire N__4190;
    wire N__4187;
    wire N__4184;
    wire N__4181;
    wire N__4178;
    wire N__4175;
    wire N__4172;
    wire N__4169;
    wire N__4166;
    wire N__4163;
    wire N__4160;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4148;
    wire N__4145;
    wire N__4142;
    wire N__4139;
    wire N__4136;
    wire N__4133;
    wire N__4130;
    wire N__4127;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4112;
    wire N__4109;
    wire N__4106;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4082;
    wire N__4079;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4067;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4052;
    wire N__4049;
    wire N__4046;
    wire N__4043;
    wire N__4040;
    wire N__4037;
    wire TCIn_c;
    wire VCCG0;
    wire GNDG0;
    wire TAn_in;
    wire N_267_i;
    wire RESETn_c_i;
    wire N_266_i;
    wire \U111_CYCLE_SM.CYCLE_STATE_0_0 ;
    wire N_247_i;
    wire N_249_i;
    wire N_251_i;
    wire N_253_i;
    wire N_254_i;
    wire N_252_i;
    wire U111_CYCLE_SM_A_AMIGA_0_i_1;
    wire A_040_c_0;
    wire A_AMIGA_c_0;
    wire N_264_i;
    wire N_262_i;
    wire N_258_i;
    wire N_246_i;
    wire N_248_i;
    wire D_LL_AMIGA_in_5;
    wire un2_D_LL_AMIGA_5;
    wire A_040_c_1;
    wire D_LM_AMIGA_in_6;
    wire un2_D_LM_AMIGA_6;
    wire N_242_i;
    wire N_260_i;
    wire D_LL_040_in_3;
    wire D_UM_040_in_3;
    wire un1_D_UM_040_3;
    wire N_239_i;
    wire D_UU_040_in_6;
    wire D_LM_040_in_6;
    wire un1_D_UU_040_6;
    wire N_263_i;
    wire N_265_i;
    wire N_257_i;
    wire D_LM_AMIGA_in_5;
    wire un2_D_LM_AMIGA_5;
    wire N_250_i;
    wire D_LM_AMIGA_in_7;
    wire un2_D_LM_AMIGA_7;
    wire N_238_i;
    wire N_241_i;
    wire N_261_i;
    wire N_256_i;
    wire D_LM_AMIGA_in_2;
    wire un2_D_LM_AMIGA_2;
    wire N_245_i;
    wire D_LM_AMIGA_in_4;
    wire un2_D_LM_AMIGA_4;
    wire WRITE_CYCLE_ACTIVE_rep16_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep20_i_ess;
    wire N_259_i;
    wire N_240_i;
    wire N_243_i;
    wire N_237_i;
    wire D_LM_040_in_0;
    wire D_UU_040_in_0;
    wire un1_D_UU_040_0;
    wire CONSTANT_ONE_NET;
    wire D_LL_AMIGA_in_6;
    wire un2_D_LL_AMIGA_6;
    wire D_LM_AMIGA_in_1;
    wire un2_D_LM_AMIGA_1;
    wire D_LM_AMIGA_in_3;
    wire un2_D_LM_AMIGA_3;
    wire LBENn_c_i;
    wire D_LM_040_in_2;
    wire D_UU_040_in_2;
    wire un1_D_UU_040_2;
    wire D_LM_AMIGA_in_0;
    wire un2_D_LM_AMIGA_0;
    wire N_268_i;
    wire N_255_i;
    wire TSn_c;
    wire \INVU111_CYCLE_SM.TSnC_net ;
    wire WRITE_CYCLE_ACTIVE_rep17_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep19_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep8_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep25_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep27_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep28_i_ess;
    wire WRITE_CYCLE_ACTIVE_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep18_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep10_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep26_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep22_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep0_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep21_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep2_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep14_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep1_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep23_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep29_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep3_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep4_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep12_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep7_i_ess;
    wire N_244_i;
    wire D_LM_040_in_5;
    wire D_UU_040_in_5;
    wire un1_D_UU_040_5;
    wire D_LM_040_in_3;
    wire D_UU_040_in_3;
    wire un1_D_UU_040_3;
    wire D_LL_AMIGA_in_3;
    wire un2_D_LL_AMIGA_3;
    wire WRITE_CYCLE_ACTIVE_rep30_i_ess;
    wire GB_BUFFER_CLK40_THRU_CO;
    wire WRITE_CYCLE_ACTIVE_rep24_i_ess;
    wire \U111_CYCLE_SM.A2_ENZ0 ;
    wire \U111_CYCLE_SM.N_67 ;
    wire \U111_CYCLE_SM.TS_ENZ0 ;
    wire TS_CPUn_c;
    wire BGn_c;
    wire \U111_CYCLE_SM.TS_DELAYZ0 ;
    wire WRITE_CYCLE_ACTIVE_rep11_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep5_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep15_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep9_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep13_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep6_i_ess;
    wire LBENn_c_i_0;
    wire \U111_CYCLE_SM.N_33 ;
    wire \U111_CYCLE_SM.N_49 ;
    wire \U111_CYCLE_SM.N_75 ;
    wire \U111_CYCLE_SM.N_75_cascade_ ;
    wire \U111_CYCLE_SM.LATCH_EN_5 ;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa_cascade_ ;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ;
    wire SIZ_c_1;
    wire SIZ_c_0;
    wire READ_CYCLE_ACTIVE_rep6_i_ess;
    wire N_211_i;
    wire READ_CYCLE_ACTIVE_rep2_i_ess;
    wire N_207_i;
    wire D_LL_AMIGA_in_0;
    wire un2_D_LL_AMIGA_0;
    wire D_LL_AMIGA_in_2;
    wire un2_D_LL_AMIGA_2;
    wire READ_CYCLE_ACTIVE_rep26_i_ess;
    wire N_231_i;
    wire D_LL_AMIGA_in_7;
    wire un2_D_LL_AMIGA_7;
    wire \U111_CYCLE_SM.LW_TRANSZ0 ;
    wire PORTSIZE_c;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ;
    wire \U111_CYCLE_SM.N_60_cascade_ ;
    wire \U111_CYCLE_SM.N_46_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ;
    wire \U111_CYCLE_SM.N_39 ;
    wire \U111_CYCLE_SM.N_40 ;
    wire \U111_CYCLE_SM.N_40_cascade_ ;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81_cascade_ ;
    wire TEAn_c;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ;
    wire RESETn_c;
    wire \U111_CYCLE_SM.N_55_cascade_ ;
    wire \U111_CYCLE_SM.N_73 ;
    wire \U111_CYCLE_SM.PORT_MISMATCHZ0 ;
    wire TACKn_in;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ;
    wire \U111_CYCLE_SM.N_57_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_1_0 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ;
    wire \U111_CYCLE_SM.BURST_COUNTZ0Z_1 ;
    wire \U111_CYCLE_SM.BURSTZ0 ;
    wire TBIn_c;
    wire \U111_CYCLE_SM.BURST_COUNTZ0Z_0 ;
    wire \U111_CYCLE_SM.N_42 ;
    wire CLK80;
    wire GB_BUFFER_CLK80_THRU_CO;
    wire READ_CYCLE_ACTIVE_rep5_i_ess;
    wire N_210_i;
    wire D_UM_040_in_1;
    wire D_LL_040_in_1;
    wire un1_D_UM_040_1;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ;
    wire D_UU_AMIGA_in_1;
    wire un1_D_UU_AMIGA_1;
    wire D_UM_AMIGA_in_3;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ;
    wire un1_D_UM_AMIGA_3;
    wire D_UM_AMIGA_in_5;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ;
    wire un1_D_UM_AMIGA_5;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ;
    wire D_UU_AMIGA_in_2;
    wire un1_D_UU_AMIGA_2;
    wire READ_CYCLE_ACTIVE_rep1_i_ess;
    wire N_206_i;
    wire \U111_CYCLE_SM.TA_DISZ0 ;
    wire LBENn_c;
    wire TAn_1_i;
    wire D_LM_040_in_4;
    wire D_UU_040_in_4;
    wire un1_D_UU_040_4;
    wire D_LL_AMIGA_in_1;
    wire un2_D_LL_AMIGA_1;
    wire D_LL_AMIGA_in_4;
    wire un2_D_LL_AMIGA_4;
    wire D_LL_040_in_0;
    wire D_UM_040_in_0;
    wire un1_D_UM_040_0;
    wire un1_D_UM_AMIGA_2;
    wire D_UM_AMIGA_in_2;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ;
    wire \U111_CYCLE_SM.N_40_i_0 ;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81 ;
    wire D_UU_AMIGA_in_0;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ;
    wire un1_D_UU_AMIGA_0;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ;
    wire D_UU_AMIGA_in_6;
    wire un1_D_UU_AMIGA_6;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ;
    wire D_UU_AMIGA_in_3;
    wire un1_D_UU_AMIGA_3;
    wire D_UM_AMIGA_in_7;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ;
    wire un1_D_UM_AMIGA_7;
    wire D_UU_040_in_7;
    wire D_LM_040_in_7;
    wire un1_D_UU_040_7;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ;
    wire D_UM_AMIGA_in_4;
    wire un1_D_UM_AMIGA_4;
    wire D_UU_AMIGA_in_4;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ;
    wire un1_D_UU_AMIGA_4;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ;
    wire D_UU_AMIGA_in_5;
    wire un1_D_UU_AMIGA_5;
    wire N_224_i;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ;
    wire D_UM_AMIGA_in_0;
    wire un1_D_UM_AMIGA_0;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ;
    wire D_UM_AMIGA_in_6;
    wire un1_D_UM_AMIGA_6;
    wire READ_CYCLE_ACTIVE_rep19_i_ess;
    wire D_UM_AMIGA_in_1;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ;
    wire un1_D_UM_AMIGA_1;
    wire READ_CYCLE_ACTIVE_rep11_i_ess;
    wire N_216_i;
    wire D_LM_040_in_1;
    wire D_UU_040_in_1;
    wire un1_D_UU_040_1;
    wire D_UU_AMIGA_in_7;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ;
    wire \U111_CYCLE_SM.LATCH_ENZ0 ;
    wire un1_D_UU_AMIGA_7;
    wire READ_CYCLE_ACTIVE_rep14_i_ess;
    wire N_219_i;
    wire READ_CYCLE_ACTIVE_rep15_i_ess;
    wire N_220_i;
    wire READ_CYCLE_ACTIVE_rep29_i_ess;
    wire N_234_i;
    wire D_LL_040_in_6;
    wire D_UM_040_in_6;
    wire un1_D_UM_040_6;
    wire RnW_c;
    wire \U111_CYCLE_SM.N_44 ;
    wire CLK40;
    wire \U111_CYCLE_SM.CYCLE_STATE_0_g_0 ;
    wire RESETn_c_i_g;
    wire READ_CYCLE_ACTIVE_rep27_i_ess;
    wire N_232_i;
    wire READ_CYCLE_ACTIVE_rep18_i_ess;
    wire N_223_i;
    wire READ_CYCLE_ACTIVE_rep0_i_ess;
    wire N_205_i;
    wire READ_CYCLE_ACTIVE_rep7_i_ess;
    wire N_212_i;
    wire D_UM_040_in_2;
    wire D_LL_040_in_2;
    wire un1_D_UM_040_2;
    wire READ_CYCLE_ACTIVE_rep31_i_ess;
    wire N_236_i;
    wire READ_CYCLE_ACTIVE_rep22_i_ess;
    wire N_227_i;
    wire READ_CYCLE_ACTIVE_rep13_i_ess;
    wire N_218_i;
    wire READ_CYCLE_ACTIVE_rep4_i_ess;
    wire N_209_i;
    wire D_UM_040_in_7;
    wire D_LL_040_in_7;
    wire un1_D_UM_040_7;
    wire READ_CYCLE_ACTIVE_rep28_i_ess;
    wire N_233_i;
    wire READ_CYCLE_ACTIVE_rep30_i_ess;
    wire N_235_i;
    wire READ_CYCLE_ACTIVE_rep17_i_ess;
    wire N_222_i;
    wire D_UM_040_in_4;
    wire D_LL_040_in_4;
    wire un1_D_UM_040_4;
    wire D_LL_040_in_5;
    wire D_UM_040_in_5;
    wire \U111_CYCLE_SM.FLIP_WORDZ0 ;
    wire un1_D_UM_040_5;
    wire READ_CYCLE_ACTIVE_rep25_i_ess;
    wire N_230_i;
    wire READ_CYCLE_ACTIVE_rep10_i_ess;
    wire N_215_i;
    wire READ_CYCLE_ACTIVE_rep21_i_ess;
    wire N_226_i;
    wire READ_CYCLE_ACTIVE_rep24_i_ess;
    wire N_229_i;
    wire READ_CYCLE_ACTIVE_rep9_i_ess;
    wire N_214_i;
    wire READ_CYCLE_ACTIVE_rep12_i_ess;
    wire N_217_i;
    wire READ_CYCLE_ACTIVE_rep8_i_ess;
    wire N_213_i;
    wire READ_CYCLE_ACTIVE_rep23_i_ess;
    wire N_228_i;
    wire READ_CYCLE_ACTIVE_rep20_i_ess;
    wire N_225_i;
    wire READ_CYCLE_ACTIVE_rep3_i_ess;
    wire N_208_i;
    wire READ_CYCLE_ACTIVE_rep16_i_ess;
    wire N_221_i;
    wire _gnd_net_;

    defparam pll_pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll_pll.TEST_MODE=1'b0;
    defparam pll_pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll_pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll_pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll_pll.FILTER_RANGE=3'b011;
    defparam pll_pll.FEEDBACK_PATH="SIMPLE";
    defparam pll_pll.FDA_RELATIVE=4'b0000;
    defparam pll_pll.FDA_FEEDBACK=4'b0000;
    defparam pll_pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll_pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll_pll.DIVR=4'b0000;
    defparam pll_pll.DIVQ=3'b011;
    defparam pll_pll.DIVF=7'b0001111;
    defparam pll_pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40_2F pll_pll (
            .SCLK(),
            .PLLOUTGLOBALA(CLK80),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALB(CLK40),
            .SDI(),
            .PLLOUTCOREA(),
            .BYPASS(),
            .RESETB(N__5291),
            .PLLOUTCOREB(),
            .LOCK(),
            .SDO(),
            .EXTFEEDBACK(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__12664));
    IO_PAD pll_iopad (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__12664),
            .PACKAGEPIN(CLK40_IN));
    IO_PAD LBENn_ibuf_iopad (
            .OE(N__12648),
            .DIN(N__12647),
            .DOUT(N__12646),
            .PACKAGEPIN(LBENn));
    defparam LBENn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam LBENn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO LBENn_ibuf_preio (
            .PADOEN(N__12648),
            .PADOUT(N__12647),
            .PADIN(N__12646),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(LBENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TAn_iobuf_iopad (
            .OE(N__12639),
            .DIN(N__12638),
            .DOUT(N__12637),
            .PACKAGEPIN(TAn));
    defparam TAn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TAn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TAn_iobuf_preio (
            .PADOEN(N__12639),
            .PADOUT(N__12638),
            .PADIN(N__12637),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7982),
            .DIN0(TAn_in),
            .DOUT0(N__7205),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_1_iopad (
            .OE(N__12630),
            .DIN(N__12629),
            .DOUT(N__12628),
            .PACKAGEPIN(D_LL_AMIGA[1]));
    defparam D_LL_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_1_preio (
            .PADOEN(N__12630),
            .PADOUT(N__12629),
            .PADIN(N__12628),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4238),
            .DIN0(D_LL_AMIGA_in_1),
            .DOUT0(N__7613),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_6_iopad (
            .OE(N__12621),
            .DIN(N__12620),
            .DOUT(N__12619),
            .PACKAGEPIN(D_UU_040[6]));
    defparam D_UU_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_6_preio (
            .PADOEN(N__12621),
            .PADOUT(N__12620),
            .PADIN(N__12619),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6392),
            .DIN0(D_UU_040_in_6),
            .DOUT0(N__8786),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam CPUBGn_obuf_iopad.PULLUP=1'b1;
    IO_PAD CPUBGn_obuf_iopad (
            .OE(N__12612),
            .DIN(N__12611),
            .DOUT(N__12610),
            .PACKAGEPIN(CPUBGn));
    defparam CPUBGn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CPUBGn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CPUBGn_obuf_preio (
            .PADOEN(N__12612),
            .PADOUT(N__12611),
            .PADIN(N__12610),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_3_iopad (
            .OE(N__12603),
            .DIN(N__12602),
            .DOUT(N__12601),
            .PACKAGEPIN(D_UM_AMIGA[3]));
    defparam D_UM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_3_preio (
            .PADOEN(N__12603),
            .PADOUT(N__12602),
            .PADIN(N__12601),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4697),
            .DIN0(D_UM_AMIGA_in_3),
            .DOUT0(N__4463),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_1_iopad (
            .OE(N__12594),
            .DIN(N__12593),
            .DOUT(N__12592),
            .PACKAGEPIN(A_040[1]));
    defparam A_040_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_1_preio (
            .PADOEN(N__12594),
            .PADOUT(N__12593),
            .PADIN(N__12592),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_4_iopad (
            .OE(N__12585),
            .DIN(N__12584),
            .DOUT(N__12583),
            .PACKAGEPIN(D_LM_AMIGA[4]));
    defparam D_LM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_4_preio (
            .PADOEN(N__12585),
            .PADOUT(N__12584),
            .PADIN(N__12583),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4835),
            .DIN0(D_LM_AMIGA_in_4),
            .DOUT0(N__7967),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_7_iopad (
            .OE(N__12576),
            .DIN(N__12575),
            .DOUT(N__12574),
            .PACKAGEPIN(D_LM_040[7]));
    defparam D_LM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_7_preio (
            .PADOEN(N__12576),
            .PADOUT(N__12575),
            .PADIN(N__12574),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__11576),
            .DIN0(D_LM_040_in_7),
            .DOUT0(N__4763),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_obuf_iopad (
            .OE(N__12567),
            .DIN(N__12566),
            .DOUT(N__12565),
            .PACKAGEPIN(CLK40B));
    defparam CLK40B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_obuf_preio (
            .PADOEN(N__12567),
            .PADOUT(N__12566),
            .PADIN(N__12565),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6123),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_1_iopad (
            .OE(N__12558),
            .DIN(N__12557),
            .DOUT(N__12556),
            .PACKAGEPIN(D_UM_040[1]));
    defparam D_UM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_1_preio (
            .PADOEN(N__12558),
            .PADOUT(N__12557),
            .PADIN(N__12556),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__11678),
            .DIN0(D_UM_040_in_1),
            .DOUT0(N__8972),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_ibuf_iopad (
            .OE(N__12549),
            .DIN(N__12548),
            .DOUT(N__12547),
            .PACKAGEPIN(TBIn));
    defparam TBIn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TBIn_ibuf_preio (
            .PADOEN(N__12549),
            .PADOUT(N__12548),
            .PADIN(N__12547),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TBIn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_7_iopad (
            .OE(N__12540),
            .DIN(N__12539),
            .DOUT(N__12538),
            .PACKAGEPIN(D_UU_AMIGA[7]));
    defparam D_UU_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_7_preio (
            .PADOEN(N__12540),
            .PADOUT(N__12539),
            .PADIN(N__12538),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5675),
            .DIN0(D_UU_AMIGA_in_7),
            .DOUT0(N__8561),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFDIR_obuf_iopad (
            .OE(N__12531),
            .DIN(N__12530),
            .DOUT(N__12529),
            .PACKAGEPIN(BUFDIR));
    defparam BUFDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFDIR_obuf_preio (
            .PADOEN(N__12531),
            .PADOUT(N__12530),
            .PADIN(N__12529),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10094),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__12522),
            .DIN(N__12521),
            .DOUT(N__12520),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__12522),
            .PADOUT(N__12521),
            .PADIN(N__12520),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TS_CPUn_ibuf_iopad (
            .OE(N__12513),
            .DIN(N__12512),
            .DOUT(N__12511),
            .PACKAGEPIN(TS_CPUn));
    defparam TS_CPUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TS_CPUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TS_CPUn_ibuf_preio (
            .PADOEN(N__12513),
            .PADOUT(N__12512),
            .PADIN(N__12511),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TS_CPUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_1_iopad (
            .OE(N__12504),
            .DIN(N__12503),
            .DOUT(N__12502),
            .PACKAGEPIN(D_LL_040[1]));
    defparam D_LL_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_1_preio (
            .PADOEN(N__12504),
            .PADOUT(N__12503),
            .PADIN(N__12502),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10835),
            .DIN0(D_LL_040_in_1),
            .DOUT0(N__7877),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_1_iopad (
            .OE(N__12495),
            .DIN(N__12494),
            .DOUT(N__12493),
            .PACKAGEPIN(D_UU_040[1]));
    defparam D_UU_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_1_preio (
            .PADOEN(N__12495),
            .PADOUT(N__12494),
            .PADIN(N__12493),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8096),
            .DIN0(D_UU_040_in_1),
            .DOUT0(N__7514),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_1_iopad (
            .OE(N__12486),
            .DIN(N__12485),
            .DOUT(N__12484),
            .PACKAGEPIN(D_LM_AMIGA[1]));
    defparam D_LM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_1_preio (
            .PADOEN(N__12486),
            .PADOUT(N__12485),
            .PADIN(N__12484),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4331),
            .DIN0(D_LM_AMIGA_in_1),
            .DOUT0(N__8924),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_2_iopad (
            .OE(N__12477),
            .DIN(N__12476),
            .DOUT(N__12475),
            .PACKAGEPIN(D_LM_040[2]));
    defparam D_LM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_2_preio (
            .PADOEN(N__12477),
            .PADOUT(N__12476),
            .PADIN(N__12475),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10751),
            .DIN0(D_LM_040_in_2),
            .DOUT0(N__5018),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TACKn_iobuf_iopad.PULLUP=1'b1;
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__12468),
            .DIN(N__12467),
            .DOUT(N__12466),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__12468),
            .PADOUT(N__12467),
            .PADIN(N__12466),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6248),
            .DIN0(TACKn_in),
            .DOUT0(N__4187),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_2_iopad (
            .OE(N__12459),
            .DIN(N__12458),
            .DOUT(N__12457),
            .PACKAGEPIN(D_UM_040[2]));
    defparam D_UM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_2_preio (
            .PADOEN(N__12459),
            .PADOUT(N__12458),
            .PADIN(N__12457),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10802),
            .DIN0(D_UM_040_in_2),
            .DOUT0(N__7736),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMB_obuf_iopad (
            .OE(N__12450),
            .DIN(N__12449),
            .DOUT(N__12448),
            .PACKAGEPIN(CLKRAMB));
    defparam CLKRAMB_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMB_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMB_obuf_preio (
            .PADOEN(N__12450),
            .PADOUT(N__12449),
            .PADIN(N__12448),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7703),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_2_iopad (
            .OE(N__12441),
            .DIN(N__12440),
            .DOUT(N__12439),
            .PACKAGEPIN(D_LL_AMIGA[2]));
    defparam D_LL_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_2_preio (
            .PADOEN(N__12441),
            .PADOUT(N__12440),
            .PADIN(N__12439),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4874),
            .DIN0(D_LL_AMIGA_in_2),
            .DOUT0(N__10649),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_2_iopad (
            .OE(N__12432),
            .DIN(N__12431),
            .DOUT(N__12430),
            .PACKAGEPIN(D_UU_AMIGA[2]));
    defparam D_UU_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_2_preio (
            .PADOEN(N__12432),
            .PADOUT(N__12431),
            .PADIN(N__12430),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4445),
            .DIN0(D_UU_AMIGA_in_2),
            .DOUT0(N__5075),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TEAn_ibuf_iopad.PULLUP=1'b1;
    IO_PAD TEAn_ibuf_iopad (
            .OE(N__12423),
            .DIN(N__12422),
            .DOUT(N__12421),
            .PACKAGEPIN(TEAn));
    defparam TEAn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TEAn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TEAn_ibuf_preio (
            .PADOEN(N__12423),
            .PADOUT(N__12422),
            .PADIN(N__12421),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TEAn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__12414),
            .DIN(N__12413),
            .DOUT(N__12412),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__12414),
            .PADOUT(N__12413),
            .PADIN(N__12412),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5159),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMAn_obuf_iopad (
            .OE(N__12405),
            .DIN(N__12404),
            .DOUT(N__12403),
            .PACKAGEPIN(DMAn));
    defparam DMAn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMAn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMAn_obuf_preio (
            .PADOEN(N__12405),
            .PADOUT(N__12404),
            .PADIN(N__12403),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5284),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_6_iopad (
            .OE(N__12396),
            .DIN(N__12395),
            .DOUT(N__12394),
            .PACKAGEPIN(D_LL_040[6]));
    defparam D_LL_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_6_preio (
            .PADOEN(N__12396),
            .PADOUT(N__12395),
            .PADIN(N__12394),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__11369),
            .DIN0(D_LL_040_in_6),
            .DOUT0(N__5249),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_5_iopad (
            .OE(N__12387),
            .DIN(N__12386),
            .DOUT(N__12385),
            .PACKAGEPIN(D_LL_AMIGA[5]));
    defparam D_LL_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_5_preio (
            .PADOEN(N__12387),
            .PADOUT(N__12386),
            .PADIN(N__12385),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4139),
            .DIN0(D_LL_AMIGA_in_5),
            .DOUT0(N__11234),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_0_iopad (
            .OE(N__12378),
            .DIN(N__12377),
            .DOUT(N__12376),
            .PACKAGEPIN(D_UM_AMIGA[0]));
    defparam D_UM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_0_preio (
            .PADOEN(N__12378),
            .PADOUT(N__12377),
            .PADIN(N__12376),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4997),
            .DIN0(D_UM_AMIGA_in_0),
            .DOUT0(N__7760),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_2_iopad (
            .OE(N__12369),
            .DIN(N__12368),
            .DOUT(N__12367),
            .PACKAGEPIN(D_UU_040[2]));
    defparam D_UU_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_2_preio (
            .PADOEN(N__12369),
            .PADOUT(N__12368),
            .PADIN(N__12367),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6665),
            .DIN0(D_UU_040_in_2),
            .DOUT0(N__7280),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_2_iopad (
            .OE(N__12360),
            .DIN(N__12359),
            .DOUT(N__12358),
            .PACKAGEPIN(D_LM_AMIGA[2]));
    defparam D_LM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_2_preio (
            .PADOEN(N__12360),
            .PADOUT(N__12359),
            .PADIN(N__12358),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5495),
            .DIN0(D_LM_AMIGA_in_2),
            .DOUT0(N__5137),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK80_CPU_obuf_iopad (
            .OE(N__12351),
            .DIN(N__12350),
            .DOUT(N__12349),
            .PACKAGEPIN(CLK80_CPU));
    defparam CLK80_CPU_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK80_CPU_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK80_CPU_obuf_preio (
            .PADOEN(N__12351),
            .PADOUT(N__12350),
            .PADIN(N__12349),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7699),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_3_iopad (
            .OE(N__12342),
            .DIN(N__12341),
            .DOUT(N__12340),
            .PACKAGEPIN(D_LL_040[3]));
    defparam D_LL_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_3_preio (
            .PADOEN(N__12342),
            .PADOUT(N__12341),
            .PADIN(N__12340),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10781),
            .DIN0(D_LL_040_in_3),
            .DOUT0(N__5810),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_1_iopad (
            .OE(N__12333),
            .DIN(N__12332),
            .DOUT(N__12331),
            .PACKAGEPIN(D_LM_040[1]));
    defparam D_LM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_1_preio (
            .PADOEN(N__12333),
            .PADOUT(N__12332),
            .PADIN(N__12331),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__11333),
            .DIN0(D_LM_040_in_1),
            .DOUT0(N__5216),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_obuf_iopad (
            .OE(N__12324),
            .DIN(N__12323),
            .DOUT(N__12322),
            .PACKAGEPIN(TSn));
    defparam TSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TSn_obuf_preio (
            .PADOEN(N__12324),
            .PADOUT(N__12323),
            .PADIN(N__12322),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5483),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_7_iopad (
            .OE(N__12315),
            .DIN(N__12314),
            .DOUT(N__12313),
            .PACKAGEPIN(D_UM_AMIGA[7]));
    defparam D_UM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_7_preio (
            .PADOEN(N__12315),
            .PADOUT(N__12314),
            .PADIN(N__12313),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4313),
            .DIN0(D_UM_AMIGA_in_7),
            .DOUT0(N__11435),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_7_iopad (
            .OE(N__12306),
            .DIN(N__12305),
            .DOUT(N__12304),
            .PACKAGEPIN(D_LM_AMIGA[7]));
    defparam D_LM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_7_preio (
            .PADOEN(N__12306),
            .PADOUT(N__12305),
            .PADIN(N__12304),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4553),
            .DIN0(D_LM_AMIGA_in_7),
            .DOUT0(N__8603),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORTSIZE_ibuf_iopad (
            .OE(N__12297),
            .DIN(N__12296),
            .DOUT(N__12295),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO PORTSIZE_ibuf_preio (
            .PADOEN(N__12297),
            .PADOUT(N__12296),
            .PADIN(N__12295),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(PORTSIZE_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_0_iopad (
            .OE(N__12288),
            .DIN(N__12287),
            .DOUT(N__12286),
            .PACKAGEPIN(A_AMIGA[0]));
    defparam A_AMIGA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_0_preio (
            .PADOEN(N__12288),
            .PADOUT(N__12287),
            .PADIN(N__12286),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4271),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_4_iopad (
            .OE(N__12279),
            .DIN(N__12278),
            .DOUT(N__12277),
            .PACKAGEPIN(D_LM_040[4]));
    defparam D_LM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_4_preio (
            .PADOEN(N__12279),
            .PADOUT(N__12278),
            .PADIN(N__12277),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__11549),
            .DIN0(D_LM_040_in_4),
            .DOUT0(N__4970),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_7_iopad (
            .OE(N__12270),
            .DIN(N__12269),
            .DOUT(N__12268),
            .PACKAGEPIN(D_UM_040[7]));
    defparam D_UM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_7_preio (
            .PADOEN(N__12270),
            .PADOUT(N__12269),
            .PADIN(N__12268),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10229),
            .DIN0(D_UM_040_in_7),
            .DOUT0(N__8633),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__12261),
            .DIN(N__12260),
            .DOUT(N__12259),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__12261),
            .PADOUT(N__12260),
            .PADIN(N__12259),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_1_iopad (
            .OE(N__12252),
            .DIN(N__12251),
            .DOUT(N__12250),
            .PACKAGEPIN(D_UU_AMIGA[1]));
    defparam D_UU_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_1_preio (
            .PADOEN(N__12252),
            .PADOUT(N__12251),
            .PADIN(N__12250),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4742),
            .DIN0(D_UU_AMIGA_in_1),
            .DOUT0(N__8858),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_obuf_iopad (
            .OE(N__12243),
            .DIN(N__12242),
            .DOUT(N__12241),
            .PACKAGEPIN(CLK40C));
    defparam CLK40C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_obuf_preio (
            .PADOEN(N__12243),
            .PADOUT(N__12242),
            .PADIN(N__12241),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6122),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_0_iopad (
            .OE(N__12234),
            .DIN(N__12233),
            .DOUT(N__12232),
            .PACKAGEPIN(D_UM_040[0]));
    defparam D_UM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_0_preio (
            .PADOEN(N__12234),
            .PADOUT(N__12233),
            .PADIN(N__12232),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__11606),
            .DIN0(D_UM_040_in_0),
            .DOUT0(N__9122),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_0_iopad (
            .OE(N__12225),
            .DIN(N__12224),
            .DOUT(N__12223),
            .PACKAGEPIN(D_LL_AMIGA[0]));
    defparam D_LL_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_0_preio (
            .PADOEN(N__12225),
            .PADOUT(N__12224),
            .PADIN(N__12223),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4709),
            .DIN0(D_LL_AMIGA_in_0),
            .DOUT0(N__7817),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_4_iopad (
            .OE(N__12216),
            .DIN(N__12215),
            .DOUT(N__12214),
            .PACKAGEPIN(D_UU_AMIGA[4]));
    defparam D_UU_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_4_preio (
            .PADOEN(N__12216),
            .PADOUT(N__12215),
            .PADIN(N__12214),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4724),
            .DIN0(D_UU_AMIGA_in_4),
            .DOUT0(N__7913),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_7_iopad (
            .OE(N__12207),
            .DIN(N__12206),
            .DOUT(N__12205),
            .PACKAGEPIN(D_UU_040[7]));
    defparam D_UU_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_7_preio (
            .PADOEN(N__12207),
            .PADOUT(N__12206),
            .PADIN(N__12205),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10679),
            .DIN0(D_UU_040_in_7),
            .DOUT0(N__10289),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__12198),
            .DIN(N__12197),
            .DOUT(N__12196),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__12198),
            .PADOUT(N__12197),
            .PADIN(N__12196),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam BGn_ibuf_iopad.PULLUP=1'b1;
    IO_PAD BGn_ibuf_iopad (
            .OE(N__12189),
            .DIN(N__12188),
            .DOUT(N__12187),
            .PACKAGEPIN(BGn));
    defparam BGn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BGn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BGn_ibuf_preio (
            .PADOEN(N__12189),
            .PADOUT(N__12188),
            .PADIN(N__12187),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(BGn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_0_iopad (
            .OE(N__12180),
            .DIN(N__12179),
            .DOUT(N__12178),
            .PACKAGEPIN(D_LL_040[0]));
    defparam D_LL_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_0_preio (
            .PADOEN(N__12180),
            .PADOUT(N__12179),
            .PADIN(N__12178),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__11714),
            .DIN0(D_LL_040_in_0),
            .DOUT0(N__6632),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_2_iopad (
            .OE(N__12171),
            .DIN(N__12170),
            .DOUT(N__12169),
            .PACKAGEPIN(D_UM_AMIGA[2]));
    defparam D_UM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_2_preio (
            .PADOEN(N__12171),
            .PADOUT(N__12170),
            .PADIN(N__12169),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4112),
            .DIN0(D_UM_AMIGA_in_2),
            .DOUT0(N__10610),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_0_iopad (
            .OE(N__12162),
            .DIN(N__12161),
            .DOUT(N__12160),
            .PACKAGEPIN(D_UU_040[0]));
    defparam D_UU_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_0_preio (
            .PADOEN(N__12162),
            .PADOUT(N__12161),
            .PADIN(N__12160),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10715),
            .DIN0(D_UU_040_in_0),
            .DOUT0(N__8117),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_ibuf_iopad (
            .OE(N__12153),
            .DIN(N__12152),
            .DOUT(N__12151),
            .PACKAGEPIN(TCIn));
    defparam TCIn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TCIn_ibuf_preio (
            .PADOEN(N__12153),
            .PADOUT(N__12152),
            .PADIN(N__12151),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TCIn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_0_iopad (
            .OE(N__12144),
            .DIN(N__12143),
            .DOUT(N__12142),
            .PACKAGEPIN(A_040[0]));
    defparam A_040_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_0_preio (
            .PADOEN(N__12144),
            .PADOUT(N__12143),
            .PADIN(N__12142),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_0_iopad (
            .OE(N__12135),
            .DIN(N__12134),
            .DOUT(N__12133),
            .PACKAGEPIN(D_LM_AMIGA[0]));
    defparam D_LM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_0_preio (
            .PADOEN(N__12135),
            .PADOUT(N__12134),
            .PADIN(N__12133),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4349),
            .DIN0(D_LM_AMIGA_in_0),
            .DOUT0(N__5381),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBI_CPUn_obuf_iopad (
            .OE(N__12126),
            .DIN(N__12125),
            .DOUT(N__12124),
            .PACKAGEPIN(TBI_CPUn));
    defparam TBI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TBI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TBI_CPUn_obuf_preio (
            .PADOEN(N__12126),
            .PADOUT(N__12125),
            .PADIN(N__12124),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7003),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40A_obuf_iopad (
            .OE(N__12117),
            .DIN(N__12116),
            .DOUT(N__12115),
            .PACKAGEPIN(CLK40A));
    defparam CLK40A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40A_obuf_preio (
            .PADOEN(N__12117),
            .PADOUT(N__12116),
            .PADIN(N__12115),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6133),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_3_iopad (
            .OE(N__12108),
            .DIN(N__12107),
            .DOUT(N__12106),
            .PACKAGEPIN(D_LM_040[3]));
    defparam D_LM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_3_preio (
            .PADOEN(N__12108),
            .PADOUT(N__12107),
            .PADIN(N__12106),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8300),
            .DIN0(D_LM_040_in_3),
            .DOUT0(N__5183),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_5_iopad (
            .OE(N__12099),
            .DIN(N__12098),
            .DOUT(N__12097),
            .PACKAGEPIN(D_LM_AMIGA[5]));
    defparam D_LM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_5_preio (
            .PADOEN(N__12099),
            .PADOUT(N__12098),
            .PADIN(N__12097),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4217),
            .DIN0(D_LM_AMIGA_in_5),
            .DOUT0(N__5996),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_6_iopad (
            .OE(N__12090),
            .DIN(N__12089),
            .DOUT(N__12088),
            .PACKAGEPIN(D_LM_040[6]));
    defparam D_LM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_6_preio (
            .PADOEN(N__12090),
            .PADOUT(N__12089),
            .PADIN(N__12088),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10556),
            .DIN0(D_LM_040_in_6),
            .DOUT0(N__4595),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_5_iopad (
            .OE(N__12081),
            .DIN(N__12080),
            .DOUT(N__12079),
            .PACKAGEPIN(D_UM_040[5]));
    defparam D_UM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_5_preio (
            .PADOEN(N__12081),
            .PADOUT(N__12080),
            .PADIN(N__12079),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10523),
            .DIN0(D_UM_040_in_5),
            .DOUT0(N__7352),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_3_iopad (
            .OE(N__12072),
            .DIN(N__12071),
            .DOUT(N__12070),
            .PACKAGEPIN(D_LL_AMIGA[3]));
    defparam D_LL_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_3_preio (
            .PADOEN(N__12072),
            .PADOUT(N__12071),
            .PADIN(N__12070),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4256),
            .DIN0(D_LL_AMIGA_in_3),
            .DOUT0(N__4531),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_3_iopad (
            .OE(N__12063),
            .DIN(N__12062),
            .DOUT(N__12061),
            .PACKAGEPIN(D_UU_AMIGA[3]));
    defparam D_UU_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_3_preio (
            .PADOEN(N__12063),
            .PADOUT(N__12062),
            .PADIN(N__12061),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4907),
            .DIN0(D_UU_AMIGA_in_3),
            .DOUT0(N__5846),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_5_iopad (
            .OE(N__12054),
            .DIN(N__12053),
            .DOUT(N__12052),
            .PACKAGEPIN(D_LL_040[5]));
    defparam D_LL_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_5_preio (
            .PADOEN(N__12054),
            .PADOUT(N__12053),
            .PADIN(N__12052),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10196),
            .DIN0(D_LL_040_in_5),
            .DOUT0(N__4664),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_6_iopad (
            .OE(N__12045),
            .DIN(N__12044),
            .DOUT(N__12043),
            .PACKAGEPIN(D_LL_AMIGA[6]));
    defparam D_LL_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_6_preio (
            .PADOEN(N__12045),
            .PADOUT(N__12044),
            .PADIN(N__12043),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4163),
            .DIN0(D_LL_AMIGA_in_6),
            .DOUT0(N__10181),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_6_iopad (
            .OE(N__12036),
            .DIN(N__12035),
            .DOUT(N__12034),
            .PACKAGEPIN(D_UU_AMIGA[6]));
    defparam D_UU_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_6_preio (
            .PADOEN(N__12036),
            .PADOUT(N__12035),
            .PADIN(N__12034),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4886),
            .DIN0(D_UU_AMIGA_in_6),
            .DOUT0(N__4367),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_1_iopad (
            .OE(N__12027),
            .DIN(N__12026),
            .DOUT(N__12025),
            .PACKAGEPIN(D_UM_AMIGA[1]));
    defparam D_UM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_1_preio (
            .PADOEN(N__12027),
            .PADOUT(N__12026),
            .PADIN(N__12025),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4202),
            .DIN0(D_UM_AMIGA_in_1),
            .DOUT0(N__7577),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_5_iopad (
            .OE(N__12018),
            .DIN(N__12017),
            .DOUT(N__12016),
            .PACKAGEPIN(D_UU_040[5]));
    defparam D_UU_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_5_preio (
            .PADOEN(N__12018),
            .PADOUT(N__12017),
            .PADIN(N__12016),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7655),
            .DIN0(D_UU_040_in_5),
            .DOUT0(N__8321),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMA_obuf_iopad (
            .OE(N__12009),
            .DIN(N__12008),
            .DOUT(N__12007),
            .PACKAGEPIN(CLKRAMA));
    defparam CLKRAMA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMA_obuf_preio (
            .PADOEN(N__12009),
            .PADOUT(N__12008),
            .PADIN(N__12007),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6134),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_2_iopad (
            .OE(N__12000),
            .DIN(N__11999),
            .DOUT(N__11998),
            .PACKAGEPIN(D_LL_040[2]));
    defparam D_LL_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_2_preio (
            .PADOEN(N__12000),
            .PADOUT(N__11999),
            .PADIN(N__11998),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6557),
            .DIN0(D_LL_040_in_2),
            .DOUT0(N__6593),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCI_CPUn_obuf_iopad (
            .OE(N__11991),
            .DIN(N__11990),
            .DOUT(N__11989),
            .PACKAGEPIN(TCI_CPUn));
    defparam TCI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TCI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TCI_CPUn_obuf_preio (
            .PADOEN(N__11991),
            .PADOUT(N__11990),
            .PADIN(N__11989),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4064),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_4_iopad (
            .OE(N__11982),
            .DIN(N__11981),
            .DOUT(N__11980),
            .PACKAGEPIN(D_UM_AMIGA[4]));
    defparam D_UM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_4_preio (
            .PADOEN(N__11982),
            .PADOUT(N__11981),
            .PADIN(N__11980),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4100),
            .DIN0(D_UM_AMIGA_in_4),
            .DOUT0(N__11255),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_6_iopad (
            .OE(N__11973),
            .DIN(N__11972),
            .DOUT(N__11971),
            .PACKAGEPIN(D_LM_AMIGA[6]));
    defparam D_LM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_6_preio (
            .PADOEN(N__11973),
            .PADOUT(N__11972),
            .PADIN(N__11971),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4928),
            .DIN0(D_LM_AMIGA_in_6),
            .DOUT0(N__4409),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__11964),
            .DIN(N__11963),
            .DOUT(N__11962),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__11964),
            .PADOUT(N__11963),
            .PADIN(N__11962),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_5_iopad (
            .OE(N__11955),
            .DIN(N__11954),
            .DOUT(N__11953),
            .PACKAGEPIN(D_LM_040[5]));
    defparam D_LM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_5_preio (
            .PADOEN(N__11955),
            .PADOUT(N__11954),
            .PADIN(N__11953),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__11738),
            .DIN0(D_LM_040_in_5),
            .DOUT0(N__4808),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_6_iopad (
            .OE(N__11946),
            .DIN(N__11945),
            .DOUT(N__11944),
            .PACKAGEPIN(D_UM_040[6]));
    defparam D_UM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_6_preio (
            .PADOEN(N__11946),
            .PADOUT(N__11945),
            .PADIN(N__11944),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10259),
            .DIN0(D_UM_040_in_6),
            .DOUT0(N__9050),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_3_iopad (
            .OE(N__11937),
            .DIN(N__11936),
            .DOUT(N__11935),
            .PACKAGEPIN(D_UM_040[3]));
    defparam D_UM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_3_preio (
            .PADOEN(N__11937),
            .PADOUT(N__11936),
            .PADIN(N__11935),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8939),
            .DIN0(D_UM_040_in_3),
            .DOUT0(N__7433),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_5_iopad (
            .OE(N__11928),
            .DIN(N__11927),
            .DOUT(N__11926),
            .PACKAGEPIN(D_UU_AMIGA[5]));
    defparam D_UU_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_5_preio (
            .PADOEN(N__11928),
            .PADOUT(N__11927),
            .PADIN(N__11926),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4574),
            .DIN0(D_UU_AMIGA_in_5),
            .DOUT0(N__5930),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_7_iopad (
            .OE(N__11919),
            .DIN(N__11918),
            .DOUT(N__11917),
            .PACKAGEPIN(D_LL_040[7]));
    defparam D_LL_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_7_preio (
            .PADOEN(N__11919),
            .PADOUT(N__11918),
            .PADIN(N__11917),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10580),
            .DIN0(D_LL_040_in_7),
            .DOUT0(N__6527),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_4_iopad (
            .OE(N__11910),
            .DIN(N__11909),
            .DOUT(N__11908),
            .PACKAGEPIN(D_LL_AMIGA[4]));
    defparam D_LL_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_4_preio (
            .PADOEN(N__11910),
            .PADOUT(N__11909),
            .PADIN(N__11908),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4856),
            .DIN0(D_LL_AMIGA_in_4),
            .DOUT0(N__11303),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_3_iopad (
            .OE(N__11901),
            .DIN(N__11900),
            .DOUT(N__11899),
            .PACKAGEPIN(D_UU_040[3]));
    defparam D_UU_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_3_preio (
            .PADOEN(N__11901),
            .PADOUT(N__11900),
            .PADIN(N__11899),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__11516),
            .DIN0(D_UU_040_in_3),
            .DOUT0(N__8711),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TEA_CPUn_obuf_iopad (
            .OE(N__11892),
            .DIN(N__11891),
            .DOUT(N__11890),
            .PACKAGEPIN(TEA_CPUn));
    defparam TEA_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TEA_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TEA_CPUn_obuf_preio (
            .PADOEN(N__11892),
            .PADOUT(N__11891),
            .PADIN(N__11890),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6851),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_3_iopad (
            .OE(N__11883),
            .DIN(N__11882),
            .DOUT(N__11881),
            .PACKAGEPIN(D_LM_AMIGA[3]));
    defparam D_LM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_3_preio (
            .PADOEN(N__11883),
            .PADOUT(N__11882),
            .PADIN(N__11881),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5039),
            .DIN0(D_LM_AMIGA_in_3),
            .DOUT0(N__5909),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_0_iopad (
            .OE(N__11874),
            .DIN(N__11873),
            .DOUT(N__11872),
            .PACKAGEPIN(D_LM_040[0]));
    defparam D_LM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_0_preio (
            .PADOEN(N__11874),
            .PADOUT(N__11873),
            .PADIN(N__11872),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__11765),
            .DIN0(D_LM_040_in_0),
            .DOUT0(N__5537),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_6_iopad (
            .OE(N__11865),
            .DIN(N__11864),
            .DOUT(N__11863),
            .PACKAGEPIN(D_UM_AMIGA[6]));
    defparam D_UM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_6_preio (
            .PADOEN(N__11865),
            .PADOUT(N__11864),
            .PADIN(N__11863),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4082),
            .DIN0(D_UM_AMIGA_in_6),
            .DOUT0(N__10118),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_1_iopad (
            .OE(N__11856),
            .DIN(N__11855),
            .DOUT(N__11854),
            .PACKAGEPIN(A_AMIGA[1]));
    defparam A_AMIGA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_1_preio (
            .PADOEN(N__11856),
            .PADOUT(N__11855),
            .PADIN(N__11854),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4295),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_4_iopad (
            .OE(N__11847),
            .DIN(N__11846),
            .DOUT(N__11845),
            .PACKAGEPIN(D_UM_040[4]));
    defparam D_UM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_4_preio (
            .PADOEN(N__11847),
            .PADOUT(N__11846),
            .PADIN(N__11845),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__11642),
            .DIN0(D_UM_040_in_4),
            .DOUT0(N__8480),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_0_iopad (
            .OE(N__11838),
            .DIN(N__11837),
            .DOUT(N__11836),
            .PACKAGEPIN(D_UU_AMIGA[0]));
    defparam D_UU_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_0_preio (
            .PADOEN(N__11838),
            .PADOUT(N__11837),
            .PADIN(N__11836),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5399),
            .DIN0(D_UU_AMIGA_in_0),
            .DOUT0(N__5309),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_4_iopad (
            .OE(N__11829),
            .DIN(N__11828),
            .DOUT(N__11827),
            .PACKAGEPIN(D_LL_040[4]));
    defparam D_LL_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_4_preio (
            .PADOEN(N__11829),
            .PADOUT(N__11828),
            .PADIN(N__11827),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__11402),
            .DIN0(D_LL_040_in_4),
            .DOUT0(N__7838),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_7_iopad (
            .OE(N__11820),
            .DIN(N__11819),
            .DOUT(N__11818),
            .PACKAGEPIN(D_LL_AMIGA[7]));
    defparam D_LL_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_7_preio (
            .PADOEN(N__11820),
            .PADOUT(N__11819),
            .PADIN(N__11818),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5516),
            .DIN0(D_LL_AMIGA_in_7),
            .DOUT0(N__11486),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_4_iopad (
            .OE(N__11811),
            .DIN(N__11810),
            .DOUT(N__11809),
            .PACKAGEPIN(D_UU_040[4]));
    defparam D_UU_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_4_preio (
            .PADOEN(N__11811),
            .PADOUT(N__11810),
            .PADIN(N__11809),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10490),
            .DIN0(D_UU_040_in_4),
            .DOUT0(N__8399),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_5_iopad (
            .OE(N__11802),
            .DIN(N__11801),
            .DOUT(N__11800),
            .PACKAGEPIN(D_UM_AMIGA[5]));
    defparam D_UM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_5_preio (
            .PADOEN(N__11802),
            .PADOUT(N__11801),
            .PADIN(N__11800),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4793),
            .DIN0(D_UM_AMIGA_in_5),
            .DOUT0(N__10865),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2923 (
            .O(N__11783),
            .I(N__11780));
    LocalMux I__2922 (
            .O(N__11780),
            .I(N__11777));
    Span4Mux_v I__2921 (
            .O(N__11777),
            .I(N__11774));
    Sp12to4 I__2920 (
            .O(N__11774),
            .I(N__11771));
    Span12Mux_h I__2919 (
            .O(N__11771),
            .I(N__11768));
    Odrv12 I__2918 (
            .O(N__11768),
            .I(READ_CYCLE_ACTIVE_rep16_i_ess));
    IoInMux I__2917 (
            .O(N__11765),
            .I(N__11762));
    LocalMux I__2916 (
            .O(N__11762),
            .I(N__11759));
    Span4Mux_s3_h I__2915 (
            .O(N__11759),
            .I(N__11756));
    Span4Mux_v I__2914 (
            .O(N__11756),
            .I(N__11753));
    Odrv4 I__2913 (
            .O(N__11753),
            .I(N_221_i));
    InMux I__2912 (
            .O(N__11750),
            .I(N__11747));
    LocalMux I__2911 (
            .O(N__11747),
            .I(N__11744));
    Span12Mux_h I__2910 (
            .O(N__11744),
            .I(N__11741));
    Odrv12 I__2909 (
            .O(N__11741),
            .I(READ_CYCLE_ACTIVE_rep21_i_ess));
    IoInMux I__2908 (
            .O(N__11738),
            .I(N__11735));
    LocalMux I__2907 (
            .O(N__11735),
            .I(N__11732));
    Span12Mux_s8_h I__2906 (
            .O(N__11732),
            .I(N__11729));
    Odrv12 I__2905 (
            .O(N__11729),
            .I(N_226_i));
    InMux I__2904 (
            .O(N__11726),
            .I(N__11723));
    LocalMux I__2903 (
            .O(N__11723),
            .I(N__11720));
    Span12Mux_s10_h I__2902 (
            .O(N__11720),
            .I(N__11717));
    Odrv12 I__2901 (
            .O(N__11717),
            .I(READ_CYCLE_ACTIVE_rep24_i_ess));
    IoInMux I__2900 (
            .O(N__11714),
            .I(N__11711));
    LocalMux I__2899 (
            .O(N__11711),
            .I(N__11708));
    Span4Mux_s3_h I__2898 (
            .O(N__11708),
            .I(N__11705));
    Span4Mux_v I__2897 (
            .O(N__11705),
            .I(N__11702));
    Sp12to4 I__2896 (
            .O(N__11702),
            .I(N__11699));
    Span12Mux_s9_h I__2895 (
            .O(N__11699),
            .I(N__11696));
    Span12Mux_v I__2894 (
            .O(N__11696),
            .I(N__11693));
    Odrv12 I__2893 (
            .O(N__11693),
            .I(N_229_i));
    InMux I__2892 (
            .O(N__11690),
            .I(N__11687));
    LocalMux I__2891 (
            .O(N__11687),
            .I(N__11684));
    Span12Mux_s10_h I__2890 (
            .O(N__11684),
            .I(N__11681));
    Odrv12 I__2889 (
            .O(N__11681),
            .I(READ_CYCLE_ACTIVE_rep9_i_ess));
    IoInMux I__2888 (
            .O(N__11678),
            .I(N__11675));
    LocalMux I__2887 (
            .O(N__11675),
            .I(N__11672));
    Span4Mux_s1_h I__2886 (
            .O(N__11672),
            .I(N__11669));
    Span4Mux_h I__2885 (
            .O(N__11669),
            .I(N__11666));
    Span4Mux_v I__2884 (
            .O(N__11666),
            .I(N__11663));
    Span4Mux_v I__2883 (
            .O(N__11663),
            .I(N__11660));
    Odrv4 I__2882 (
            .O(N__11660),
            .I(N_214_i));
    InMux I__2881 (
            .O(N__11657),
            .I(N__11654));
    LocalMux I__2880 (
            .O(N__11654),
            .I(N__11651));
    Span4Mux_v I__2879 (
            .O(N__11651),
            .I(N__11648));
    Sp12to4 I__2878 (
            .O(N__11648),
            .I(N__11645));
    Odrv12 I__2877 (
            .O(N__11645),
            .I(READ_CYCLE_ACTIVE_rep12_i_ess));
    IoInMux I__2876 (
            .O(N__11642),
            .I(N__11639));
    LocalMux I__2875 (
            .O(N__11639),
            .I(N__11636));
    Span4Mux_s0_v I__2874 (
            .O(N__11636),
            .I(N__11633));
    Span4Mux_h I__2873 (
            .O(N__11633),
            .I(N__11630));
    Span4Mux_v I__2872 (
            .O(N__11630),
            .I(N__11627));
    Span4Mux_v I__2871 (
            .O(N__11627),
            .I(N__11624));
    Odrv4 I__2870 (
            .O(N__11624),
            .I(N_217_i));
    InMux I__2869 (
            .O(N__11621),
            .I(N__11618));
    LocalMux I__2868 (
            .O(N__11618),
            .I(N__11615));
    Span4Mux_v I__2867 (
            .O(N__11615),
            .I(N__11612));
    Sp12to4 I__2866 (
            .O(N__11612),
            .I(N__11609));
    Odrv12 I__2865 (
            .O(N__11609),
            .I(READ_CYCLE_ACTIVE_rep8_i_ess));
    IoInMux I__2864 (
            .O(N__11606),
            .I(N__11603));
    LocalMux I__2863 (
            .O(N__11603),
            .I(N__11600));
    Span4Mux_s2_h I__2862 (
            .O(N__11600),
            .I(N__11597));
    Span4Mux_h I__2861 (
            .O(N__11597),
            .I(N__11594));
    Odrv4 I__2860 (
            .O(N__11594),
            .I(N_213_i));
    InMux I__2859 (
            .O(N__11591),
            .I(N__11588));
    LocalMux I__2858 (
            .O(N__11588),
            .I(N__11585));
    Span12Mux_v I__2857 (
            .O(N__11585),
            .I(N__11582));
    Span12Mux_h I__2856 (
            .O(N__11582),
            .I(N__11579));
    Odrv12 I__2855 (
            .O(N__11579),
            .I(READ_CYCLE_ACTIVE_rep23_i_ess));
    IoInMux I__2854 (
            .O(N__11576),
            .I(N__11573));
    LocalMux I__2853 (
            .O(N__11573),
            .I(N__11570));
    Span4Mux_s2_h I__2852 (
            .O(N__11570),
            .I(N__11567));
    Span4Mux_h I__2851 (
            .O(N__11567),
            .I(N__11564));
    Odrv4 I__2850 (
            .O(N__11564),
            .I(N_228_i));
    InMux I__2849 (
            .O(N__11561),
            .I(N__11558));
    LocalMux I__2848 (
            .O(N__11558),
            .I(N__11555));
    Span4Mux_h I__2847 (
            .O(N__11555),
            .I(N__11552));
    Odrv4 I__2846 (
            .O(N__11552),
            .I(READ_CYCLE_ACTIVE_rep20_i_ess));
    IoInMux I__2845 (
            .O(N__11549),
            .I(N__11546));
    LocalMux I__2844 (
            .O(N__11546),
            .I(N__11543));
    IoSpan4Mux I__2843 (
            .O(N__11543),
            .I(N__11540));
    IoSpan4Mux I__2842 (
            .O(N__11540),
            .I(N__11537));
    Span4Mux_s1_h I__2841 (
            .O(N__11537),
            .I(N__11534));
    Odrv4 I__2840 (
            .O(N__11534),
            .I(N_225_i));
    InMux I__2839 (
            .O(N__11531),
            .I(N__11528));
    LocalMux I__2838 (
            .O(N__11528),
            .I(N__11525));
    Span4Mux_v I__2837 (
            .O(N__11525),
            .I(N__11522));
    Sp12to4 I__2836 (
            .O(N__11522),
            .I(N__11519));
    Odrv12 I__2835 (
            .O(N__11519),
            .I(READ_CYCLE_ACTIVE_rep3_i_ess));
    IoInMux I__2834 (
            .O(N__11516),
            .I(N__11513));
    LocalMux I__2833 (
            .O(N__11513),
            .I(N__11510));
    Span12Mux_s7_v I__2832 (
            .O(N__11510),
            .I(N__11507));
    Odrv12 I__2831 (
            .O(N__11507),
            .I(N_208_i));
    InMux I__2830 (
            .O(N__11504),
            .I(N__11501));
    LocalMux I__2829 (
            .O(N__11501),
            .I(N__11498));
    Span4Mux_v I__2828 (
            .O(N__11498),
            .I(N__11495));
    Span4Mux_v I__2827 (
            .O(N__11495),
            .I(N__11492));
    Sp12to4 I__2826 (
            .O(N__11492),
            .I(N__11489));
    Odrv12 I__2825 (
            .O(N__11489),
            .I(D_UM_040_in_7));
    IoInMux I__2824 (
            .O(N__11486),
            .I(N__11483));
    LocalMux I__2823 (
            .O(N__11483),
            .I(N__11479));
    InMux I__2822 (
            .O(N__11482),
            .I(N__11476));
    IoSpan4Mux I__2821 (
            .O(N__11479),
            .I(N__11473));
    LocalMux I__2820 (
            .O(N__11476),
            .I(N__11470));
    Span4Mux_s3_h I__2819 (
            .O(N__11473),
            .I(N__11467));
    Span4Mux_h I__2818 (
            .O(N__11470),
            .I(N__11464));
    Sp12to4 I__2817 (
            .O(N__11467),
            .I(N__11461));
    Sp12to4 I__2816 (
            .O(N__11464),
            .I(N__11458));
    Span12Mux_v I__2815 (
            .O(N__11461),
            .I(N__11455));
    Span12Mux_v I__2814 (
            .O(N__11458),
            .I(N__11452));
    Span12Mux_h I__2813 (
            .O(N__11455),
            .I(N__11449));
    Span12Mux_v I__2812 (
            .O(N__11452),
            .I(N__11446));
    Span12Mux_h I__2811 (
            .O(N__11449),
            .I(N__11443));
    Span12Mux_h I__2810 (
            .O(N__11446),
            .I(N__11440));
    Odrv12 I__2809 (
            .O(N__11443),
            .I(D_LL_040_in_7));
    Odrv12 I__2808 (
            .O(N__11440),
            .I(D_LL_040_in_7));
    IoInMux I__2807 (
            .O(N__11435),
            .I(N__11432));
    LocalMux I__2806 (
            .O(N__11432),
            .I(N__11429));
    IoSpan4Mux I__2805 (
            .O(N__11429),
            .I(N__11426));
    Span4Mux_s2_h I__2804 (
            .O(N__11426),
            .I(N__11423));
    Span4Mux_h I__2803 (
            .O(N__11423),
            .I(N__11420));
    Sp12to4 I__2802 (
            .O(N__11420),
            .I(N__11417));
    Span12Mux_h I__2801 (
            .O(N__11417),
            .I(N__11414));
    Odrv12 I__2800 (
            .O(N__11414),
            .I(un1_D_UM_040_7));
    InMux I__2799 (
            .O(N__11411),
            .I(N__11408));
    LocalMux I__2798 (
            .O(N__11408),
            .I(N__11405));
    Odrv12 I__2797 (
            .O(N__11405),
            .I(READ_CYCLE_ACTIVE_rep28_i_ess));
    IoInMux I__2796 (
            .O(N__11402),
            .I(N__11399));
    LocalMux I__2795 (
            .O(N__11399),
            .I(N__11396));
    Span4Mux_s1_h I__2794 (
            .O(N__11396),
            .I(N__11393));
    Sp12to4 I__2793 (
            .O(N__11393),
            .I(N__11390));
    Span12Mux_s11_v I__2792 (
            .O(N__11390),
            .I(N__11387));
    Odrv12 I__2791 (
            .O(N__11387),
            .I(N_233_i));
    InMux I__2790 (
            .O(N__11384),
            .I(N__11381));
    LocalMux I__2789 (
            .O(N__11381),
            .I(N__11378));
    Span4Mux_v I__2788 (
            .O(N__11378),
            .I(N__11375));
    Sp12to4 I__2787 (
            .O(N__11375),
            .I(N__11372));
    Odrv12 I__2786 (
            .O(N__11372),
            .I(READ_CYCLE_ACTIVE_rep30_i_ess));
    IoInMux I__2785 (
            .O(N__11369),
            .I(N__11366));
    LocalMux I__2784 (
            .O(N__11366),
            .I(N__11363));
    Span4Mux_s3_h I__2783 (
            .O(N__11363),
            .I(N__11360));
    Sp12to4 I__2782 (
            .O(N__11360),
            .I(N__11357));
    Span12Mux_s11_v I__2781 (
            .O(N__11357),
            .I(N__11354));
    Odrv12 I__2780 (
            .O(N__11354),
            .I(N_235_i));
    InMux I__2779 (
            .O(N__11351),
            .I(N__11348));
    LocalMux I__2778 (
            .O(N__11348),
            .I(N__11345));
    Span4Mux_v I__2777 (
            .O(N__11345),
            .I(N__11342));
    Sp12to4 I__2776 (
            .O(N__11342),
            .I(N__11339));
    Span12Mux_h I__2775 (
            .O(N__11339),
            .I(N__11336));
    Odrv12 I__2774 (
            .O(N__11336),
            .I(READ_CYCLE_ACTIVE_rep17_i_ess));
    IoInMux I__2773 (
            .O(N__11333),
            .I(N__11330));
    LocalMux I__2772 (
            .O(N__11330),
            .I(N__11327));
    Span12Mux_s9_h I__2771 (
            .O(N__11327),
            .I(N__11324));
    Odrv12 I__2770 (
            .O(N__11324),
            .I(N_222_i));
    InMux I__2769 (
            .O(N__11321),
            .I(N__11318));
    LocalMux I__2768 (
            .O(N__11318),
            .I(N__11315));
    Span4Mux_h I__2767 (
            .O(N__11315),
            .I(N__11312));
    Span4Mux_v I__2766 (
            .O(N__11312),
            .I(N__11309));
    Span4Mux_h I__2765 (
            .O(N__11309),
            .I(N__11306));
    Odrv4 I__2764 (
            .O(N__11306),
            .I(D_UM_040_in_4));
    IoInMux I__2763 (
            .O(N__11303),
            .I(N__11299));
    InMux I__2762 (
            .O(N__11302),
            .I(N__11296));
    LocalMux I__2761 (
            .O(N__11299),
            .I(N__11293));
    LocalMux I__2760 (
            .O(N__11296),
            .I(N__11290));
    Span4Mux_s2_h I__2759 (
            .O(N__11293),
            .I(N__11287));
    Span4Mux_v I__2758 (
            .O(N__11290),
            .I(N__11284));
    Span4Mux_v I__2757 (
            .O(N__11287),
            .I(N__11281));
    Sp12to4 I__2756 (
            .O(N__11284),
            .I(N__11278));
    Sp12to4 I__2755 (
            .O(N__11281),
            .I(N__11275));
    Span12Mux_h I__2754 (
            .O(N__11278),
            .I(N__11272));
    Span12Mux_h I__2753 (
            .O(N__11275),
            .I(N__11269));
    Span12Mux_v I__2752 (
            .O(N__11272),
            .I(N__11266));
    Span12Mux_h I__2751 (
            .O(N__11269),
            .I(N__11263));
    Span12Mux_v I__2750 (
            .O(N__11266),
            .I(N__11260));
    Odrv12 I__2749 (
            .O(N__11263),
            .I(D_LL_040_in_4));
    Odrv12 I__2748 (
            .O(N__11260),
            .I(D_LL_040_in_4));
    IoInMux I__2747 (
            .O(N__11255),
            .I(N__11252));
    LocalMux I__2746 (
            .O(N__11252),
            .I(N__11249));
    Span4Mux_s1_h I__2745 (
            .O(N__11249),
            .I(N__11246));
    Sp12to4 I__2744 (
            .O(N__11246),
            .I(N__11243));
    Span12Mux_s7_v I__2743 (
            .O(N__11243),
            .I(N__11240));
    Span12Mux_h I__2742 (
            .O(N__11240),
            .I(N__11237));
    Odrv12 I__2741 (
            .O(N__11237),
            .I(un1_D_UM_040_4));
    IoInMux I__2740 (
            .O(N__11234),
            .I(N__11231));
    LocalMux I__2739 (
            .O(N__11231),
            .I(N__11228));
    IoSpan4Mux I__2738 (
            .O(N__11228),
            .I(N__11225));
    Span4Mux_s3_h I__2737 (
            .O(N__11225),
            .I(N__11221));
    InMux I__2736 (
            .O(N__11224),
            .I(N__11218));
    Sp12to4 I__2735 (
            .O(N__11221),
            .I(N__11215));
    LocalMux I__2734 (
            .O(N__11218),
            .I(N__11212));
    Span12Mux_v I__2733 (
            .O(N__11215),
            .I(N__11209));
    Sp12to4 I__2732 (
            .O(N__11212),
            .I(N__11206));
    Span12Mux_h I__2731 (
            .O(N__11209),
            .I(N__11203));
    Span12Mux_v I__2730 (
            .O(N__11206),
            .I(N__11200));
    Span12Mux_h I__2729 (
            .O(N__11203),
            .I(N__11197));
    Span12Mux_v I__2728 (
            .O(N__11200),
            .I(N__11194));
    Odrv12 I__2727 (
            .O(N__11197),
            .I(D_LL_040_in_5));
    Odrv12 I__2726 (
            .O(N__11194),
            .I(D_LL_040_in_5));
    InMux I__2725 (
            .O(N__11189),
            .I(N__11186));
    LocalMux I__2724 (
            .O(N__11186),
            .I(N__11183));
    Span4Mux_v I__2723 (
            .O(N__11183),
            .I(N__11180));
    Span4Mux_h I__2722 (
            .O(N__11180),
            .I(N__11177));
    IoSpan4Mux I__2721 (
            .O(N__11177),
            .I(N__11174));
    Odrv4 I__2720 (
            .O(N__11174),
            .I(D_UM_040_in_5));
    InMux I__2719 (
            .O(N__11171),
            .I(N__11158));
    InMux I__2718 (
            .O(N__11170),
            .I(N__11155));
    InMux I__2717 (
            .O(N__11169),
            .I(N__11152));
    InMux I__2716 (
            .O(N__11168),
            .I(N__11148));
    InMux I__2715 (
            .O(N__11167),
            .I(N__11145));
    InMux I__2714 (
            .O(N__11166),
            .I(N__11140));
    InMux I__2713 (
            .O(N__11165),
            .I(N__11134));
    InMux I__2712 (
            .O(N__11164),
            .I(N__11134));
    InMux I__2711 (
            .O(N__11163),
            .I(N__11131));
    InMux I__2710 (
            .O(N__11162),
            .I(N__11126));
    InMux I__2709 (
            .O(N__11161),
            .I(N__11123));
    LocalMux I__2708 (
            .O(N__11158),
            .I(N__11112));
    LocalMux I__2707 (
            .O(N__11155),
            .I(N__11112));
    LocalMux I__2706 (
            .O(N__11152),
            .I(N__11108));
    InMux I__2705 (
            .O(N__11151),
            .I(N__11105));
    LocalMux I__2704 (
            .O(N__11148),
            .I(N__11102));
    LocalMux I__2703 (
            .O(N__11145),
            .I(N__11099));
    InMux I__2702 (
            .O(N__11144),
            .I(N__11094));
    InMux I__2701 (
            .O(N__11143),
            .I(N__11094));
    LocalMux I__2700 (
            .O(N__11140),
            .I(N__11090));
    InMux I__2699 (
            .O(N__11139),
            .I(N__11087));
    LocalMux I__2698 (
            .O(N__11134),
            .I(N__11083));
    LocalMux I__2697 (
            .O(N__11131),
            .I(N__11080));
    InMux I__2696 (
            .O(N__11130),
            .I(N__11077));
    InMux I__2695 (
            .O(N__11129),
            .I(N__11073));
    LocalMux I__2694 (
            .O(N__11126),
            .I(N__11068));
    LocalMux I__2693 (
            .O(N__11123),
            .I(N__11068));
    InMux I__2692 (
            .O(N__11122),
            .I(N__11065));
    InMux I__2691 (
            .O(N__11121),
            .I(N__11062));
    InMux I__2690 (
            .O(N__11120),
            .I(N__11058));
    InMux I__2689 (
            .O(N__11119),
            .I(N__11055));
    InMux I__2688 (
            .O(N__11118),
            .I(N__11052));
    InMux I__2687 (
            .O(N__11117),
            .I(N__11049));
    Span4Mux_v I__2686 (
            .O(N__11112),
            .I(N__11043));
    InMux I__2685 (
            .O(N__11111),
            .I(N__11040));
    Span4Mux_v I__2684 (
            .O(N__11108),
            .I(N__11037));
    LocalMux I__2683 (
            .O(N__11105),
            .I(N__11034));
    Span4Mux_v I__2682 (
            .O(N__11102),
            .I(N__11031));
    Span4Mux_h I__2681 (
            .O(N__11099),
            .I(N__11026));
    LocalMux I__2680 (
            .O(N__11094),
            .I(N__11026));
    InMux I__2679 (
            .O(N__11093),
            .I(N__11023));
    Span4Mux_v I__2678 (
            .O(N__11090),
            .I(N__11018));
    LocalMux I__2677 (
            .O(N__11087),
            .I(N__11018));
    InMux I__2676 (
            .O(N__11086),
            .I(N__11015));
    Span4Mux_v I__2675 (
            .O(N__11083),
            .I(N__11012));
    Span4Mux_h I__2674 (
            .O(N__11080),
            .I(N__11007));
    LocalMux I__2673 (
            .O(N__11077),
            .I(N__11007));
    InMux I__2672 (
            .O(N__11076),
            .I(N__11004));
    LocalMux I__2671 (
            .O(N__11073),
            .I(N__11001));
    Span4Mux_v I__2670 (
            .O(N__11068),
            .I(N__10996));
    LocalMux I__2669 (
            .O(N__11065),
            .I(N__10996));
    LocalMux I__2668 (
            .O(N__11062),
            .I(N__10993));
    InMux I__2667 (
            .O(N__11061),
            .I(N__10990));
    LocalMux I__2666 (
            .O(N__11058),
            .I(N__10985));
    LocalMux I__2665 (
            .O(N__11055),
            .I(N__10985));
    LocalMux I__2664 (
            .O(N__11052),
            .I(N__10980));
    LocalMux I__2663 (
            .O(N__11049),
            .I(N__10980));
    InMux I__2662 (
            .O(N__11048),
            .I(N__10977));
    InMux I__2661 (
            .O(N__11047),
            .I(N__10972));
    InMux I__2660 (
            .O(N__11046),
            .I(N__10972));
    Span4Mux_v I__2659 (
            .O(N__11043),
            .I(N__10967));
    LocalMux I__2658 (
            .O(N__11040),
            .I(N__10964));
    Span4Mux_v I__2657 (
            .O(N__11037),
            .I(N__10959));
    Span4Mux_v I__2656 (
            .O(N__11034),
            .I(N__10959));
    Span4Mux_h I__2655 (
            .O(N__11031),
            .I(N__10954));
    Span4Mux_v I__2654 (
            .O(N__11026),
            .I(N__10954));
    LocalMux I__2653 (
            .O(N__11023),
            .I(N__10951));
    Span4Mux_v I__2652 (
            .O(N__11018),
            .I(N__10946));
    LocalMux I__2651 (
            .O(N__11015),
            .I(N__10946));
    Span4Mux_h I__2650 (
            .O(N__11012),
            .I(N__10939));
    Span4Mux_h I__2649 (
            .O(N__11007),
            .I(N__10939));
    LocalMux I__2648 (
            .O(N__11004),
            .I(N__10939));
    Span4Mux_v I__2647 (
            .O(N__11001),
            .I(N__10936));
    Span4Mux_v I__2646 (
            .O(N__10996),
            .I(N__10933));
    Span4Mux_v I__2645 (
            .O(N__10993),
            .I(N__10928));
    LocalMux I__2644 (
            .O(N__10990),
            .I(N__10928));
    Span4Mux_v I__2643 (
            .O(N__10985),
            .I(N__10921));
    Span4Mux_h I__2642 (
            .O(N__10980),
            .I(N__10921));
    LocalMux I__2641 (
            .O(N__10977),
            .I(N__10921));
    LocalMux I__2640 (
            .O(N__10972),
            .I(N__10918));
    InMux I__2639 (
            .O(N__10971),
            .I(N__10915));
    CascadeMux I__2638 (
            .O(N__10970),
            .I(N__10912));
    Sp12to4 I__2637 (
            .O(N__10967),
            .I(N__10907));
    Span12Mux_v I__2636 (
            .O(N__10964),
            .I(N__10907));
    Span4Mux_h I__2635 (
            .O(N__10959),
            .I(N__10900));
    Span4Mux_v I__2634 (
            .O(N__10954),
            .I(N__10900));
    Span4Mux_v I__2633 (
            .O(N__10951),
            .I(N__10900));
    Span4Mux_h I__2632 (
            .O(N__10946),
            .I(N__10895));
    Span4Mux_v I__2631 (
            .O(N__10939),
            .I(N__10895));
    Span4Mux_h I__2630 (
            .O(N__10936),
            .I(N__10884));
    Span4Mux_v I__2629 (
            .O(N__10933),
            .I(N__10884));
    Span4Mux_v I__2628 (
            .O(N__10928),
            .I(N__10884));
    Span4Mux_v I__2627 (
            .O(N__10921),
            .I(N__10884));
    Span4Mux_v I__2626 (
            .O(N__10918),
            .I(N__10884));
    LocalMux I__2625 (
            .O(N__10915),
            .I(N__10881));
    InMux I__2624 (
            .O(N__10912),
            .I(N__10878));
    Odrv12 I__2623 (
            .O(N__10907),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv4 I__2622 (
            .O(N__10900),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv4 I__2621 (
            .O(N__10895),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv4 I__2620 (
            .O(N__10884),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv4 I__2619 (
            .O(N__10881),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    LocalMux I__2618 (
            .O(N__10878),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    IoInMux I__2617 (
            .O(N__10865),
            .I(N__10862));
    LocalMux I__2616 (
            .O(N__10862),
            .I(N__10859));
    Span12Mux_s6_v I__2615 (
            .O(N__10859),
            .I(N__10856));
    Span12Mux_h I__2614 (
            .O(N__10856),
            .I(N__10853));
    Odrv12 I__2613 (
            .O(N__10853),
            .I(un1_D_UM_040_5));
    InMux I__2612 (
            .O(N__10850),
            .I(N__10847));
    LocalMux I__2611 (
            .O(N__10847),
            .I(N__10844));
    Span4Mux_v I__2610 (
            .O(N__10844),
            .I(N__10841));
    Sp12to4 I__2609 (
            .O(N__10841),
            .I(N__10838));
    Odrv12 I__2608 (
            .O(N__10838),
            .I(READ_CYCLE_ACTIVE_rep25_i_ess));
    IoInMux I__2607 (
            .O(N__10835),
            .I(N__10832));
    LocalMux I__2606 (
            .O(N__10832),
            .I(N__10829));
    IoSpan4Mux I__2605 (
            .O(N__10829),
            .I(N__10826));
    Span4Mux_s2_h I__2604 (
            .O(N__10826),
            .I(N__10823));
    Sp12to4 I__2603 (
            .O(N__10823),
            .I(N__10820));
    Span12Mux_v I__2602 (
            .O(N__10820),
            .I(N__10817));
    Odrv12 I__2601 (
            .O(N__10817),
            .I(N_230_i));
    InMux I__2600 (
            .O(N__10814),
            .I(N__10811));
    LocalMux I__2599 (
            .O(N__10811),
            .I(N__10808));
    Span4Mux_h I__2598 (
            .O(N__10808),
            .I(N__10805));
    Odrv4 I__2597 (
            .O(N__10805),
            .I(READ_CYCLE_ACTIVE_rep10_i_ess));
    IoInMux I__2596 (
            .O(N__10802),
            .I(N__10799));
    LocalMux I__2595 (
            .O(N__10799),
            .I(N__10796));
    Odrv12 I__2594 (
            .O(N__10796),
            .I(N_215_i));
    InMux I__2593 (
            .O(N__10793),
            .I(N__10790));
    LocalMux I__2592 (
            .O(N__10790),
            .I(N__10787));
    Span12Mux_h I__2591 (
            .O(N__10787),
            .I(N__10784));
    Odrv12 I__2590 (
            .O(N__10784),
            .I(READ_CYCLE_ACTIVE_rep27_i_ess));
    IoInMux I__2589 (
            .O(N__10781),
            .I(N__10778));
    LocalMux I__2588 (
            .O(N__10778),
            .I(N__10775));
    IoSpan4Mux I__2587 (
            .O(N__10775),
            .I(N__10772));
    Span4Mux_s2_v I__2586 (
            .O(N__10772),
            .I(N__10769));
    Span4Mux_v I__2585 (
            .O(N__10769),
            .I(N__10766));
    Span4Mux_h I__2584 (
            .O(N__10766),
            .I(N__10763));
    Odrv4 I__2583 (
            .O(N__10763),
            .I(N_232_i));
    InMux I__2582 (
            .O(N__10760),
            .I(N__10757));
    LocalMux I__2581 (
            .O(N__10757),
            .I(N__10754));
    Odrv12 I__2580 (
            .O(N__10754),
            .I(READ_CYCLE_ACTIVE_rep18_i_ess));
    IoInMux I__2579 (
            .O(N__10751),
            .I(N__10748));
    LocalMux I__2578 (
            .O(N__10748),
            .I(N__10745));
    IoSpan4Mux I__2577 (
            .O(N__10745),
            .I(N__10742));
    Span4Mux_s3_h I__2576 (
            .O(N__10742),
            .I(N__10739));
    Span4Mux_v I__2575 (
            .O(N__10739),
            .I(N__10736));
    Span4Mux_h I__2574 (
            .O(N__10736),
            .I(N__10733));
    Odrv4 I__2573 (
            .O(N__10733),
            .I(N_223_i));
    InMux I__2572 (
            .O(N__10730),
            .I(N__10727));
    LocalMux I__2571 (
            .O(N__10727),
            .I(N__10724));
    Span4Mux_v I__2570 (
            .O(N__10724),
            .I(N__10721));
    Span4Mux_h I__2569 (
            .O(N__10721),
            .I(N__10718));
    Odrv4 I__2568 (
            .O(N__10718),
            .I(READ_CYCLE_ACTIVE_rep0_i_ess));
    IoInMux I__2567 (
            .O(N__10715),
            .I(N__10712));
    LocalMux I__2566 (
            .O(N__10712),
            .I(N__10709));
    Span4Mux_s1_v I__2565 (
            .O(N__10709),
            .I(N__10706));
    Span4Mux_h I__2564 (
            .O(N__10706),
            .I(N__10703));
    Span4Mux_v I__2563 (
            .O(N__10703),
            .I(N__10700));
    Span4Mux_v I__2562 (
            .O(N__10700),
            .I(N__10697));
    Odrv4 I__2561 (
            .O(N__10697),
            .I(N_205_i));
    InMux I__2560 (
            .O(N__10694),
            .I(N__10691));
    LocalMux I__2559 (
            .O(N__10691),
            .I(N__10688));
    Span4Mux_v I__2558 (
            .O(N__10688),
            .I(N__10685));
    Span4Mux_h I__2557 (
            .O(N__10685),
            .I(N__10682));
    Odrv4 I__2556 (
            .O(N__10682),
            .I(READ_CYCLE_ACTIVE_rep7_i_ess));
    IoInMux I__2555 (
            .O(N__10679),
            .I(N__10676));
    LocalMux I__2554 (
            .O(N__10676),
            .I(N__10673));
    Span4Mux_s3_v I__2553 (
            .O(N__10673),
            .I(N__10670));
    Sp12to4 I__2552 (
            .O(N__10670),
            .I(N__10667));
    Span12Mux_s11_h I__2551 (
            .O(N__10667),
            .I(N__10664));
    Odrv12 I__2550 (
            .O(N__10664),
            .I(N_212_i));
    InMux I__2549 (
            .O(N__10661),
            .I(N__10658));
    LocalMux I__2548 (
            .O(N__10658),
            .I(N__10655));
    Span12Mux_h I__2547 (
            .O(N__10655),
            .I(N__10652));
    Odrv12 I__2546 (
            .O(N__10652),
            .I(D_UM_040_in_2));
    IoInMux I__2545 (
            .O(N__10649),
            .I(N__10646));
    LocalMux I__2544 (
            .O(N__10646),
            .I(N__10643));
    IoSpan4Mux I__2543 (
            .O(N__10643),
            .I(N__10640));
    Span4Mux_s2_h I__2542 (
            .O(N__10640),
            .I(N__10636));
    InMux I__2541 (
            .O(N__10639),
            .I(N__10633));
    Sp12to4 I__2540 (
            .O(N__10636),
            .I(N__10630));
    LocalMux I__2539 (
            .O(N__10633),
            .I(N__10627));
    Span12Mux_h I__2538 (
            .O(N__10630),
            .I(N__10624));
    Span12Mux_v I__2537 (
            .O(N__10627),
            .I(N__10621));
    Span12Mux_h I__2536 (
            .O(N__10624),
            .I(N__10618));
    Span12Mux_v I__2535 (
            .O(N__10621),
            .I(N__10615));
    Odrv12 I__2534 (
            .O(N__10618),
            .I(D_LL_040_in_2));
    Odrv12 I__2533 (
            .O(N__10615),
            .I(D_LL_040_in_2));
    IoInMux I__2532 (
            .O(N__10610),
            .I(N__10607));
    LocalMux I__2531 (
            .O(N__10607),
            .I(N__10604));
    Span4Mux_s2_h I__2530 (
            .O(N__10604),
            .I(N__10601));
    Span4Mux_v I__2529 (
            .O(N__10601),
            .I(N__10598));
    Sp12to4 I__2528 (
            .O(N__10598),
            .I(N__10595));
    Span12Mux_h I__2527 (
            .O(N__10595),
            .I(N__10592));
    Odrv12 I__2526 (
            .O(N__10592),
            .I(un1_D_UM_040_2));
    InMux I__2525 (
            .O(N__10589),
            .I(N__10586));
    LocalMux I__2524 (
            .O(N__10586),
            .I(N__10583));
    Odrv12 I__2523 (
            .O(N__10583),
            .I(READ_CYCLE_ACTIVE_rep31_i_ess));
    IoInMux I__2522 (
            .O(N__10580),
            .I(N__10577));
    LocalMux I__2521 (
            .O(N__10577),
            .I(N__10574));
    Span12Mux_s10_h I__2520 (
            .O(N__10574),
            .I(N__10571));
    Span12Mux_v I__2519 (
            .O(N__10571),
            .I(N__10568));
    Odrv12 I__2518 (
            .O(N__10568),
            .I(N_236_i));
    InMux I__2517 (
            .O(N__10565),
            .I(N__10562));
    LocalMux I__2516 (
            .O(N__10562),
            .I(N__10559));
    Odrv12 I__2515 (
            .O(N__10559),
            .I(READ_CYCLE_ACTIVE_rep22_i_ess));
    IoInMux I__2514 (
            .O(N__10556),
            .I(N__10553));
    LocalMux I__2513 (
            .O(N__10553),
            .I(N__10550));
    IoSpan4Mux I__2512 (
            .O(N__10550),
            .I(N__10547));
    Span4Mux_s2_h I__2511 (
            .O(N__10547),
            .I(N__10544));
    Span4Mux_h I__2510 (
            .O(N__10544),
            .I(N__10541));
    Odrv4 I__2509 (
            .O(N__10541),
            .I(N_227_i));
    InMux I__2508 (
            .O(N__10538),
            .I(N__10535));
    LocalMux I__2507 (
            .O(N__10535),
            .I(N__10532));
    Span4Mux_v I__2506 (
            .O(N__10532),
            .I(N__10529));
    Span4Mux_h I__2505 (
            .O(N__10529),
            .I(N__10526));
    Odrv4 I__2504 (
            .O(N__10526),
            .I(READ_CYCLE_ACTIVE_rep13_i_ess));
    IoInMux I__2503 (
            .O(N__10523),
            .I(N__10520));
    LocalMux I__2502 (
            .O(N__10520),
            .I(N__10517));
    Span4Mux_s0_v I__2501 (
            .O(N__10517),
            .I(N__10514));
    Sp12to4 I__2500 (
            .O(N__10514),
            .I(N__10511));
    Span12Mux_s10_h I__2499 (
            .O(N__10511),
            .I(N__10508));
    Odrv12 I__2498 (
            .O(N__10508),
            .I(N_218_i));
    InMux I__2497 (
            .O(N__10505),
            .I(N__10502));
    LocalMux I__2496 (
            .O(N__10502),
            .I(N__10499));
    Span4Mux_v I__2495 (
            .O(N__10499),
            .I(N__10496));
    Sp12to4 I__2494 (
            .O(N__10496),
            .I(N__10493));
    Odrv12 I__2493 (
            .O(N__10493),
            .I(READ_CYCLE_ACTIVE_rep4_i_ess));
    IoInMux I__2492 (
            .O(N__10490),
            .I(N__10487));
    LocalMux I__2491 (
            .O(N__10487),
            .I(N__10484));
    Span4Mux_s2_v I__2490 (
            .O(N__10484),
            .I(N__10481));
    Span4Mux_h I__2489 (
            .O(N__10481),
            .I(N__10478));
    Span4Mux_v I__2488 (
            .O(N__10478),
            .I(N__10475));
    Odrv4 I__2487 (
            .O(N__10475),
            .I(N_209_i));
    InMux I__2486 (
            .O(N__10472),
            .I(N__10468));
    InMux I__2485 (
            .O(N__10471),
            .I(N__10465));
    LocalMux I__2484 (
            .O(N__10468),
            .I(N__10462));
    LocalMux I__2483 (
            .O(N__10465),
            .I(N__10458));
    Span4Mux_v I__2482 (
            .O(N__10462),
            .I(N__10455));
    InMux I__2481 (
            .O(N__10461),
            .I(N__10452));
    Span4Mux_v I__2480 (
            .O(N__10458),
            .I(N__10449));
    Span4Mux_v I__2479 (
            .O(N__10455),
            .I(N__10446));
    LocalMux I__2478 (
            .O(N__10452),
            .I(N__10443));
    Span4Mux_v I__2477 (
            .O(N__10449),
            .I(N__10440));
    Sp12to4 I__2476 (
            .O(N__10446),
            .I(N__10435));
    Span12Mux_h I__2475 (
            .O(N__10443),
            .I(N__10435));
    Span4Mux_h I__2474 (
            .O(N__10440),
            .I(N__10432));
    Span12Mux_h I__2473 (
            .O(N__10435),
            .I(N__10429));
    IoSpan4Mux I__2472 (
            .O(N__10432),
            .I(N__10426));
    Odrv12 I__2471 (
            .O(N__10429),
            .I(D_UU_AMIGA_in_7));
    Odrv4 I__2470 (
            .O(N__10426),
            .I(D_UU_AMIGA_in_7));
    InMux I__2469 (
            .O(N__10421),
            .I(N__10418));
    LocalMux I__2468 (
            .O(N__10418),
            .I(N__10415));
    Span4Mux_v I__2467 (
            .O(N__10415),
            .I(N__10412));
    Odrv4 I__2466 (
            .O(N__10412),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ));
    InMux I__2465 (
            .O(N__10409),
            .I(N__10396));
    InMux I__2464 (
            .O(N__10408),
            .I(N__10396));
    InMux I__2463 (
            .O(N__10407),
            .I(N__10396));
    InMux I__2462 (
            .O(N__10406),
            .I(N__10390));
    InMux I__2461 (
            .O(N__10405),
            .I(N__10385));
    InMux I__2460 (
            .O(N__10404),
            .I(N__10385));
    InMux I__2459 (
            .O(N__10403),
            .I(N__10382));
    LocalMux I__2458 (
            .O(N__10396),
            .I(N__10376));
    InMux I__2457 (
            .O(N__10395),
            .I(N__10371));
    InMux I__2456 (
            .O(N__10394),
            .I(N__10371));
    InMux I__2455 (
            .O(N__10393),
            .I(N__10368));
    LocalMux I__2454 (
            .O(N__10390),
            .I(N__10360));
    LocalMux I__2453 (
            .O(N__10385),
            .I(N__10360));
    LocalMux I__2452 (
            .O(N__10382),
            .I(N__10360));
    InMux I__2451 (
            .O(N__10381),
            .I(N__10357));
    InMux I__2450 (
            .O(N__10380),
            .I(N__10354));
    InMux I__2449 (
            .O(N__10379),
            .I(N__10351));
    Span4Mux_h I__2448 (
            .O(N__10376),
            .I(N__10343));
    LocalMux I__2447 (
            .O(N__10371),
            .I(N__10343));
    LocalMux I__2446 (
            .O(N__10368),
            .I(N__10343));
    InMux I__2445 (
            .O(N__10367),
            .I(N__10340));
    Span4Mux_v I__2444 (
            .O(N__10360),
            .I(N__10331));
    LocalMux I__2443 (
            .O(N__10357),
            .I(N__10331));
    LocalMux I__2442 (
            .O(N__10354),
            .I(N__10331));
    LocalMux I__2441 (
            .O(N__10351),
            .I(N__10331));
    InMux I__2440 (
            .O(N__10350),
            .I(N__10328));
    Span4Mux_v I__2439 (
            .O(N__10343),
            .I(N__10321));
    LocalMux I__2438 (
            .O(N__10340),
            .I(N__10321));
    Span4Mux_v I__2437 (
            .O(N__10331),
            .I(N__10316));
    LocalMux I__2436 (
            .O(N__10328),
            .I(N__10316));
    InMux I__2435 (
            .O(N__10327),
            .I(N__10313));
    CascadeMux I__2434 (
            .O(N__10326),
            .I(N__10310));
    Span4Mux_v I__2433 (
            .O(N__10321),
            .I(N__10307));
    Span4Mux_h I__2432 (
            .O(N__10316),
            .I(N__10304));
    LocalMux I__2431 (
            .O(N__10313),
            .I(N__10301));
    InMux I__2430 (
            .O(N__10310),
            .I(N__10298));
    Odrv4 I__2429 (
            .O(N__10307),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    Odrv4 I__2428 (
            .O(N__10304),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    Odrv12 I__2427 (
            .O(N__10301),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    LocalMux I__2426 (
            .O(N__10298),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    IoInMux I__2425 (
            .O(N__10289),
            .I(N__10286));
    LocalMux I__2424 (
            .O(N__10286),
            .I(N__10283));
    Span4Mux_s3_v I__2423 (
            .O(N__10283),
            .I(N__10280));
    Span4Mux_v I__2422 (
            .O(N__10280),
            .I(N__10277));
    Sp12to4 I__2421 (
            .O(N__10277),
            .I(N__10274));
    Odrv12 I__2420 (
            .O(N__10274),
            .I(un1_D_UU_AMIGA_7));
    InMux I__2419 (
            .O(N__10271),
            .I(N__10268));
    LocalMux I__2418 (
            .O(N__10268),
            .I(N__10265));
    Span12Mux_h I__2417 (
            .O(N__10265),
            .I(N__10262));
    Odrv12 I__2416 (
            .O(N__10262),
            .I(READ_CYCLE_ACTIVE_rep14_i_ess));
    IoInMux I__2415 (
            .O(N__10259),
            .I(N__10256));
    LocalMux I__2414 (
            .O(N__10256),
            .I(N__10253));
    IoSpan4Mux I__2413 (
            .O(N__10253),
            .I(N__10250));
    Span4Mux_s0_h I__2412 (
            .O(N__10250),
            .I(N__10247));
    Sp12to4 I__2411 (
            .O(N__10247),
            .I(N__10244));
    Odrv12 I__2410 (
            .O(N__10244),
            .I(N_219_i));
    InMux I__2409 (
            .O(N__10241),
            .I(N__10238));
    LocalMux I__2408 (
            .O(N__10238),
            .I(N__10235));
    Span4Mux_v I__2407 (
            .O(N__10235),
            .I(N__10232));
    Odrv4 I__2406 (
            .O(N__10232),
            .I(READ_CYCLE_ACTIVE_rep15_i_ess));
    IoInMux I__2405 (
            .O(N__10229),
            .I(N__10226));
    LocalMux I__2404 (
            .O(N__10226),
            .I(N__10223));
    Span4Mux_s1_h I__2403 (
            .O(N__10223),
            .I(N__10220));
    Sp12to4 I__2402 (
            .O(N__10220),
            .I(N__10217));
    Span12Mux_s11_v I__2401 (
            .O(N__10217),
            .I(N__10214));
    Span12Mux_h I__2400 (
            .O(N__10214),
            .I(N__10211));
    Odrv12 I__2399 (
            .O(N__10211),
            .I(N_220_i));
    InMux I__2398 (
            .O(N__10208),
            .I(N__10205));
    LocalMux I__2397 (
            .O(N__10205),
            .I(N__10202));
    Span12Mux_h I__2396 (
            .O(N__10202),
            .I(N__10199));
    Odrv12 I__2395 (
            .O(N__10199),
            .I(READ_CYCLE_ACTIVE_rep29_i_ess));
    IoInMux I__2394 (
            .O(N__10196),
            .I(N__10193));
    LocalMux I__2393 (
            .O(N__10193),
            .I(N__10190));
    Sp12to4 I__2392 (
            .O(N__10190),
            .I(N__10187));
    Span12Mux_h I__2391 (
            .O(N__10187),
            .I(N__10184));
    Odrv12 I__2390 (
            .O(N__10184),
            .I(N_234_i));
    IoInMux I__2389 (
            .O(N__10181),
            .I(N__10178));
    LocalMux I__2388 (
            .O(N__10178),
            .I(N__10175));
    IoSpan4Mux I__2387 (
            .O(N__10175),
            .I(N__10171));
    InMux I__2386 (
            .O(N__10174),
            .I(N__10168));
    IoSpan4Mux I__2385 (
            .O(N__10171),
            .I(N__10165));
    LocalMux I__2384 (
            .O(N__10168),
            .I(N__10162));
    Span4Mux_s2_h I__2383 (
            .O(N__10165),
            .I(N__10159));
    Span4Mux_v I__2382 (
            .O(N__10162),
            .I(N__10156));
    Sp12to4 I__2381 (
            .O(N__10159),
            .I(N__10153));
    Sp12to4 I__2380 (
            .O(N__10156),
            .I(N__10150));
    Span12Mux_h I__2379 (
            .O(N__10153),
            .I(N__10147));
    Span12Mux_h I__2378 (
            .O(N__10150),
            .I(N__10144));
    Span12Mux_h I__2377 (
            .O(N__10147),
            .I(N__10141));
    Span12Mux_v I__2376 (
            .O(N__10144),
            .I(N__10138));
    Odrv12 I__2375 (
            .O(N__10141),
            .I(D_LL_040_in_6));
    Odrv12 I__2374 (
            .O(N__10138),
            .I(D_LL_040_in_6));
    InMux I__2373 (
            .O(N__10133),
            .I(N__10130));
    LocalMux I__2372 (
            .O(N__10130),
            .I(N__10127));
    Span4Mux_v I__2371 (
            .O(N__10127),
            .I(N__10124));
    Sp12to4 I__2370 (
            .O(N__10124),
            .I(N__10121));
    Odrv12 I__2369 (
            .O(N__10121),
            .I(D_UM_040_in_6));
    IoInMux I__2368 (
            .O(N__10118),
            .I(N__10115));
    LocalMux I__2367 (
            .O(N__10115),
            .I(N__10112));
    Span4Mux_s0_h I__2366 (
            .O(N__10112),
            .I(N__10109));
    Span4Mux_h I__2365 (
            .O(N__10109),
            .I(N__10106));
    Sp12to4 I__2364 (
            .O(N__10106),
            .I(N__10103));
    Span12Mux_v I__2363 (
            .O(N__10103),
            .I(N__10100));
    Span12Mux_h I__2362 (
            .O(N__10100),
            .I(N__10097));
    Odrv12 I__2361 (
            .O(N__10097),
            .I(un1_D_UM_040_6));
    IoInMux I__2360 (
            .O(N__10094),
            .I(N__10091));
    LocalMux I__2359 (
            .O(N__10091),
            .I(N__10087));
    CascadeMux I__2358 (
            .O(N__10090),
            .I(N__10078));
    Span4Mux_s3_v I__2357 (
            .O(N__10087),
            .I(N__10074));
    InMux I__2356 (
            .O(N__10086),
            .I(N__10066));
    InMux I__2355 (
            .O(N__10085),
            .I(N__10066));
    InMux I__2354 (
            .O(N__10084),
            .I(N__10066));
    InMux I__2353 (
            .O(N__10083),
            .I(N__10059));
    InMux I__2352 (
            .O(N__10082),
            .I(N__10059));
    InMux I__2351 (
            .O(N__10081),
            .I(N__10059));
    InMux I__2350 (
            .O(N__10078),
            .I(N__10052));
    InMux I__2349 (
            .O(N__10077),
            .I(N__10052));
    Span4Mux_h I__2348 (
            .O(N__10074),
            .I(N__10044));
    CascadeMux I__2347 (
            .O(N__10073),
            .I(N__10035));
    LocalMux I__2346 (
            .O(N__10066),
            .I(N__10032));
    LocalMux I__2345 (
            .O(N__10059),
            .I(N__10029));
    InMux I__2344 (
            .O(N__10058),
            .I(N__10026));
    InMux I__2343 (
            .O(N__10057),
            .I(N__10023));
    LocalMux I__2342 (
            .O(N__10052),
            .I(N__10020));
    InMux I__2341 (
            .O(N__10051),
            .I(N__10015));
    InMux I__2340 (
            .O(N__10050),
            .I(N__10015));
    CascadeMux I__2339 (
            .O(N__10049),
            .I(N__9996));
    CascadeMux I__2338 (
            .O(N__10048),
            .I(N__9993));
    CascadeMux I__2337 (
            .O(N__10047),
            .I(N__9989));
    Span4Mux_h I__2336 (
            .O(N__10044),
            .I(N__9985));
    InMux I__2335 (
            .O(N__10043),
            .I(N__9980));
    InMux I__2334 (
            .O(N__10042),
            .I(N__9980));
    InMux I__2333 (
            .O(N__10041),
            .I(N__9975));
    InMux I__2332 (
            .O(N__10040),
            .I(N__9975));
    InMux I__2331 (
            .O(N__10039),
            .I(N__9972));
    InMux I__2330 (
            .O(N__10038),
            .I(N__9969));
    InMux I__2329 (
            .O(N__10035),
            .I(N__9966));
    Span4Mux_v I__2328 (
            .O(N__10032),
            .I(N__9957));
    Span4Mux_h I__2327 (
            .O(N__10029),
            .I(N__9957));
    LocalMux I__2326 (
            .O(N__10026),
            .I(N__9957));
    LocalMux I__2325 (
            .O(N__10023),
            .I(N__9957));
    Span4Mux_v I__2324 (
            .O(N__10020),
            .I(N__9952));
    LocalMux I__2323 (
            .O(N__10015),
            .I(N__9952));
    InMux I__2322 (
            .O(N__10014),
            .I(N__9949));
    CascadeMux I__2321 (
            .O(N__10013),
            .I(N__9946));
    CascadeMux I__2320 (
            .O(N__10012),
            .I(N__9943));
    CascadeMux I__2319 (
            .O(N__10011),
            .I(N__9940));
    InMux I__2318 (
            .O(N__10010),
            .I(N__9931));
    InMux I__2317 (
            .O(N__10009),
            .I(N__9931));
    InMux I__2316 (
            .O(N__10008),
            .I(N__9931));
    InMux I__2315 (
            .O(N__10007),
            .I(N__9914));
    InMux I__2314 (
            .O(N__10006),
            .I(N__9914));
    InMux I__2313 (
            .O(N__10005),
            .I(N__9914));
    InMux I__2312 (
            .O(N__10004),
            .I(N__9914));
    InMux I__2311 (
            .O(N__10003),
            .I(N__9914));
    InMux I__2310 (
            .O(N__10002),
            .I(N__9914));
    InMux I__2309 (
            .O(N__10001),
            .I(N__9914));
    InMux I__2308 (
            .O(N__10000),
            .I(N__9914));
    InMux I__2307 (
            .O(N__9999),
            .I(N__9901));
    InMux I__2306 (
            .O(N__9996),
            .I(N__9901));
    InMux I__2305 (
            .O(N__9993),
            .I(N__9901));
    InMux I__2304 (
            .O(N__9992),
            .I(N__9901));
    InMux I__2303 (
            .O(N__9989),
            .I(N__9901));
    InMux I__2302 (
            .O(N__9988),
            .I(N__9901));
    Span4Mux_v I__2301 (
            .O(N__9985),
            .I(N__9884));
    LocalMux I__2300 (
            .O(N__9980),
            .I(N__9884));
    LocalMux I__2299 (
            .O(N__9975),
            .I(N__9884));
    LocalMux I__2298 (
            .O(N__9972),
            .I(N__9884));
    LocalMux I__2297 (
            .O(N__9969),
            .I(N__9884));
    LocalMux I__2296 (
            .O(N__9966),
            .I(N__9881));
    Span4Mux_v I__2295 (
            .O(N__9957),
            .I(N__9874));
    Span4Mux_h I__2294 (
            .O(N__9952),
            .I(N__9874));
    LocalMux I__2293 (
            .O(N__9949),
            .I(N__9874));
    InMux I__2292 (
            .O(N__9946),
            .I(N__9865));
    InMux I__2291 (
            .O(N__9943),
            .I(N__9865));
    InMux I__2290 (
            .O(N__9940),
            .I(N__9865));
    InMux I__2289 (
            .O(N__9939),
            .I(N__9865));
    CascadeMux I__2288 (
            .O(N__9938),
            .I(N__9861));
    LocalMux I__2287 (
            .O(N__9931),
            .I(N__9857));
    LocalMux I__2286 (
            .O(N__9914),
            .I(N__9852));
    LocalMux I__2285 (
            .O(N__9901),
            .I(N__9852));
    CascadeMux I__2284 (
            .O(N__9900),
            .I(N__9847));
    CascadeMux I__2283 (
            .O(N__9899),
            .I(N__9843));
    CascadeMux I__2282 (
            .O(N__9898),
            .I(N__9831));
    CascadeMux I__2281 (
            .O(N__9897),
            .I(N__9827));
    CascadeMux I__2280 (
            .O(N__9896),
            .I(N__9824));
    CascadeMux I__2279 (
            .O(N__9895),
            .I(N__9820));
    Span4Mux_v I__2278 (
            .O(N__9884),
            .I(N__9814));
    Span4Mux_v I__2277 (
            .O(N__9881),
            .I(N__9814));
    Span4Mux_h I__2276 (
            .O(N__9874),
            .I(N__9809));
    LocalMux I__2275 (
            .O(N__9865),
            .I(N__9809));
    InMux I__2274 (
            .O(N__9864),
            .I(N__9802));
    InMux I__2273 (
            .O(N__9861),
            .I(N__9802));
    InMux I__2272 (
            .O(N__9860),
            .I(N__9802));
    Span4Mux_v I__2271 (
            .O(N__9857),
            .I(N__9797));
    Span4Mux_v I__2270 (
            .O(N__9852),
            .I(N__9797));
    InMux I__2269 (
            .O(N__9851),
            .I(N__9784));
    InMux I__2268 (
            .O(N__9850),
            .I(N__9784));
    InMux I__2267 (
            .O(N__9847),
            .I(N__9784));
    InMux I__2266 (
            .O(N__9846),
            .I(N__9784));
    InMux I__2265 (
            .O(N__9843),
            .I(N__9784));
    InMux I__2264 (
            .O(N__9842),
            .I(N__9784));
    InMux I__2263 (
            .O(N__9841),
            .I(N__9767));
    InMux I__2262 (
            .O(N__9840),
            .I(N__9767));
    InMux I__2261 (
            .O(N__9839),
            .I(N__9767));
    InMux I__2260 (
            .O(N__9838),
            .I(N__9767));
    InMux I__2259 (
            .O(N__9837),
            .I(N__9767));
    InMux I__2258 (
            .O(N__9836),
            .I(N__9767));
    InMux I__2257 (
            .O(N__9835),
            .I(N__9767));
    InMux I__2256 (
            .O(N__9834),
            .I(N__9767));
    InMux I__2255 (
            .O(N__9831),
            .I(N__9752));
    InMux I__2254 (
            .O(N__9830),
            .I(N__9752));
    InMux I__2253 (
            .O(N__9827),
            .I(N__9752));
    InMux I__2252 (
            .O(N__9824),
            .I(N__9752));
    InMux I__2251 (
            .O(N__9823),
            .I(N__9752));
    InMux I__2250 (
            .O(N__9820),
            .I(N__9752));
    InMux I__2249 (
            .O(N__9819),
            .I(N__9752));
    Span4Mux_h I__2248 (
            .O(N__9814),
            .I(N__9747));
    Span4Mux_v I__2247 (
            .O(N__9809),
            .I(N__9747));
    LocalMux I__2246 (
            .O(N__9802),
            .I(N__9744));
    Sp12to4 I__2245 (
            .O(N__9797),
            .I(N__9733));
    LocalMux I__2244 (
            .O(N__9784),
            .I(N__9733));
    LocalMux I__2243 (
            .O(N__9767),
            .I(N__9733));
    LocalMux I__2242 (
            .O(N__9752),
            .I(N__9733));
    Sp12to4 I__2241 (
            .O(N__9747),
            .I(N__9733));
    Span12Mux_v I__2240 (
            .O(N__9744),
            .I(N__9730));
    Span12Mux_h I__2239 (
            .O(N__9733),
            .I(N__9727));
    Span12Mux_h I__2238 (
            .O(N__9730),
            .I(N__9724));
    Odrv12 I__2237 (
            .O(N__9727),
            .I(RnW_c));
    Odrv12 I__2236 (
            .O(N__9724),
            .I(RnW_c));
    InMux I__2235 (
            .O(N__9719),
            .I(N__9710));
    InMux I__2234 (
            .O(N__9718),
            .I(N__9710));
    InMux I__2233 (
            .O(N__9717),
            .I(N__9710));
    LocalMux I__2232 (
            .O(N__9710),
            .I(N__9687));
    InMux I__2231 (
            .O(N__9709),
            .I(N__9684));
    InMux I__2230 (
            .O(N__9708),
            .I(N__9676));
    InMux I__2229 (
            .O(N__9707),
            .I(N__9671));
    InMux I__2228 (
            .O(N__9706),
            .I(N__9664));
    InMux I__2227 (
            .O(N__9705),
            .I(N__9664));
    InMux I__2226 (
            .O(N__9704),
            .I(N__9664));
    InMux I__2225 (
            .O(N__9703),
            .I(N__9655));
    InMux I__2224 (
            .O(N__9702),
            .I(N__9655));
    InMux I__2223 (
            .O(N__9701),
            .I(N__9655));
    InMux I__2222 (
            .O(N__9700),
            .I(N__9655));
    InMux I__2221 (
            .O(N__9699),
            .I(N__9652));
    InMux I__2220 (
            .O(N__9698),
            .I(N__9649));
    InMux I__2219 (
            .O(N__9697),
            .I(N__9639));
    InMux I__2218 (
            .O(N__9696),
            .I(N__9632));
    InMux I__2217 (
            .O(N__9695),
            .I(N__9632));
    InMux I__2216 (
            .O(N__9694),
            .I(N__9632));
    InMux I__2215 (
            .O(N__9693),
            .I(N__9627));
    InMux I__2214 (
            .O(N__9692),
            .I(N__9627));
    InMux I__2213 (
            .O(N__9691),
            .I(N__9622));
    InMux I__2212 (
            .O(N__9690),
            .I(N__9622));
    Span4Mux_v I__2211 (
            .O(N__9687),
            .I(N__9603));
    LocalMux I__2210 (
            .O(N__9684),
            .I(N__9603));
    InMux I__2209 (
            .O(N__9683),
            .I(N__9598));
    InMux I__2208 (
            .O(N__9682),
            .I(N__9598));
    InMux I__2207 (
            .O(N__9681),
            .I(N__9591));
    InMux I__2206 (
            .O(N__9680),
            .I(N__9591));
    InMux I__2205 (
            .O(N__9679),
            .I(N__9591));
    LocalMux I__2204 (
            .O(N__9676),
            .I(N__9588));
    InMux I__2203 (
            .O(N__9675),
            .I(N__9583));
    InMux I__2202 (
            .O(N__9674),
            .I(N__9583));
    LocalMux I__2201 (
            .O(N__9671),
            .I(N__9564));
    LocalMux I__2200 (
            .O(N__9664),
            .I(N__9559));
    LocalMux I__2199 (
            .O(N__9655),
            .I(N__9559));
    LocalMux I__2198 (
            .O(N__9652),
            .I(N__9554));
    LocalMux I__2197 (
            .O(N__9649),
            .I(N__9554));
    InMux I__2196 (
            .O(N__9648),
            .I(N__9539));
    InMux I__2195 (
            .O(N__9647),
            .I(N__9539));
    InMux I__2194 (
            .O(N__9646),
            .I(N__9539));
    InMux I__2193 (
            .O(N__9645),
            .I(N__9539));
    InMux I__2192 (
            .O(N__9644),
            .I(N__9539));
    InMux I__2191 (
            .O(N__9643),
            .I(N__9539));
    InMux I__2190 (
            .O(N__9642),
            .I(N__9539));
    LocalMux I__2189 (
            .O(N__9639),
            .I(N__9534));
    LocalMux I__2188 (
            .O(N__9632),
            .I(N__9534));
    LocalMux I__2187 (
            .O(N__9627),
            .I(N__9531));
    LocalMux I__2186 (
            .O(N__9622),
            .I(N__9528));
    InMux I__2185 (
            .O(N__9621),
            .I(N__9515));
    InMux I__2184 (
            .O(N__9620),
            .I(N__9515));
    InMux I__2183 (
            .O(N__9619),
            .I(N__9515));
    InMux I__2182 (
            .O(N__9618),
            .I(N__9515));
    InMux I__2181 (
            .O(N__9617),
            .I(N__9515));
    InMux I__2180 (
            .O(N__9616),
            .I(N__9515));
    InMux I__2179 (
            .O(N__9615),
            .I(N__9498));
    InMux I__2178 (
            .O(N__9614),
            .I(N__9498));
    InMux I__2177 (
            .O(N__9613),
            .I(N__9498));
    InMux I__2176 (
            .O(N__9612),
            .I(N__9498));
    InMux I__2175 (
            .O(N__9611),
            .I(N__9498));
    InMux I__2174 (
            .O(N__9610),
            .I(N__9498));
    InMux I__2173 (
            .O(N__9609),
            .I(N__9498));
    InMux I__2172 (
            .O(N__9608),
            .I(N__9498));
    Span4Mux_v I__2171 (
            .O(N__9603),
            .I(N__9487));
    LocalMux I__2170 (
            .O(N__9598),
            .I(N__9487));
    LocalMux I__2169 (
            .O(N__9591),
            .I(N__9487));
    Span4Mux_h I__2168 (
            .O(N__9588),
            .I(N__9487));
    LocalMux I__2167 (
            .O(N__9583),
            .I(N__9487));
    InMux I__2166 (
            .O(N__9582),
            .I(N__9470));
    InMux I__2165 (
            .O(N__9581),
            .I(N__9470));
    InMux I__2164 (
            .O(N__9580),
            .I(N__9470));
    InMux I__2163 (
            .O(N__9579),
            .I(N__9470));
    InMux I__2162 (
            .O(N__9578),
            .I(N__9470));
    InMux I__2161 (
            .O(N__9577),
            .I(N__9470));
    InMux I__2160 (
            .O(N__9576),
            .I(N__9470));
    InMux I__2159 (
            .O(N__9575),
            .I(N__9470));
    InMux I__2158 (
            .O(N__9574),
            .I(N__9457));
    InMux I__2157 (
            .O(N__9573),
            .I(N__9457));
    InMux I__2156 (
            .O(N__9572),
            .I(N__9457));
    InMux I__2155 (
            .O(N__9571),
            .I(N__9457));
    InMux I__2154 (
            .O(N__9570),
            .I(N__9457));
    InMux I__2153 (
            .O(N__9569),
            .I(N__9457));
    InMux I__2152 (
            .O(N__9568),
            .I(N__9454));
    InMux I__2151 (
            .O(N__9567),
            .I(N__9451));
    Odrv4 I__2150 (
            .O(N__9564),
            .I(\U111_CYCLE_SM.N_44 ));
    Odrv12 I__2149 (
            .O(N__9559),
            .I(\U111_CYCLE_SM.N_44 ));
    Odrv4 I__2148 (
            .O(N__9554),
            .I(\U111_CYCLE_SM.N_44 ));
    LocalMux I__2147 (
            .O(N__9539),
            .I(\U111_CYCLE_SM.N_44 ));
    Odrv12 I__2146 (
            .O(N__9534),
            .I(\U111_CYCLE_SM.N_44 ));
    Odrv4 I__2145 (
            .O(N__9531),
            .I(\U111_CYCLE_SM.N_44 ));
    Odrv4 I__2144 (
            .O(N__9528),
            .I(\U111_CYCLE_SM.N_44 ));
    LocalMux I__2143 (
            .O(N__9515),
            .I(\U111_CYCLE_SM.N_44 ));
    LocalMux I__2142 (
            .O(N__9498),
            .I(\U111_CYCLE_SM.N_44 ));
    Odrv4 I__2141 (
            .O(N__9487),
            .I(\U111_CYCLE_SM.N_44 ));
    LocalMux I__2140 (
            .O(N__9470),
            .I(\U111_CYCLE_SM.N_44 ));
    LocalMux I__2139 (
            .O(N__9457),
            .I(\U111_CYCLE_SM.N_44 ));
    LocalMux I__2138 (
            .O(N__9454),
            .I(\U111_CYCLE_SM.N_44 ));
    LocalMux I__2137 (
            .O(N__9451),
            .I(\U111_CYCLE_SM.N_44 ));
    InMux I__2136 (
            .O(N__9422),
            .I(N__9419));
    LocalMux I__2135 (
            .O(N__9419),
            .I(N__9413));
    ClkMux I__2134 (
            .O(N__9418),
            .I(N__9317));
    ClkMux I__2133 (
            .O(N__9417),
            .I(N__9317));
    ClkMux I__2132 (
            .O(N__9416),
            .I(N__9317));
    Glb2LocalMux I__2131 (
            .O(N__9413),
            .I(N__9317));
    ClkMux I__2130 (
            .O(N__9412),
            .I(N__9317));
    ClkMux I__2129 (
            .O(N__9411),
            .I(N__9317));
    ClkMux I__2128 (
            .O(N__9410),
            .I(N__9317));
    ClkMux I__2127 (
            .O(N__9409),
            .I(N__9317));
    ClkMux I__2126 (
            .O(N__9408),
            .I(N__9317));
    ClkMux I__2125 (
            .O(N__9407),
            .I(N__9317));
    ClkMux I__2124 (
            .O(N__9406),
            .I(N__9317));
    ClkMux I__2123 (
            .O(N__9405),
            .I(N__9317));
    ClkMux I__2122 (
            .O(N__9404),
            .I(N__9317));
    ClkMux I__2121 (
            .O(N__9403),
            .I(N__9317));
    ClkMux I__2120 (
            .O(N__9402),
            .I(N__9317));
    ClkMux I__2119 (
            .O(N__9401),
            .I(N__9317));
    ClkMux I__2118 (
            .O(N__9400),
            .I(N__9317));
    ClkMux I__2117 (
            .O(N__9399),
            .I(N__9317));
    ClkMux I__2116 (
            .O(N__9398),
            .I(N__9317));
    ClkMux I__2115 (
            .O(N__9397),
            .I(N__9317));
    ClkMux I__2114 (
            .O(N__9396),
            .I(N__9317));
    ClkMux I__2113 (
            .O(N__9395),
            .I(N__9317));
    ClkMux I__2112 (
            .O(N__9394),
            .I(N__9317));
    ClkMux I__2111 (
            .O(N__9393),
            .I(N__9317));
    ClkMux I__2110 (
            .O(N__9392),
            .I(N__9317));
    ClkMux I__2109 (
            .O(N__9391),
            .I(N__9317));
    ClkMux I__2108 (
            .O(N__9390),
            .I(N__9317));
    ClkMux I__2107 (
            .O(N__9389),
            .I(N__9317));
    ClkMux I__2106 (
            .O(N__9388),
            .I(N__9317));
    ClkMux I__2105 (
            .O(N__9387),
            .I(N__9317));
    ClkMux I__2104 (
            .O(N__9386),
            .I(N__9317));
    ClkMux I__2103 (
            .O(N__9385),
            .I(N__9317));
    ClkMux I__2102 (
            .O(N__9384),
            .I(N__9317));
    GlobalMux I__2101 (
            .O(N__9317),
            .I(CLK40));
    CEMux I__2100 (
            .O(N__9314),
            .I(N__9257));
    CEMux I__2099 (
            .O(N__9313),
            .I(N__9257));
    CEMux I__2098 (
            .O(N__9312),
            .I(N__9257));
    CEMux I__2097 (
            .O(N__9311),
            .I(N__9257));
    CEMux I__2096 (
            .O(N__9310),
            .I(N__9257));
    CEMux I__2095 (
            .O(N__9309),
            .I(N__9257));
    CEMux I__2094 (
            .O(N__9308),
            .I(N__9257));
    CEMux I__2093 (
            .O(N__9307),
            .I(N__9257));
    CEMux I__2092 (
            .O(N__9306),
            .I(N__9257));
    CEMux I__2091 (
            .O(N__9305),
            .I(N__9257));
    CEMux I__2090 (
            .O(N__9304),
            .I(N__9257));
    CEMux I__2089 (
            .O(N__9303),
            .I(N__9257));
    CEMux I__2088 (
            .O(N__9302),
            .I(N__9257));
    CEMux I__2087 (
            .O(N__9301),
            .I(N__9257));
    CEMux I__2086 (
            .O(N__9300),
            .I(N__9257));
    CEMux I__2085 (
            .O(N__9299),
            .I(N__9257));
    CEMux I__2084 (
            .O(N__9298),
            .I(N__9257));
    CEMux I__2083 (
            .O(N__9297),
            .I(N__9257));
    CEMux I__2082 (
            .O(N__9296),
            .I(N__9257));
    GlobalMux I__2081 (
            .O(N__9257),
            .I(N__9254));
    gio2CtrlBuf I__2080 (
            .O(N__9254),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_g_0 ));
    InMux I__2079 (
            .O(N__9251),
            .I(N__9248));
    LocalMux I__2078 (
            .O(N__9248),
            .I(N__9221));
    SRMux I__2077 (
            .O(N__9247),
            .I(N__9170));
    SRMux I__2076 (
            .O(N__9246),
            .I(N__9170));
    SRMux I__2075 (
            .O(N__9245),
            .I(N__9170));
    SRMux I__2074 (
            .O(N__9244),
            .I(N__9170));
    SRMux I__2073 (
            .O(N__9243),
            .I(N__9170));
    SRMux I__2072 (
            .O(N__9242),
            .I(N__9170));
    SRMux I__2071 (
            .O(N__9241),
            .I(N__9170));
    SRMux I__2070 (
            .O(N__9240),
            .I(N__9170));
    SRMux I__2069 (
            .O(N__9239),
            .I(N__9170));
    SRMux I__2068 (
            .O(N__9238),
            .I(N__9170));
    SRMux I__2067 (
            .O(N__9237),
            .I(N__9170));
    SRMux I__2066 (
            .O(N__9236),
            .I(N__9170));
    SRMux I__2065 (
            .O(N__9235),
            .I(N__9170));
    SRMux I__2064 (
            .O(N__9234),
            .I(N__9170));
    SRMux I__2063 (
            .O(N__9233),
            .I(N__9170));
    SRMux I__2062 (
            .O(N__9232),
            .I(N__9170));
    SRMux I__2061 (
            .O(N__9231),
            .I(N__9170));
    SRMux I__2060 (
            .O(N__9230),
            .I(N__9170));
    SRMux I__2059 (
            .O(N__9229),
            .I(N__9170));
    SRMux I__2058 (
            .O(N__9228),
            .I(N__9170));
    SRMux I__2057 (
            .O(N__9227),
            .I(N__9170));
    SRMux I__2056 (
            .O(N__9226),
            .I(N__9170));
    SRMux I__2055 (
            .O(N__9225),
            .I(N__9170));
    SRMux I__2054 (
            .O(N__9224),
            .I(N__9170));
    Glb2LocalMux I__2053 (
            .O(N__9221),
            .I(N__9170));
    GlobalMux I__2052 (
            .O(N__9170),
            .I(N__9167));
    gio2CtrlBuf I__2051 (
            .O(N__9167),
            .I(RESETn_c_i_g));
    InMux I__2050 (
            .O(N__9164),
            .I(N__9161));
    LocalMux I__2049 (
            .O(N__9161),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ));
    InMux I__2048 (
            .O(N__9158),
            .I(N__9155));
    LocalMux I__2047 (
            .O(N__9155),
            .I(N__9152));
    Span4Mux_v I__2046 (
            .O(N__9152),
            .I(N__9149));
    Span4Mux_v I__2045 (
            .O(N__9149),
            .I(N__9146));
    Span4Mux_v I__2044 (
            .O(N__9146),
            .I(N__9141));
    InMux I__2043 (
            .O(N__9145),
            .I(N__9138));
    InMux I__2042 (
            .O(N__9144),
            .I(N__9135));
    Sp12to4 I__2041 (
            .O(N__9141),
            .I(N__9128));
    LocalMux I__2040 (
            .O(N__9138),
            .I(N__9128));
    LocalMux I__2039 (
            .O(N__9135),
            .I(N__9128));
    Span12Mux_h I__2038 (
            .O(N__9128),
            .I(N__9125));
    Odrv12 I__2037 (
            .O(N__9125),
            .I(D_UM_AMIGA_in_0));
    IoInMux I__2036 (
            .O(N__9122),
            .I(N__9119));
    LocalMux I__2035 (
            .O(N__9119),
            .I(N__9116));
    IoSpan4Mux I__2034 (
            .O(N__9116),
            .I(N__9113));
    Span4Mux_s3_h I__2033 (
            .O(N__9113),
            .I(N__9110));
    Span4Mux_h I__2032 (
            .O(N__9110),
            .I(N__9107));
    Span4Mux_h I__2031 (
            .O(N__9107),
            .I(N__9104));
    Odrv4 I__2030 (
            .O(N__9104),
            .I(un1_D_UM_AMIGA_0));
    InMux I__2029 (
            .O(N__9101),
            .I(N__9098));
    LocalMux I__2028 (
            .O(N__9098),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ));
    InMux I__2027 (
            .O(N__9095),
            .I(N__9091));
    InMux I__2026 (
            .O(N__9094),
            .I(N__9087));
    LocalMux I__2025 (
            .O(N__9091),
            .I(N__9084));
    InMux I__2024 (
            .O(N__9090),
            .I(N__9081));
    LocalMux I__2023 (
            .O(N__9087),
            .I(N__9078));
    Span4Mux_v I__2022 (
            .O(N__9084),
            .I(N__9075));
    LocalMux I__2021 (
            .O(N__9081),
            .I(N__9072));
    Span4Mux_v I__2020 (
            .O(N__9078),
            .I(N__9069));
    Span4Mux_v I__2019 (
            .O(N__9075),
            .I(N__9064));
    Span4Mux_v I__2018 (
            .O(N__9072),
            .I(N__9064));
    Sp12to4 I__2017 (
            .O(N__9069),
            .I(N__9059));
    Sp12to4 I__2016 (
            .O(N__9064),
            .I(N__9059));
    Span12Mux_h I__2015 (
            .O(N__9059),
            .I(N__9056));
    Span12Mux_v I__2014 (
            .O(N__9056),
            .I(N__9053));
    Odrv12 I__2013 (
            .O(N__9053),
            .I(D_UM_AMIGA_in_6));
    IoInMux I__2012 (
            .O(N__9050),
            .I(N__9047));
    LocalMux I__2011 (
            .O(N__9047),
            .I(N__9044));
    Span12Mux_s6_h I__2010 (
            .O(N__9044),
            .I(N__9041));
    Odrv12 I__2009 (
            .O(N__9041),
            .I(un1_D_UM_AMIGA_6));
    InMux I__2008 (
            .O(N__9038),
            .I(N__9035));
    LocalMux I__2007 (
            .O(N__9035),
            .I(N__9032));
    Odrv4 I__2006 (
            .O(N__9032),
            .I(READ_CYCLE_ACTIVE_rep19_i_ess));
    InMux I__2005 (
            .O(N__9029),
            .I(N__9026));
    LocalMux I__2004 (
            .O(N__9026),
            .I(N__9021));
    InMux I__2003 (
            .O(N__9025),
            .I(N__9018));
    InMux I__2002 (
            .O(N__9024),
            .I(N__9015));
    Span4Mux_v I__2001 (
            .O(N__9021),
            .I(N__9012));
    LocalMux I__2000 (
            .O(N__9018),
            .I(N__9009));
    LocalMux I__1999 (
            .O(N__9015),
            .I(N__9006));
    Sp12to4 I__1998 (
            .O(N__9012),
            .I(N__9003));
    Span4Mux_v I__1997 (
            .O(N__9009),
            .I(N__9000));
    Span4Mux_v I__1996 (
            .O(N__9006),
            .I(N__8997));
    Span12Mux_h I__1995 (
            .O(N__9003),
            .I(N__8994));
    Sp12to4 I__1994 (
            .O(N__9000),
            .I(N__8989));
    Sp12to4 I__1993 (
            .O(N__8997),
            .I(N__8989));
    Span12Mux_v I__1992 (
            .O(N__8994),
            .I(N__8986));
    Span12Mux_h I__1991 (
            .O(N__8989),
            .I(N__8983));
    Odrv12 I__1990 (
            .O(N__8986),
            .I(D_UM_AMIGA_in_1));
    Odrv12 I__1989 (
            .O(N__8983),
            .I(D_UM_AMIGA_in_1));
    InMux I__1988 (
            .O(N__8978),
            .I(N__8975));
    LocalMux I__1987 (
            .O(N__8975),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ));
    IoInMux I__1986 (
            .O(N__8972),
            .I(N__8969));
    LocalMux I__1985 (
            .O(N__8969),
            .I(N__8966));
    Span4Mux_s2_h I__1984 (
            .O(N__8966),
            .I(N__8963));
    Sp12to4 I__1983 (
            .O(N__8963),
            .I(N__8960));
    Span12Mux_v I__1982 (
            .O(N__8960),
            .I(N__8957));
    Span12Mux_h I__1981 (
            .O(N__8957),
            .I(N__8954));
    Odrv12 I__1980 (
            .O(N__8954),
            .I(un1_D_UM_AMIGA_1));
    InMux I__1979 (
            .O(N__8951),
            .I(N__8948));
    LocalMux I__1978 (
            .O(N__8948),
            .I(N__8945));
    Span4Mux_v I__1977 (
            .O(N__8945),
            .I(N__8942));
    Odrv4 I__1976 (
            .O(N__8942),
            .I(READ_CYCLE_ACTIVE_rep11_i_ess));
    IoInMux I__1975 (
            .O(N__8939),
            .I(N__8936));
    LocalMux I__1974 (
            .O(N__8936),
            .I(N__8933));
    Span12Mux_s2_h I__1973 (
            .O(N__8933),
            .I(N__8930));
    Span12Mux_h I__1972 (
            .O(N__8930),
            .I(N__8927));
    Odrv12 I__1971 (
            .O(N__8927),
            .I(N_216_i));
    IoInMux I__1970 (
            .O(N__8924),
            .I(N__8921));
    LocalMux I__1969 (
            .O(N__8921),
            .I(N__8917));
    InMux I__1968 (
            .O(N__8920),
            .I(N__8914));
    Span4Mux_s3_h I__1967 (
            .O(N__8917),
            .I(N__8911));
    LocalMux I__1966 (
            .O(N__8914),
            .I(N__8908));
    Span4Mux_h I__1965 (
            .O(N__8911),
            .I(N__8905));
    Span4Mux_h I__1964 (
            .O(N__8908),
            .I(N__8902));
    Sp12to4 I__1963 (
            .O(N__8905),
            .I(N__8899));
    Sp12to4 I__1962 (
            .O(N__8902),
            .I(N__8896));
    Span12Mux_v I__1961 (
            .O(N__8899),
            .I(N__8893));
    Span12Mux_v I__1960 (
            .O(N__8896),
            .I(N__8890));
    Span12Mux_h I__1959 (
            .O(N__8893),
            .I(N__8885));
    Span12Mux_v I__1958 (
            .O(N__8890),
            .I(N__8885));
    Span12Mux_h I__1957 (
            .O(N__8885),
            .I(N__8882));
    Odrv12 I__1956 (
            .O(N__8882),
            .I(D_LM_040_in_1));
    InMux I__1955 (
            .O(N__8879),
            .I(N__8876));
    LocalMux I__1954 (
            .O(N__8876),
            .I(N__8873));
    Span4Mux_v I__1953 (
            .O(N__8873),
            .I(N__8870));
    Span4Mux_v I__1952 (
            .O(N__8870),
            .I(N__8867));
    Sp12to4 I__1951 (
            .O(N__8867),
            .I(N__8864));
    Span12Mux_h I__1950 (
            .O(N__8864),
            .I(N__8861));
    Odrv12 I__1949 (
            .O(N__8861),
            .I(D_UU_040_in_1));
    IoInMux I__1948 (
            .O(N__8858),
            .I(N__8855));
    LocalMux I__1947 (
            .O(N__8855),
            .I(N__8852));
    Span4Mux_s1_h I__1946 (
            .O(N__8852),
            .I(N__8849));
    Span4Mux_h I__1945 (
            .O(N__8849),
            .I(N__8846));
    Span4Mux_h I__1944 (
            .O(N__8846),
            .I(N__8843));
    Span4Mux_h I__1943 (
            .O(N__8843),
            .I(N__8840));
    Span4Mux_h I__1942 (
            .O(N__8840),
            .I(N__8837));
    Odrv4 I__1941 (
            .O(N__8837),
            .I(un1_D_UU_040_1));
    InMux I__1940 (
            .O(N__8834),
            .I(N__8831));
    LocalMux I__1939 (
            .O(N__8831),
            .I(N__8828));
    Odrv12 I__1938 (
            .O(N__8828),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ));
    InMux I__1937 (
            .O(N__8825),
            .I(N__8820));
    InMux I__1936 (
            .O(N__8824),
            .I(N__8817));
    InMux I__1935 (
            .O(N__8823),
            .I(N__8814));
    LocalMux I__1934 (
            .O(N__8820),
            .I(N__8811));
    LocalMux I__1933 (
            .O(N__8817),
            .I(N__8808));
    LocalMux I__1932 (
            .O(N__8814),
            .I(N__8805));
    Span4Mux_v I__1931 (
            .O(N__8811),
            .I(N__8800));
    Span4Mux_v I__1930 (
            .O(N__8808),
            .I(N__8800));
    Span4Mux_v I__1929 (
            .O(N__8805),
            .I(N__8797));
    Sp12to4 I__1928 (
            .O(N__8800),
            .I(N__8792));
    Sp12to4 I__1927 (
            .O(N__8797),
            .I(N__8792));
    Span12Mux_h I__1926 (
            .O(N__8792),
            .I(N__8789));
    Odrv12 I__1925 (
            .O(N__8789),
            .I(D_UU_AMIGA_in_6));
    IoInMux I__1924 (
            .O(N__8786),
            .I(N__8783));
    LocalMux I__1923 (
            .O(N__8783),
            .I(N__8780));
    Span12Mux_s8_v I__1922 (
            .O(N__8780),
            .I(N__8777));
    Odrv12 I__1921 (
            .O(N__8777),
            .I(un1_D_UU_AMIGA_6));
    InMux I__1920 (
            .O(N__8774),
            .I(N__8771));
    LocalMux I__1919 (
            .O(N__8771),
            .I(N__8768));
    Odrv12 I__1918 (
            .O(N__8768),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ));
    InMux I__1917 (
            .O(N__8765),
            .I(N__8762));
    LocalMux I__1916 (
            .O(N__8762),
            .I(N__8757));
    InMux I__1915 (
            .O(N__8761),
            .I(N__8754));
    InMux I__1914 (
            .O(N__8760),
            .I(N__8751));
    Span4Mux_v I__1913 (
            .O(N__8757),
            .I(N__8748));
    LocalMux I__1912 (
            .O(N__8754),
            .I(N__8745));
    LocalMux I__1911 (
            .O(N__8751),
            .I(N__8742));
    Span4Mux_h I__1910 (
            .O(N__8748),
            .I(N__8739));
    Span4Mux_v I__1909 (
            .O(N__8745),
            .I(N__8736));
    Span4Mux_h I__1908 (
            .O(N__8742),
            .I(N__8733));
    Sp12to4 I__1907 (
            .O(N__8739),
            .I(N__8728));
    Sp12to4 I__1906 (
            .O(N__8736),
            .I(N__8728));
    Sp12to4 I__1905 (
            .O(N__8733),
            .I(N__8725));
    Span12Mux_h I__1904 (
            .O(N__8728),
            .I(N__8722));
    Span12Mux_v I__1903 (
            .O(N__8725),
            .I(N__8719));
    Span12Mux_v I__1902 (
            .O(N__8722),
            .I(N__8714));
    Span12Mux_h I__1901 (
            .O(N__8719),
            .I(N__8714));
    Odrv12 I__1900 (
            .O(N__8714),
            .I(D_UU_AMIGA_in_3));
    IoInMux I__1899 (
            .O(N__8711),
            .I(N__8708));
    LocalMux I__1898 (
            .O(N__8708),
            .I(N__8705));
    IoSpan4Mux I__1897 (
            .O(N__8705),
            .I(N__8702));
    IoSpan4Mux I__1896 (
            .O(N__8702),
            .I(N__8699));
    Span4Mux_s3_v I__1895 (
            .O(N__8699),
            .I(N__8696));
    Span4Mux_h I__1894 (
            .O(N__8696),
            .I(N__8693));
    Span4Mux_v I__1893 (
            .O(N__8693),
            .I(N__8690));
    Odrv4 I__1892 (
            .O(N__8690),
            .I(un1_D_UU_AMIGA_3));
    InMux I__1891 (
            .O(N__8687),
            .I(N__8683));
    InMux I__1890 (
            .O(N__8686),
            .I(N__8679));
    LocalMux I__1889 (
            .O(N__8683),
            .I(N__8676));
    InMux I__1888 (
            .O(N__8682),
            .I(N__8673));
    LocalMux I__1887 (
            .O(N__8679),
            .I(N__8670));
    Span12Mux_v I__1886 (
            .O(N__8676),
            .I(N__8665));
    LocalMux I__1885 (
            .O(N__8673),
            .I(N__8665));
    Span4Mux_v I__1884 (
            .O(N__8670),
            .I(N__8662));
    Span12Mux_v I__1883 (
            .O(N__8665),
            .I(N__8659));
    Sp12to4 I__1882 (
            .O(N__8662),
            .I(N__8656));
    Span12Mux_h I__1881 (
            .O(N__8659),
            .I(N__8653));
    Span12Mux_h I__1880 (
            .O(N__8656),
            .I(N__8650));
    Odrv12 I__1879 (
            .O(N__8653),
            .I(D_UM_AMIGA_in_7));
    Odrv12 I__1878 (
            .O(N__8650),
            .I(D_UM_AMIGA_in_7));
    InMux I__1877 (
            .O(N__8645),
            .I(N__8642));
    LocalMux I__1876 (
            .O(N__8642),
            .I(N__8639));
    Span4Mux_v I__1875 (
            .O(N__8639),
            .I(N__8636));
    Odrv4 I__1874 (
            .O(N__8636),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ));
    IoInMux I__1873 (
            .O(N__8633),
            .I(N__8630));
    LocalMux I__1872 (
            .O(N__8630),
            .I(N__8627));
    Span12Mux_s3_h I__1871 (
            .O(N__8627),
            .I(N__8624));
    Span12Mux_h I__1870 (
            .O(N__8624),
            .I(N__8621));
    Odrv12 I__1869 (
            .O(N__8621),
            .I(un1_D_UM_AMIGA_7));
    InMux I__1868 (
            .O(N__8618),
            .I(N__8615));
    LocalMux I__1867 (
            .O(N__8615),
            .I(N__8612));
    Span12Mux_s7_v I__1866 (
            .O(N__8612),
            .I(N__8609));
    Span12Mux_h I__1865 (
            .O(N__8609),
            .I(N__8606));
    Odrv12 I__1864 (
            .O(N__8606),
            .I(D_UU_040_in_7));
    IoInMux I__1863 (
            .O(N__8603),
            .I(N__8600));
    LocalMux I__1862 (
            .O(N__8600),
            .I(N__8597));
    IoSpan4Mux I__1861 (
            .O(N__8597),
            .I(N__8593));
    InMux I__1860 (
            .O(N__8596),
            .I(N__8590));
    Span4Mux_s2_h I__1859 (
            .O(N__8593),
            .I(N__8587));
    LocalMux I__1858 (
            .O(N__8590),
            .I(N__8584));
    Sp12to4 I__1857 (
            .O(N__8587),
            .I(N__8581));
    Sp12to4 I__1856 (
            .O(N__8584),
            .I(N__8578));
    Span12Mux_h I__1855 (
            .O(N__8581),
            .I(N__8575));
    Span12Mux_s9_v I__1854 (
            .O(N__8578),
            .I(N__8572));
    Span12Mux_h I__1853 (
            .O(N__8575),
            .I(N__8569));
    Span12Mux_h I__1852 (
            .O(N__8572),
            .I(N__8566));
    Odrv12 I__1851 (
            .O(N__8569),
            .I(D_LM_040_in_7));
    Odrv12 I__1850 (
            .O(N__8566),
            .I(D_LM_040_in_7));
    IoInMux I__1849 (
            .O(N__8561),
            .I(N__8558));
    LocalMux I__1848 (
            .O(N__8558),
            .I(N__8555));
    Span4Mux_s2_v I__1847 (
            .O(N__8555),
            .I(N__8552));
    Span4Mux_v I__1846 (
            .O(N__8552),
            .I(N__8549));
    Sp12to4 I__1845 (
            .O(N__8549),
            .I(N__8546));
    Span12Mux_s11_h I__1844 (
            .O(N__8546),
            .I(N__8543));
    Odrv12 I__1843 (
            .O(N__8543),
            .I(un1_D_UU_040_7));
    InMux I__1842 (
            .O(N__8540),
            .I(N__8537));
    LocalMux I__1841 (
            .O(N__8537),
            .I(N__8534));
    Span4Mux_v I__1840 (
            .O(N__8534),
            .I(N__8531));
    Odrv4 I__1839 (
            .O(N__8531),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ));
    InMux I__1838 (
            .O(N__8528),
            .I(N__8524));
    InMux I__1837 (
            .O(N__8527),
            .I(N__8521));
    LocalMux I__1836 (
            .O(N__8524),
            .I(N__8518));
    LocalMux I__1835 (
            .O(N__8521),
            .I(N__8514));
    Span4Mux_h I__1834 (
            .O(N__8518),
            .I(N__8511));
    InMux I__1833 (
            .O(N__8517),
            .I(N__8508));
    Sp12to4 I__1832 (
            .O(N__8514),
            .I(N__8505));
    Span4Mux_v I__1831 (
            .O(N__8511),
            .I(N__8500));
    LocalMux I__1830 (
            .O(N__8508),
            .I(N__8500));
    Span12Mux_v I__1829 (
            .O(N__8505),
            .I(N__8497));
    Span4Mux_v I__1828 (
            .O(N__8500),
            .I(N__8494));
    Span12Mux_h I__1827 (
            .O(N__8497),
            .I(N__8491));
    Sp12to4 I__1826 (
            .O(N__8494),
            .I(N__8488));
    Span12Mux_v I__1825 (
            .O(N__8491),
            .I(N__8483));
    Span12Mux_h I__1824 (
            .O(N__8488),
            .I(N__8483));
    Odrv12 I__1823 (
            .O(N__8483),
            .I(D_UM_AMIGA_in_4));
    IoInMux I__1822 (
            .O(N__8480),
            .I(N__8477));
    LocalMux I__1821 (
            .O(N__8477),
            .I(N__8474));
    IoSpan4Mux I__1820 (
            .O(N__8474),
            .I(N__8471));
    IoSpan4Mux I__1819 (
            .O(N__8471),
            .I(N__8468));
    IoSpan4Mux I__1818 (
            .O(N__8468),
            .I(N__8465));
    Span4Mux_s2_v I__1817 (
            .O(N__8465),
            .I(N__8462));
    Span4Mux_v I__1816 (
            .O(N__8462),
            .I(N__8459));
    Odrv4 I__1815 (
            .O(N__8459),
            .I(un1_D_UM_AMIGA_4));
    InMux I__1814 (
            .O(N__8456),
            .I(N__8453));
    LocalMux I__1813 (
            .O(N__8453),
            .I(N__8449));
    InMux I__1812 (
            .O(N__8452),
            .I(N__8445));
    Span4Mux_v I__1811 (
            .O(N__8449),
            .I(N__8442));
    InMux I__1810 (
            .O(N__8448),
            .I(N__8439));
    LocalMux I__1809 (
            .O(N__8445),
            .I(N__8436));
    Span4Mux_v I__1808 (
            .O(N__8442),
            .I(N__8431));
    LocalMux I__1807 (
            .O(N__8439),
            .I(N__8431));
    Span4Mux_v I__1806 (
            .O(N__8436),
            .I(N__8428));
    Span4Mux_v I__1805 (
            .O(N__8431),
            .I(N__8425));
    Span4Mux_h I__1804 (
            .O(N__8428),
            .I(N__8422));
    Sp12to4 I__1803 (
            .O(N__8425),
            .I(N__8419));
    Sp12to4 I__1802 (
            .O(N__8422),
            .I(N__8416));
    Span12Mux_h I__1801 (
            .O(N__8419),
            .I(N__8413));
    Odrv12 I__1800 (
            .O(N__8416),
            .I(D_UU_AMIGA_in_4));
    Odrv12 I__1799 (
            .O(N__8413),
            .I(D_UU_AMIGA_in_4));
    InMux I__1798 (
            .O(N__8408),
            .I(N__8405));
    LocalMux I__1797 (
            .O(N__8405),
            .I(N__8402));
    Odrv12 I__1796 (
            .O(N__8402),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ));
    IoInMux I__1795 (
            .O(N__8399),
            .I(N__8396));
    LocalMux I__1794 (
            .O(N__8396),
            .I(N__8393));
    Span4Mux_s3_v I__1793 (
            .O(N__8393),
            .I(N__8390));
    Span4Mux_h I__1792 (
            .O(N__8390),
            .I(N__8387));
    Span4Mux_h I__1791 (
            .O(N__8387),
            .I(N__8384));
    Odrv4 I__1790 (
            .O(N__8384),
            .I(un1_D_UU_AMIGA_4));
    InMux I__1789 (
            .O(N__8381),
            .I(N__8378));
    LocalMux I__1788 (
            .O(N__8378),
            .I(N__8375));
    Odrv12 I__1787 (
            .O(N__8375),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ));
    InMux I__1786 (
            .O(N__8372),
            .I(N__8368));
    InMux I__1785 (
            .O(N__8371),
            .I(N__8365));
    LocalMux I__1784 (
            .O(N__8368),
            .I(N__8362));
    LocalMux I__1783 (
            .O(N__8365),
            .I(N__8359));
    Span4Mux_h I__1782 (
            .O(N__8362),
            .I(N__8356));
    Span4Mux_h I__1781 (
            .O(N__8359),
            .I(N__8353));
    Sp12to4 I__1780 (
            .O(N__8356),
            .I(N__8349));
    Span4Mux_v I__1779 (
            .O(N__8353),
            .I(N__8346));
    InMux I__1778 (
            .O(N__8352),
            .I(N__8343));
    Span12Mux_v I__1777 (
            .O(N__8349),
            .I(N__8340));
    Span4Mux_h I__1776 (
            .O(N__8346),
            .I(N__8337));
    LocalMux I__1775 (
            .O(N__8343),
            .I(N__8334));
    Span12Mux_h I__1774 (
            .O(N__8340),
            .I(N__8331));
    Sp12to4 I__1773 (
            .O(N__8337),
            .I(N__8326));
    Span12Mux_v I__1772 (
            .O(N__8334),
            .I(N__8326));
    Odrv12 I__1771 (
            .O(N__8331),
            .I(D_UU_AMIGA_in_5));
    Odrv12 I__1770 (
            .O(N__8326),
            .I(D_UU_AMIGA_in_5));
    IoInMux I__1769 (
            .O(N__8321),
            .I(N__8318));
    LocalMux I__1768 (
            .O(N__8318),
            .I(N__8315));
    Span4Mux_s3_v I__1767 (
            .O(N__8315),
            .I(N__8312));
    Span4Mux_h I__1766 (
            .O(N__8312),
            .I(N__8309));
    Span4Mux_h I__1765 (
            .O(N__8309),
            .I(N__8306));
    Span4Mux_h I__1764 (
            .O(N__8306),
            .I(N__8303));
    Odrv4 I__1763 (
            .O(N__8303),
            .I(un1_D_UU_AMIGA_5));
    IoInMux I__1762 (
            .O(N__8300),
            .I(N__8297));
    LocalMux I__1761 (
            .O(N__8297),
            .I(N__8294));
    IoSpan4Mux I__1760 (
            .O(N__8294),
            .I(N__8291));
    Span4Mux_s3_h I__1759 (
            .O(N__8291),
            .I(N__8288));
    Sp12to4 I__1758 (
            .O(N__8288),
            .I(N__8285));
    Span12Mux_h I__1757 (
            .O(N__8285),
            .I(N__8282));
    Odrv12 I__1756 (
            .O(N__8282),
            .I(N_224_i));
    InMux I__1755 (
            .O(N__8279),
            .I(N__8276));
    LocalMux I__1754 (
            .O(N__8276),
            .I(N__8273));
    Span4Mux_v I__1753 (
            .O(N__8273),
            .I(N__8268));
    InMux I__1752 (
            .O(N__8272),
            .I(N__8265));
    InMux I__1751 (
            .O(N__8271),
            .I(N__8262));
    Span4Mux_v I__1750 (
            .O(N__8268),
            .I(N__8255));
    LocalMux I__1749 (
            .O(N__8265),
            .I(N__8255));
    LocalMux I__1748 (
            .O(N__8262),
            .I(N__8255));
    Span4Mux_v I__1747 (
            .O(N__8255),
            .I(N__8252));
    Sp12to4 I__1746 (
            .O(N__8252),
            .I(N__8249));
    Span12Mux_h I__1745 (
            .O(N__8249),
            .I(N__8246));
    Odrv12 I__1744 (
            .O(N__8246),
            .I(D_UM_AMIGA_in_2));
    InMux I__1743 (
            .O(N__8243),
            .I(N__8240));
    LocalMux I__1742 (
            .O(N__8240),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ));
    CEMux I__1741 (
            .O(N__8237),
            .I(N__8231));
    CEMux I__1740 (
            .O(N__8236),
            .I(N__8228));
    CEMux I__1739 (
            .O(N__8235),
            .I(N__8225));
    CEMux I__1738 (
            .O(N__8234),
            .I(N__8222));
    LocalMux I__1737 (
            .O(N__8231),
            .I(\U111_CYCLE_SM.N_40_i_0 ));
    LocalMux I__1736 (
            .O(N__8228),
            .I(\U111_CYCLE_SM.N_40_i_0 ));
    LocalMux I__1735 (
            .O(N__8225),
            .I(\U111_CYCLE_SM.N_40_i_0 ));
    LocalMux I__1734 (
            .O(N__8222),
            .I(\U111_CYCLE_SM.N_40_i_0 ));
    SRMux I__1733 (
            .O(N__8213),
            .I(N__8208));
    SRMux I__1732 (
            .O(N__8212),
            .I(N__8205));
    SRMux I__1731 (
            .O(N__8211),
            .I(N__8202));
    LocalMux I__1730 (
            .O(N__8208),
            .I(N__8198));
    LocalMux I__1729 (
            .O(N__8205),
            .I(N__8195));
    LocalMux I__1728 (
            .O(N__8202),
            .I(N__8192));
    SRMux I__1727 (
            .O(N__8201),
            .I(N__8189));
    Span4Mux_v I__1726 (
            .O(N__8198),
            .I(N__8184));
    Span4Mux_v I__1725 (
            .O(N__8195),
            .I(N__8184));
    Span4Mux_h I__1724 (
            .O(N__8192),
            .I(N__8179));
    LocalMux I__1723 (
            .O(N__8189),
            .I(N__8179));
    Span4Mux_h I__1722 (
            .O(N__8184),
            .I(N__8176));
    Span4Mux_v I__1721 (
            .O(N__8179),
            .I(N__8173));
    Odrv4 I__1720 (
            .O(N__8176),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81 ));
    Odrv4 I__1719 (
            .O(N__8173),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81 ));
    InMux I__1718 (
            .O(N__8168),
            .I(N__8165));
    LocalMux I__1717 (
            .O(N__8165),
            .I(N__8160));
    InMux I__1716 (
            .O(N__8164),
            .I(N__8157));
    InMux I__1715 (
            .O(N__8163),
            .I(N__8154));
    Span4Mux_v I__1714 (
            .O(N__8160),
            .I(N__8151));
    LocalMux I__1713 (
            .O(N__8157),
            .I(N__8146));
    LocalMux I__1712 (
            .O(N__8154),
            .I(N__8146));
    Sp12to4 I__1711 (
            .O(N__8151),
            .I(N__8143));
    Sp12to4 I__1710 (
            .O(N__8146),
            .I(N__8140));
    Span12Mux_h I__1709 (
            .O(N__8143),
            .I(N__8137));
    Span12Mux_v I__1708 (
            .O(N__8140),
            .I(N__8134));
    Span12Mux_v I__1707 (
            .O(N__8137),
            .I(N__8131));
    Span12Mux_h I__1706 (
            .O(N__8134),
            .I(N__8128));
    Odrv12 I__1705 (
            .O(N__8131),
            .I(D_UU_AMIGA_in_0));
    Odrv12 I__1704 (
            .O(N__8128),
            .I(D_UU_AMIGA_in_0));
    InMux I__1703 (
            .O(N__8123),
            .I(N__8120));
    LocalMux I__1702 (
            .O(N__8120),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ));
    IoInMux I__1701 (
            .O(N__8117),
            .I(N__8114));
    LocalMux I__1700 (
            .O(N__8114),
            .I(N__8111));
    Span4Mux_s2_v I__1699 (
            .O(N__8111),
            .I(N__8108));
    Span4Mux_h I__1698 (
            .O(N__8108),
            .I(N__8105));
    Sp12to4 I__1697 (
            .O(N__8105),
            .I(N__8102));
    Span12Mux_s11_v I__1696 (
            .O(N__8102),
            .I(N__8099));
    Odrv12 I__1695 (
            .O(N__8099),
            .I(un1_D_UU_AMIGA_0));
    IoInMux I__1694 (
            .O(N__8096),
            .I(N__8093));
    LocalMux I__1693 (
            .O(N__8093),
            .I(N__8090));
    Span4Mux_s3_h I__1692 (
            .O(N__8090),
            .I(N__8087));
    Span4Mux_h I__1691 (
            .O(N__8087),
            .I(N__8084));
    Sp12to4 I__1690 (
            .O(N__8084),
            .I(N__8081));
    Span12Mux_s8_v I__1689 (
            .O(N__8081),
            .I(N__8078));
    Odrv12 I__1688 (
            .O(N__8078),
            .I(N_206_i));
    InMux I__1687 (
            .O(N__8075),
            .I(N__8072));
    LocalMux I__1686 (
            .O(N__8072),
            .I(N__8069));
    Span4Mux_v I__1685 (
            .O(N__8069),
            .I(N__8065));
    CascadeMux I__1684 (
            .O(N__8068),
            .I(N__8062));
    Span4Mux_v I__1683 (
            .O(N__8065),
            .I(N__8059));
    InMux I__1682 (
            .O(N__8062),
            .I(N__8056));
    Odrv4 I__1681 (
            .O(N__8059),
            .I(\U111_CYCLE_SM.TA_DISZ0 ));
    LocalMux I__1680 (
            .O(N__8056),
            .I(\U111_CYCLE_SM.TA_DISZ0 ));
    InMux I__1679 (
            .O(N__8051),
            .I(N__8046));
    CascadeMux I__1678 (
            .O(N__8050),
            .I(N__8043));
    InMux I__1677 (
            .O(N__8049),
            .I(N__8040));
    LocalMux I__1676 (
            .O(N__8046),
            .I(N__8037));
    InMux I__1675 (
            .O(N__8043),
            .I(N__8034));
    LocalMux I__1674 (
            .O(N__8040),
            .I(N__8030));
    Span4Mux_v I__1673 (
            .O(N__8037),
            .I(N__8025));
    LocalMux I__1672 (
            .O(N__8034),
            .I(N__8025));
    InMux I__1671 (
            .O(N__8033),
            .I(N__8022));
    Span4Mux_v I__1670 (
            .O(N__8030),
            .I(N__8019));
    Span4Mux_v I__1669 (
            .O(N__8025),
            .I(N__8016));
    LocalMux I__1668 (
            .O(N__8022),
            .I(N__8012));
    Sp12to4 I__1667 (
            .O(N__8019),
            .I(N__8009));
    Sp12to4 I__1666 (
            .O(N__8016),
            .I(N__8006));
    InMux I__1665 (
            .O(N__8015),
            .I(N__8003));
    Span12Mux_v I__1664 (
            .O(N__8012),
            .I(N__7996));
    Span12Mux_h I__1663 (
            .O(N__8009),
            .I(N__7996));
    Span12Mux_h I__1662 (
            .O(N__8006),
            .I(N__7996));
    LocalMux I__1661 (
            .O(N__8003),
            .I(N__7993));
    Span12Mux_v I__1660 (
            .O(N__7996),
            .I(N__7990));
    Span4Mux_v I__1659 (
            .O(N__7993),
            .I(N__7987));
    Odrv12 I__1658 (
            .O(N__7990),
            .I(LBENn_c));
    Odrv4 I__1657 (
            .O(N__7987),
            .I(LBENn_c));
    IoInMux I__1656 (
            .O(N__7982),
            .I(N__7979));
    LocalMux I__1655 (
            .O(N__7979),
            .I(N__7976));
    Span4Mux_s3_v I__1654 (
            .O(N__7976),
            .I(N__7973));
    Span4Mux_v I__1653 (
            .O(N__7973),
            .I(N__7970));
    Odrv4 I__1652 (
            .O(N__7970),
            .I(TAn_1_i));
    IoInMux I__1651 (
            .O(N__7967),
            .I(N__7964));
    LocalMux I__1650 (
            .O(N__7964),
            .I(N__7961));
    Span4Mux_s1_h I__1649 (
            .O(N__7961),
            .I(N__7958));
    Sp12to4 I__1648 (
            .O(N__7958),
            .I(N__7954));
    InMux I__1647 (
            .O(N__7957),
            .I(N__7951));
    Span12Mux_v I__1646 (
            .O(N__7954),
            .I(N__7948));
    LocalMux I__1645 (
            .O(N__7951),
            .I(N__7945));
    Span12Mux_h I__1644 (
            .O(N__7948),
            .I(N__7942));
    Span12Mux_h I__1643 (
            .O(N__7945),
            .I(N__7939));
    Span12Mux_h I__1642 (
            .O(N__7942),
            .I(N__7934));
    Span12Mux_v I__1641 (
            .O(N__7939),
            .I(N__7934));
    Odrv12 I__1640 (
            .O(N__7934),
            .I(D_LM_040_in_4));
    InMux I__1639 (
            .O(N__7931),
            .I(N__7928));
    LocalMux I__1638 (
            .O(N__7928),
            .I(N__7925));
    Span4Mux_v I__1637 (
            .O(N__7925),
            .I(N__7922));
    Sp12to4 I__1636 (
            .O(N__7922),
            .I(N__7919));
    Span12Mux_h I__1635 (
            .O(N__7919),
            .I(N__7916));
    Odrv12 I__1634 (
            .O(N__7916),
            .I(D_UU_040_in_4));
    IoInMux I__1633 (
            .O(N__7913),
            .I(N__7910));
    LocalMux I__1632 (
            .O(N__7910),
            .I(N__7907));
    Span4Mux_s2_v I__1631 (
            .O(N__7907),
            .I(N__7904));
    Span4Mux_v I__1630 (
            .O(N__7904),
            .I(N__7901));
    Sp12to4 I__1629 (
            .O(N__7901),
            .I(N__7898));
    Odrv12 I__1628 (
            .O(N__7898),
            .I(un1_D_UU_040_4));
    InMux I__1627 (
            .O(N__7895),
            .I(N__7892));
    LocalMux I__1626 (
            .O(N__7892),
            .I(N__7889));
    Span4Mux_v I__1625 (
            .O(N__7889),
            .I(N__7886));
    Sp12to4 I__1624 (
            .O(N__7886),
            .I(N__7883));
    Span12Mux_h I__1623 (
            .O(N__7883),
            .I(N__7880));
    Odrv12 I__1622 (
            .O(N__7880),
            .I(D_LL_AMIGA_in_1));
    IoInMux I__1621 (
            .O(N__7877),
            .I(N__7874));
    LocalMux I__1620 (
            .O(N__7874),
            .I(N__7871));
    Span4Mux_s3_h I__1619 (
            .O(N__7871),
            .I(N__7868));
    Span4Mux_v I__1618 (
            .O(N__7868),
            .I(N__7865));
    Sp12to4 I__1617 (
            .O(N__7865),
            .I(N__7862));
    Span12Mux_h I__1616 (
            .O(N__7862),
            .I(N__7859));
    Odrv12 I__1615 (
            .O(N__7859),
            .I(un2_D_LL_AMIGA_1));
    InMux I__1614 (
            .O(N__7856),
            .I(N__7853));
    LocalMux I__1613 (
            .O(N__7853),
            .I(N__7850));
    Span4Mux_v I__1612 (
            .O(N__7850),
            .I(N__7847));
    Sp12to4 I__1611 (
            .O(N__7847),
            .I(N__7844));
    Span12Mux_h I__1610 (
            .O(N__7844),
            .I(N__7841));
    Odrv12 I__1609 (
            .O(N__7841),
            .I(D_LL_AMIGA_in_4));
    IoInMux I__1608 (
            .O(N__7838),
            .I(N__7835));
    LocalMux I__1607 (
            .O(N__7835),
            .I(N__7832));
    IoSpan4Mux I__1606 (
            .O(N__7832),
            .I(N__7829));
    Span4Mux_s2_h I__1605 (
            .O(N__7829),
            .I(N__7826));
    Sp12to4 I__1604 (
            .O(N__7826),
            .I(N__7823));
    Span12Mux_h I__1603 (
            .O(N__7823),
            .I(N__7820));
    Odrv12 I__1602 (
            .O(N__7820),
            .I(un2_D_LL_AMIGA_4));
    IoInMux I__1601 (
            .O(N__7817),
            .I(N__7814));
    LocalMux I__1600 (
            .O(N__7814),
            .I(N__7810));
    InMux I__1599 (
            .O(N__7813),
            .I(N__7807));
    IoSpan4Mux I__1598 (
            .O(N__7810),
            .I(N__7804));
    LocalMux I__1597 (
            .O(N__7807),
            .I(N__7801));
    Span4Mux_s2_h I__1596 (
            .O(N__7804),
            .I(N__7798));
    Span4Mux_v I__1595 (
            .O(N__7801),
            .I(N__7795));
    Sp12to4 I__1594 (
            .O(N__7798),
            .I(N__7792));
    Sp12to4 I__1593 (
            .O(N__7795),
            .I(N__7789));
    Span12Mux_h I__1592 (
            .O(N__7792),
            .I(N__7786));
    Span12Mux_v I__1591 (
            .O(N__7789),
            .I(N__7783));
    Span12Mux_h I__1590 (
            .O(N__7786),
            .I(N__7780));
    Span12Mux_h I__1589 (
            .O(N__7783),
            .I(N__7777));
    Odrv12 I__1588 (
            .O(N__7780),
            .I(D_LL_040_in_0));
    Odrv12 I__1587 (
            .O(N__7777),
            .I(D_LL_040_in_0));
    InMux I__1586 (
            .O(N__7772),
            .I(N__7769));
    LocalMux I__1585 (
            .O(N__7769),
            .I(N__7766));
    Span12Mux_h I__1584 (
            .O(N__7766),
            .I(N__7763));
    Odrv12 I__1583 (
            .O(N__7763),
            .I(D_UM_040_in_0));
    IoInMux I__1582 (
            .O(N__7760),
            .I(N__7757));
    LocalMux I__1581 (
            .O(N__7757),
            .I(N__7754));
    IoSpan4Mux I__1580 (
            .O(N__7754),
            .I(N__7751));
    Span4Mux_s2_h I__1579 (
            .O(N__7751),
            .I(N__7748));
    Span4Mux_h I__1578 (
            .O(N__7748),
            .I(N__7745));
    Span4Mux_h I__1577 (
            .O(N__7745),
            .I(N__7742));
    Span4Mux_h I__1576 (
            .O(N__7742),
            .I(N__7739));
    Odrv4 I__1575 (
            .O(N__7739),
            .I(un1_D_UM_040_0));
    IoInMux I__1574 (
            .O(N__7736),
            .I(N__7733));
    LocalMux I__1573 (
            .O(N__7733),
            .I(N__7730));
    IoSpan4Mux I__1572 (
            .O(N__7730),
            .I(N__7727));
    Span4Mux_s3_h I__1571 (
            .O(N__7727),
            .I(N__7724));
    Span4Mux_h I__1570 (
            .O(N__7724),
            .I(N__7721));
    Span4Mux_h I__1569 (
            .O(N__7721),
            .I(N__7718));
    Odrv4 I__1568 (
            .O(N__7718),
            .I(un1_D_UM_AMIGA_2));
    InMux I__1567 (
            .O(N__7715),
            .I(N__7712));
    LocalMux I__1566 (
            .O(N__7712),
            .I(N__7709));
    Glb2LocalMux I__1565 (
            .O(N__7709),
            .I(N__7706));
    GlobalMux I__1564 (
            .O(N__7706),
            .I(CLK80));
    IoInMux I__1563 (
            .O(N__7703),
            .I(N__7700));
    LocalMux I__1562 (
            .O(N__7700),
            .I(N__7696));
    IoInMux I__1561 (
            .O(N__7699),
            .I(N__7693));
    Span4Mux_s0_v I__1560 (
            .O(N__7696),
            .I(N__7690));
    LocalMux I__1559 (
            .O(N__7693),
            .I(N__7687));
    Sp12to4 I__1558 (
            .O(N__7690),
            .I(N__7684));
    Span4Mux_s3_h I__1557 (
            .O(N__7687),
            .I(N__7681));
    Span12Mux_h I__1556 (
            .O(N__7684),
            .I(N__7678));
    Span4Mux_v I__1555 (
            .O(N__7681),
            .I(N__7675));
    Span12Mux_v I__1554 (
            .O(N__7678),
            .I(N__7672));
    Sp12to4 I__1553 (
            .O(N__7675),
            .I(N__7669));
    Odrv12 I__1552 (
            .O(N__7672),
            .I(GB_BUFFER_CLK80_THRU_CO));
    Odrv12 I__1551 (
            .O(N__7669),
            .I(GB_BUFFER_CLK80_THRU_CO));
    InMux I__1550 (
            .O(N__7664),
            .I(N__7661));
    LocalMux I__1549 (
            .O(N__7661),
            .I(N__7658));
    Odrv4 I__1548 (
            .O(N__7658),
            .I(READ_CYCLE_ACTIVE_rep5_i_ess));
    IoInMux I__1547 (
            .O(N__7655),
            .I(N__7652));
    LocalMux I__1546 (
            .O(N__7652),
            .I(N__7649));
    IoSpan4Mux I__1545 (
            .O(N__7649),
            .I(N__7646));
    Span4Mux_s0_v I__1544 (
            .O(N__7646),
            .I(N__7643));
    Sp12to4 I__1543 (
            .O(N__7643),
            .I(N__7640));
    Span12Mux_s11_v I__1542 (
            .O(N__7640),
            .I(N__7637));
    Odrv12 I__1541 (
            .O(N__7637),
            .I(N_210_i));
    InMux I__1540 (
            .O(N__7634),
            .I(N__7631));
    LocalMux I__1539 (
            .O(N__7631),
            .I(N__7628));
    Span4Mux_v I__1538 (
            .O(N__7628),
            .I(N__7625));
    Sp12to4 I__1537 (
            .O(N__7625),
            .I(N__7622));
    Span12Mux_h I__1536 (
            .O(N__7622),
            .I(N__7619));
    Span12Mux_v I__1535 (
            .O(N__7619),
            .I(N__7616));
    Odrv12 I__1534 (
            .O(N__7616),
            .I(D_UM_040_in_1));
    IoInMux I__1533 (
            .O(N__7613),
            .I(N__7610));
    LocalMux I__1532 (
            .O(N__7610),
            .I(N__7607));
    Span4Mux_s3_h I__1531 (
            .O(N__7607),
            .I(N__7603));
    InMux I__1530 (
            .O(N__7606),
            .I(N__7600));
    Sp12to4 I__1529 (
            .O(N__7603),
            .I(N__7597));
    LocalMux I__1528 (
            .O(N__7600),
            .I(N__7594));
    Span12Mux_v I__1527 (
            .O(N__7597),
            .I(N__7591));
    Span12Mux_v I__1526 (
            .O(N__7594),
            .I(N__7588));
    Span12Mux_h I__1525 (
            .O(N__7591),
            .I(N__7583));
    Span12Mux_v I__1524 (
            .O(N__7588),
            .I(N__7583));
    Span12Mux_h I__1523 (
            .O(N__7583),
            .I(N__7580));
    Odrv12 I__1522 (
            .O(N__7580),
            .I(D_LL_040_in_1));
    IoInMux I__1521 (
            .O(N__7577),
            .I(N__7574));
    LocalMux I__1520 (
            .O(N__7574),
            .I(N__7571));
    Span4Mux_s3_h I__1519 (
            .O(N__7571),
            .I(N__7568));
    Span4Mux_h I__1518 (
            .O(N__7568),
            .I(N__7565));
    Span4Mux_h I__1517 (
            .O(N__7565),
            .I(N__7562));
    Span4Mux_h I__1516 (
            .O(N__7562),
            .I(N__7559));
    Odrv4 I__1515 (
            .O(N__7559),
            .I(un1_D_UM_040_1));
    InMux I__1514 (
            .O(N__7556),
            .I(N__7553));
    LocalMux I__1513 (
            .O(N__7553),
            .I(N__7550));
    Odrv4 I__1512 (
            .O(N__7550),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ));
    InMux I__1511 (
            .O(N__7547),
            .I(N__7542));
    InMux I__1510 (
            .O(N__7546),
            .I(N__7539));
    InMux I__1509 (
            .O(N__7545),
            .I(N__7536));
    LocalMux I__1508 (
            .O(N__7542),
            .I(N__7531));
    LocalMux I__1507 (
            .O(N__7539),
            .I(N__7531));
    LocalMux I__1506 (
            .O(N__7536),
            .I(N__7528));
    Span12Mux_v I__1505 (
            .O(N__7531),
            .I(N__7525));
    Span12Mux_v I__1504 (
            .O(N__7528),
            .I(N__7522));
    Span12Mux_h I__1503 (
            .O(N__7525),
            .I(N__7519));
    Odrv12 I__1502 (
            .O(N__7522),
            .I(D_UU_AMIGA_in_1));
    Odrv12 I__1501 (
            .O(N__7519),
            .I(D_UU_AMIGA_in_1));
    IoInMux I__1500 (
            .O(N__7514),
            .I(N__7511));
    LocalMux I__1499 (
            .O(N__7511),
            .I(N__7508));
    IoSpan4Mux I__1498 (
            .O(N__7508),
            .I(N__7505));
    Span4Mux_s3_h I__1497 (
            .O(N__7505),
            .I(N__7502));
    Span4Mux_h I__1496 (
            .O(N__7502),
            .I(N__7499));
    Sp12to4 I__1495 (
            .O(N__7499),
            .I(N__7496));
    Span12Mux_h I__1494 (
            .O(N__7496),
            .I(N__7493));
    Odrv12 I__1493 (
            .O(N__7493),
            .I(un1_D_UU_AMIGA_1));
    InMux I__1492 (
            .O(N__7490),
            .I(N__7487));
    LocalMux I__1491 (
            .O(N__7487),
            .I(N__7482));
    InMux I__1490 (
            .O(N__7486),
            .I(N__7479));
    InMux I__1489 (
            .O(N__7485),
            .I(N__7476));
    Span4Mux_v I__1488 (
            .O(N__7482),
            .I(N__7471));
    LocalMux I__1487 (
            .O(N__7479),
            .I(N__7471));
    LocalMux I__1486 (
            .O(N__7476),
            .I(N__7468));
    Span4Mux_h I__1485 (
            .O(N__7471),
            .I(N__7465));
    Span12Mux_v I__1484 (
            .O(N__7468),
            .I(N__7462));
    Span4Mux_v I__1483 (
            .O(N__7465),
            .I(N__7459));
    Span12Mux_h I__1482 (
            .O(N__7462),
            .I(N__7456));
    Span4Mux_h I__1481 (
            .O(N__7459),
            .I(N__7453));
    Span12Mux_v I__1480 (
            .O(N__7456),
            .I(N__7450));
    Sp12to4 I__1479 (
            .O(N__7453),
            .I(N__7447));
    Odrv12 I__1478 (
            .O(N__7450),
            .I(D_UM_AMIGA_in_3));
    Odrv12 I__1477 (
            .O(N__7447),
            .I(D_UM_AMIGA_in_3));
    InMux I__1476 (
            .O(N__7442),
            .I(N__7439));
    LocalMux I__1475 (
            .O(N__7439),
            .I(N__7436));
    Odrv4 I__1474 (
            .O(N__7436),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ));
    IoInMux I__1473 (
            .O(N__7433),
            .I(N__7430));
    LocalMux I__1472 (
            .O(N__7430),
            .I(N__7427));
    Span4Mux_s2_h I__1471 (
            .O(N__7427),
            .I(N__7424));
    Span4Mux_v I__1470 (
            .O(N__7424),
            .I(N__7421));
    Span4Mux_v I__1469 (
            .O(N__7421),
            .I(N__7418));
    Sp12to4 I__1468 (
            .O(N__7418),
            .I(N__7415));
    Span12Mux_h I__1467 (
            .O(N__7415),
            .I(N__7412));
    Odrv12 I__1466 (
            .O(N__7412),
            .I(un1_D_UM_AMIGA_3));
    InMux I__1465 (
            .O(N__7409),
            .I(N__7405));
    InMux I__1464 (
            .O(N__7408),
            .I(N__7402));
    LocalMux I__1463 (
            .O(N__7405),
            .I(N__7398));
    LocalMux I__1462 (
            .O(N__7402),
            .I(N__7395));
    InMux I__1461 (
            .O(N__7401),
            .I(N__7392));
    Span4Mux_v I__1460 (
            .O(N__7398),
            .I(N__7389));
    Span4Mux_v I__1459 (
            .O(N__7395),
            .I(N__7384));
    LocalMux I__1458 (
            .O(N__7392),
            .I(N__7384));
    Span4Mux_h I__1457 (
            .O(N__7389),
            .I(N__7381));
    Sp12to4 I__1456 (
            .O(N__7384),
            .I(N__7378));
    Sp12to4 I__1455 (
            .O(N__7381),
            .I(N__7375));
    Span12Mux_v I__1454 (
            .O(N__7378),
            .I(N__7372));
    Span12Mux_v I__1453 (
            .O(N__7375),
            .I(N__7367));
    Span12Mux_h I__1452 (
            .O(N__7372),
            .I(N__7367));
    Odrv12 I__1451 (
            .O(N__7367),
            .I(D_UM_AMIGA_in_5));
    InMux I__1450 (
            .O(N__7364),
            .I(N__7361));
    LocalMux I__1449 (
            .O(N__7361),
            .I(N__7358));
    Span4Mux_v I__1448 (
            .O(N__7358),
            .I(N__7355));
    Odrv4 I__1447 (
            .O(N__7355),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ));
    IoInMux I__1446 (
            .O(N__7352),
            .I(N__7349));
    LocalMux I__1445 (
            .O(N__7349),
            .I(N__7346));
    Span4Mux_s2_v I__1444 (
            .O(N__7346),
            .I(N__7343));
    Span4Mux_h I__1443 (
            .O(N__7343),
            .I(N__7340));
    Span4Mux_h I__1442 (
            .O(N__7340),
            .I(N__7337));
    Sp12to4 I__1441 (
            .O(N__7337),
            .I(N__7334));
    Span12Mux_s8_v I__1440 (
            .O(N__7334),
            .I(N__7331));
    Odrv12 I__1439 (
            .O(N__7331),
            .I(un1_D_UM_AMIGA_5));
    InMux I__1438 (
            .O(N__7328),
            .I(N__7325));
    LocalMux I__1437 (
            .O(N__7325),
            .I(N__7322));
    Odrv12 I__1436 (
            .O(N__7322),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ));
    InMux I__1435 (
            .O(N__7319),
            .I(N__7314));
    InMux I__1434 (
            .O(N__7318),
            .I(N__7311));
    InMux I__1433 (
            .O(N__7317),
            .I(N__7308));
    LocalMux I__1432 (
            .O(N__7314),
            .I(N__7305));
    LocalMux I__1431 (
            .O(N__7311),
            .I(N__7302));
    LocalMux I__1430 (
            .O(N__7308),
            .I(N__7299));
    Span4Mux_v I__1429 (
            .O(N__7305),
            .I(N__7296));
    Span4Mux_v I__1428 (
            .O(N__7302),
            .I(N__7291));
    Span4Mux_v I__1427 (
            .O(N__7299),
            .I(N__7291));
    Sp12to4 I__1426 (
            .O(N__7296),
            .I(N__7286));
    Sp12to4 I__1425 (
            .O(N__7291),
            .I(N__7286));
    Span12Mux_h I__1424 (
            .O(N__7286),
            .I(N__7283));
    Odrv12 I__1423 (
            .O(N__7283),
            .I(D_UU_AMIGA_in_2));
    IoInMux I__1422 (
            .O(N__7280),
            .I(N__7277));
    LocalMux I__1421 (
            .O(N__7277),
            .I(N__7274));
    Span4Mux_s2_v I__1420 (
            .O(N__7274),
            .I(N__7271));
    Sp12to4 I__1419 (
            .O(N__7271),
            .I(N__7268));
    Span12Mux_h I__1418 (
            .O(N__7268),
            .I(N__7265));
    Odrv12 I__1417 (
            .O(N__7265),
            .I(un1_D_UU_AMIGA_2));
    InMux I__1416 (
            .O(N__7262),
            .I(N__7259));
    LocalMux I__1415 (
            .O(N__7259),
            .I(N__7256));
    Odrv4 I__1414 (
            .O(N__7256),
            .I(READ_CYCLE_ACTIVE_rep1_i_ess));
    CascadeMux I__1413 (
            .O(N__7253),
            .I(\U111_CYCLE_SM.N_55_cascade_ ));
    InMux I__1412 (
            .O(N__7250),
            .I(N__7247));
    LocalMux I__1411 (
            .O(N__7247),
            .I(N__7243));
    InMux I__1410 (
            .O(N__7246),
            .I(N__7240));
    Odrv4 I__1409 (
            .O(N__7243),
            .I(\U111_CYCLE_SM.N_73 ));
    LocalMux I__1408 (
            .O(N__7240),
            .I(\U111_CYCLE_SM.N_73 ));
    InMux I__1407 (
            .O(N__7235),
            .I(N__7229));
    InMux I__1406 (
            .O(N__7234),
            .I(N__7226));
    InMux I__1405 (
            .O(N__7233),
            .I(N__7223));
    InMux I__1404 (
            .O(N__7232),
            .I(N__7220));
    LocalMux I__1403 (
            .O(N__7229),
            .I(N__7217));
    LocalMux I__1402 (
            .O(N__7226),
            .I(N__7212));
    LocalMux I__1401 (
            .O(N__7223),
            .I(N__7212));
    LocalMux I__1400 (
            .O(N__7220),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    Odrv12 I__1399 (
            .O(N__7217),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    Odrv4 I__1398 (
            .O(N__7212),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    IoInMux I__1397 (
            .O(N__7205),
            .I(N__7202));
    LocalMux I__1396 (
            .O(N__7202),
            .I(N__7199));
    Span4Mux_s1_v I__1395 (
            .O(N__7199),
            .I(N__7194));
    CascadeMux I__1394 (
            .O(N__7198),
            .I(N__7190));
    CascadeMux I__1393 (
            .O(N__7197),
            .I(N__7185));
    Span4Mux_v I__1392 (
            .O(N__7194),
            .I(N__7181));
    InMux I__1391 (
            .O(N__7193),
            .I(N__7178));
    InMux I__1390 (
            .O(N__7190),
            .I(N__7171));
    InMux I__1389 (
            .O(N__7189),
            .I(N__7171));
    InMux I__1388 (
            .O(N__7188),
            .I(N__7171));
    InMux I__1387 (
            .O(N__7185),
            .I(N__7166));
    InMux I__1386 (
            .O(N__7184),
            .I(N__7166));
    Span4Mux_v I__1385 (
            .O(N__7181),
            .I(N__7163));
    LocalMux I__1384 (
            .O(N__7178),
            .I(N__7156));
    LocalMux I__1383 (
            .O(N__7171),
            .I(N__7156));
    LocalMux I__1382 (
            .O(N__7166),
            .I(N__7156));
    Span4Mux_v I__1381 (
            .O(N__7163),
            .I(N__7150));
    Span4Mux_v I__1380 (
            .O(N__7156),
            .I(N__7150));
    CascadeMux I__1379 (
            .O(N__7155),
            .I(N__7147));
    Sp12to4 I__1378 (
            .O(N__7150),
            .I(N__7143));
    InMux I__1377 (
            .O(N__7147),
            .I(N__7138));
    InMux I__1376 (
            .O(N__7146),
            .I(N__7138));
    Span12Mux_h I__1375 (
            .O(N__7143),
            .I(N__7133));
    LocalMux I__1374 (
            .O(N__7138),
            .I(N__7133));
    Span12Mux_v I__1373 (
            .O(N__7133),
            .I(N__7130));
    Odrv12 I__1372 (
            .O(N__7130),
            .I(TACKn_in));
    CascadeMux I__1371 (
            .O(N__7127),
            .I(N__7120));
    InMux I__1370 (
            .O(N__7126),
            .I(N__7117));
    InMux I__1369 (
            .O(N__7125),
            .I(N__7108));
    InMux I__1368 (
            .O(N__7124),
            .I(N__7108));
    InMux I__1367 (
            .O(N__7123),
            .I(N__7108));
    InMux I__1366 (
            .O(N__7120),
            .I(N__7108));
    LocalMux I__1365 (
            .O(N__7117),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ));
    LocalMux I__1364 (
            .O(N__7108),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ));
    CascadeMux I__1363 (
            .O(N__7103),
            .I(\U111_CYCLE_SM.N_57_cascade_ ));
    InMux I__1362 (
            .O(N__7100),
            .I(N__7097));
    LocalMux I__1361 (
            .O(N__7097),
            .I(\U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_1_0 ));
    InMux I__1360 (
            .O(N__7094),
            .I(N__7091));
    LocalMux I__1359 (
            .O(N__7091),
            .I(N__7088));
    Span4Mux_h I__1358 (
            .O(N__7088),
            .I(N__7085));
    Span4Mux_h I__1357 (
            .O(N__7085),
            .I(N__7078));
    InMux I__1356 (
            .O(N__7084),
            .I(N__7075));
    InMux I__1355 (
            .O(N__7083),
            .I(N__7072));
    InMux I__1354 (
            .O(N__7082),
            .I(N__7069));
    InMux I__1353 (
            .O(N__7081),
            .I(N__7066));
    Span4Mux_h I__1352 (
            .O(N__7078),
            .I(N__7063));
    LocalMux I__1351 (
            .O(N__7075),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1350 (
            .O(N__7072),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1349 (
            .O(N__7069),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1348 (
            .O(N__7066),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    Odrv4 I__1347 (
            .O(N__7063),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    InMux I__1346 (
            .O(N__7052),
            .I(N__7048));
    InMux I__1345 (
            .O(N__7051),
            .I(N__7045));
    LocalMux I__1344 (
            .O(N__7048),
            .I(N__7040));
    LocalMux I__1343 (
            .O(N__7045),
            .I(N__7040));
    Odrv4 I__1342 (
            .O(N__7040),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_1 ));
    InMux I__1341 (
            .O(N__7037),
            .I(N__7031));
    InMux I__1340 (
            .O(N__7036),
            .I(N__7028));
    InMux I__1339 (
            .O(N__7035),
            .I(N__7025));
    InMux I__1338 (
            .O(N__7034),
            .I(N__7022));
    LocalMux I__1337 (
            .O(N__7031),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    LocalMux I__1336 (
            .O(N__7028),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    LocalMux I__1335 (
            .O(N__7025),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    LocalMux I__1334 (
            .O(N__7022),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    CascadeMux I__1333 (
            .O(N__7013),
            .I(N__7010));
    InMux I__1332 (
            .O(N__7010),
            .I(N__7007));
    LocalMux I__1331 (
            .O(N__7007),
            .I(N__7004));
    Sp12to4 I__1330 (
            .O(N__7004),
            .I(N__7000));
    IoInMux I__1329 (
            .O(N__7003),
            .I(N__6997));
    Span12Mux_h I__1328 (
            .O(N__7000),
            .I(N__6994));
    LocalMux I__1327 (
            .O(N__6997),
            .I(N__6991));
    Span12Mux_v I__1326 (
            .O(N__6994),
            .I(N__6988));
    IoSpan4Mux I__1325 (
            .O(N__6991),
            .I(N__6985));
    Odrv12 I__1324 (
            .O(N__6988),
            .I(TBIn_c));
    Odrv4 I__1323 (
            .O(N__6985),
            .I(TBIn_c));
    CascadeMux I__1322 (
            .O(N__6980),
            .I(N__6977));
    InMux I__1321 (
            .O(N__6977),
            .I(N__6972));
    InMux I__1320 (
            .O(N__6976),
            .I(N__6969));
    InMux I__1319 (
            .O(N__6975),
            .I(N__6966));
    LocalMux I__1318 (
            .O(N__6972),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ));
    LocalMux I__1317 (
            .O(N__6969),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ));
    LocalMux I__1316 (
            .O(N__6966),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ));
    InMux I__1315 (
            .O(N__6959),
            .I(N__6955));
    InMux I__1314 (
            .O(N__6958),
            .I(N__6952));
    LocalMux I__1313 (
            .O(N__6955),
            .I(\U111_CYCLE_SM.N_42 ));
    LocalMux I__1312 (
            .O(N__6952),
            .I(\U111_CYCLE_SM.N_42 ));
    CascadeMux I__1311 (
            .O(N__6947),
            .I(\U111_CYCLE_SM.N_46_cascade_ ));
    InMux I__1310 (
            .O(N__6944),
            .I(N__6936));
    InMux I__1309 (
            .O(N__6943),
            .I(N__6927));
    InMux I__1308 (
            .O(N__6942),
            .I(N__6927));
    InMux I__1307 (
            .O(N__6941),
            .I(N__6927));
    InMux I__1306 (
            .O(N__6940),
            .I(N__6927));
    InMux I__1305 (
            .O(N__6939),
            .I(N__6924));
    LocalMux I__1304 (
            .O(N__6936),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    LocalMux I__1303 (
            .O(N__6927),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    LocalMux I__1302 (
            .O(N__6924),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    CascadeMux I__1301 (
            .O(N__6917),
            .I(N__6914));
    InMux I__1300 (
            .O(N__6914),
            .I(N__6910));
    InMux I__1299 (
            .O(N__6913),
            .I(N__6907));
    LocalMux I__1298 (
            .O(N__6910),
            .I(N__6904));
    LocalMux I__1297 (
            .O(N__6907),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ));
    Odrv4 I__1296 (
            .O(N__6904),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ));
    InMux I__1295 (
            .O(N__6899),
            .I(N__6896));
    LocalMux I__1294 (
            .O(N__6896),
            .I(\U111_CYCLE_SM.N_39 ));
    InMux I__1293 (
            .O(N__6893),
            .I(N__6888));
    InMux I__1292 (
            .O(N__6892),
            .I(N__6883));
    InMux I__1291 (
            .O(N__6891),
            .I(N__6883));
    LocalMux I__1290 (
            .O(N__6888),
            .I(\U111_CYCLE_SM.N_40 ));
    LocalMux I__1289 (
            .O(N__6883),
            .I(\U111_CYCLE_SM.N_40 ));
    CascadeMux I__1288 (
            .O(N__6878),
            .I(\U111_CYCLE_SM.N_40_cascade_ ));
    InMux I__1287 (
            .O(N__6875),
            .I(N__6871));
    InMux I__1286 (
            .O(N__6874),
            .I(N__6867));
    LocalMux I__1285 (
            .O(N__6871),
            .I(N__6864));
    InMux I__1284 (
            .O(N__6870),
            .I(N__6861));
    LocalMux I__1283 (
            .O(N__6867),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    Odrv4 I__1282 (
            .O(N__6864),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    LocalMux I__1281 (
            .O(N__6861),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    CascadeMux I__1280 (
            .O(N__6854),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81_cascade_ ));
    IoInMux I__1279 (
            .O(N__6851),
            .I(N__6848));
    LocalMux I__1278 (
            .O(N__6848),
            .I(N__6844));
    CascadeMux I__1277 (
            .O(N__6847),
            .I(N__6838));
    Span4Mux_s1_v I__1276 (
            .O(N__6844),
            .I(N__6832));
    InMux I__1275 (
            .O(N__6843),
            .I(N__6825));
    InMux I__1274 (
            .O(N__6842),
            .I(N__6825));
    InMux I__1273 (
            .O(N__6841),
            .I(N__6825));
    InMux I__1272 (
            .O(N__6838),
            .I(N__6820));
    InMux I__1271 (
            .O(N__6837),
            .I(N__6820));
    InMux I__1270 (
            .O(N__6836),
            .I(N__6815));
    InMux I__1269 (
            .O(N__6835),
            .I(N__6815));
    Span4Mux_v I__1268 (
            .O(N__6832),
            .I(N__6812));
    LocalMux I__1267 (
            .O(N__6825),
            .I(N__6807));
    LocalMux I__1266 (
            .O(N__6820),
            .I(N__6807));
    LocalMux I__1265 (
            .O(N__6815),
            .I(N__6804));
    Sp12to4 I__1264 (
            .O(N__6812),
            .I(N__6801));
    Span4Mux_v I__1263 (
            .O(N__6807),
            .I(N__6798));
    Span4Mux_v I__1262 (
            .O(N__6804),
            .I(N__6795));
    Span12Mux_h I__1261 (
            .O(N__6801),
            .I(N__6792));
    Sp12to4 I__1260 (
            .O(N__6798),
            .I(N__6789));
    Span4Mux_h I__1259 (
            .O(N__6795),
            .I(N__6786));
    Span12Mux_v I__1258 (
            .O(N__6792),
            .I(N__6779));
    Span12Mux_h I__1257 (
            .O(N__6789),
            .I(N__6779));
    Sp12to4 I__1256 (
            .O(N__6786),
            .I(N__6779));
    Span12Mux_v I__1255 (
            .O(N__6779),
            .I(N__6776));
    Odrv12 I__1254 (
            .O(N__6776),
            .I(TEAn_c));
    InMux I__1253 (
            .O(N__6773),
            .I(N__6764));
    InMux I__1252 (
            .O(N__6772),
            .I(N__6764));
    InMux I__1251 (
            .O(N__6771),
            .I(N__6761));
    InMux I__1250 (
            .O(N__6770),
            .I(N__6756));
    InMux I__1249 (
            .O(N__6769),
            .I(N__6756));
    LocalMux I__1248 (
            .O(N__6764),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    LocalMux I__1247 (
            .O(N__6761),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    LocalMux I__1246 (
            .O(N__6756),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    InMux I__1245 (
            .O(N__6749),
            .I(N__6737));
    InMux I__1244 (
            .O(N__6748),
            .I(N__6737));
    InMux I__1243 (
            .O(N__6747),
            .I(N__6730));
    InMux I__1242 (
            .O(N__6746),
            .I(N__6730));
    InMux I__1241 (
            .O(N__6745),
            .I(N__6730));
    InMux I__1240 (
            .O(N__6744),
            .I(N__6725));
    InMux I__1239 (
            .O(N__6743),
            .I(N__6725));
    InMux I__1238 (
            .O(N__6742),
            .I(N__6722));
    LocalMux I__1237 (
            .O(N__6737),
            .I(N__6719));
    LocalMux I__1236 (
            .O(N__6730),
            .I(N__6716));
    LocalMux I__1235 (
            .O(N__6725),
            .I(N__6713));
    LocalMux I__1234 (
            .O(N__6722),
            .I(N__6710));
    Span4Mux_v I__1233 (
            .O(N__6719),
            .I(N__6704));
    Span4Mux_v I__1232 (
            .O(N__6716),
            .I(N__6704));
    Span4Mux_v I__1231 (
            .O(N__6713),
            .I(N__6701));
    Span4Mux_v I__1230 (
            .O(N__6710),
            .I(N__6698));
    InMux I__1229 (
            .O(N__6709),
            .I(N__6695));
    Sp12to4 I__1228 (
            .O(N__6704),
            .I(N__6688));
    Sp12to4 I__1227 (
            .O(N__6701),
            .I(N__6688));
    Sp12to4 I__1226 (
            .O(N__6698),
            .I(N__6688));
    LocalMux I__1225 (
            .O(N__6695),
            .I(N__6685));
    Span12Mux_h I__1224 (
            .O(N__6688),
            .I(N__6680));
    Span12Mux_s7_h I__1223 (
            .O(N__6685),
            .I(N__6680));
    Span12Mux_v I__1222 (
            .O(N__6680),
            .I(N__6677));
    Odrv12 I__1221 (
            .O(N__6677),
            .I(RESETn_c));
    InMux I__1220 (
            .O(N__6674),
            .I(N__6671));
    LocalMux I__1219 (
            .O(N__6671),
            .I(N__6668));
    Odrv4 I__1218 (
            .O(N__6668),
            .I(READ_CYCLE_ACTIVE_rep2_i_ess));
    IoInMux I__1217 (
            .O(N__6665),
            .I(N__6662));
    LocalMux I__1216 (
            .O(N__6662),
            .I(N__6659));
    Span12Mux_s8_v I__1215 (
            .O(N__6659),
            .I(N__6656));
    Span12Mux_h I__1214 (
            .O(N__6656),
            .I(N__6653));
    Odrv12 I__1213 (
            .O(N__6653),
            .I(N_207_i));
    InMux I__1212 (
            .O(N__6650),
            .I(N__6647));
    LocalMux I__1211 (
            .O(N__6647),
            .I(N__6644));
    Span4Mux_v I__1210 (
            .O(N__6644),
            .I(N__6641));
    Sp12to4 I__1209 (
            .O(N__6641),
            .I(N__6638));
    Span12Mux_h I__1208 (
            .O(N__6638),
            .I(N__6635));
    Odrv12 I__1207 (
            .O(N__6635),
            .I(D_LL_AMIGA_in_0));
    IoInMux I__1206 (
            .O(N__6632),
            .I(N__6629));
    LocalMux I__1205 (
            .O(N__6629),
            .I(N__6626));
    Span4Mux_s2_h I__1204 (
            .O(N__6626),
            .I(N__6623));
    Span4Mux_v I__1203 (
            .O(N__6623),
            .I(N__6620));
    Sp12to4 I__1202 (
            .O(N__6620),
            .I(N__6617));
    Span12Mux_h I__1201 (
            .O(N__6617),
            .I(N__6614));
    Odrv12 I__1200 (
            .O(N__6614),
            .I(un2_D_LL_AMIGA_0));
    InMux I__1199 (
            .O(N__6611),
            .I(N__6608));
    LocalMux I__1198 (
            .O(N__6608),
            .I(N__6605));
    Span4Mux_v I__1197 (
            .O(N__6605),
            .I(N__6602));
    Sp12to4 I__1196 (
            .O(N__6602),
            .I(N__6599));
    Span12Mux_h I__1195 (
            .O(N__6599),
            .I(N__6596));
    Odrv12 I__1194 (
            .O(N__6596),
            .I(D_LL_AMIGA_in_2));
    IoInMux I__1193 (
            .O(N__6593),
            .I(N__6590));
    LocalMux I__1192 (
            .O(N__6590),
            .I(N__6587));
    IoSpan4Mux I__1191 (
            .O(N__6587),
            .I(N__6584));
    IoSpan4Mux I__1190 (
            .O(N__6584),
            .I(N__6581));
    Span4Mux_s2_h I__1189 (
            .O(N__6581),
            .I(N__6578));
    Sp12to4 I__1188 (
            .O(N__6578),
            .I(N__6575));
    Span12Mux_h I__1187 (
            .O(N__6575),
            .I(N__6572));
    Odrv12 I__1186 (
            .O(N__6572),
            .I(un2_D_LL_AMIGA_2));
    InMux I__1185 (
            .O(N__6569),
            .I(N__6566));
    LocalMux I__1184 (
            .O(N__6566),
            .I(N__6563));
    Span4Mux_v I__1183 (
            .O(N__6563),
            .I(N__6560));
    Odrv4 I__1182 (
            .O(N__6560),
            .I(READ_CYCLE_ACTIVE_rep26_i_ess));
    IoInMux I__1181 (
            .O(N__6557),
            .I(N__6554));
    LocalMux I__1180 (
            .O(N__6554),
            .I(N__6551));
    Span12Mux_s4_h I__1179 (
            .O(N__6551),
            .I(N__6548));
    Span12Mux_h I__1178 (
            .O(N__6548),
            .I(N__6545));
    Odrv12 I__1177 (
            .O(N__6545),
            .I(N_231_i));
    InMux I__1176 (
            .O(N__6542),
            .I(N__6539));
    LocalMux I__1175 (
            .O(N__6539),
            .I(N__6536));
    Span12Mux_v I__1174 (
            .O(N__6536),
            .I(N__6533));
    Span12Mux_h I__1173 (
            .O(N__6533),
            .I(N__6530));
    Odrv12 I__1172 (
            .O(N__6530),
            .I(D_LL_AMIGA_in_7));
    IoInMux I__1171 (
            .O(N__6527),
            .I(N__6524));
    LocalMux I__1170 (
            .O(N__6524),
            .I(N__6521));
    IoSpan4Mux I__1169 (
            .O(N__6521),
            .I(N__6518));
    Sp12to4 I__1168 (
            .O(N__6518),
            .I(N__6515));
    Span12Mux_s7_h I__1167 (
            .O(N__6515),
            .I(N__6512));
    Span12Mux_v I__1166 (
            .O(N__6512),
            .I(N__6509));
    Odrv12 I__1165 (
            .O(N__6509),
            .I(un2_D_LL_AMIGA_7));
    InMux I__1164 (
            .O(N__6506),
            .I(N__6503));
    LocalMux I__1163 (
            .O(N__6503),
            .I(N__6500));
    Span4Mux_v I__1162 (
            .O(N__6500),
            .I(N__6495));
    InMux I__1161 (
            .O(N__6499),
            .I(N__6492));
    InMux I__1160 (
            .O(N__6498),
            .I(N__6489));
    Odrv4 I__1159 (
            .O(N__6495),
            .I(\U111_CYCLE_SM.LW_TRANSZ0 ));
    LocalMux I__1158 (
            .O(N__6492),
            .I(\U111_CYCLE_SM.LW_TRANSZ0 ));
    LocalMux I__1157 (
            .O(N__6489),
            .I(\U111_CYCLE_SM.LW_TRANSZ0 ));
    CascadeMux I__1156 (
            .O(N__6482),
            .I(N__6478));
    InMux I__1155 (
            .O(N__6481),
            .I(N__6475));
    InMux I__1154 (
            .O(N__6478),
            .I(N__6472));
    LocalMux I__1153 (
            .O(N__6475),
            .I(N__6469));
    LocalMux I__1152 (
            .O(N__6472),
            .I(N__6466));
    Span4Mux_v I__1151 (
            .O(N__6469),
            .I(N__6462));
    Span4Mux_v I__1150 (
            .O(N__6466),
            .I(N__6459));
    InMux I__1149 (
            .O(N__6465),
            .I(N__6456));
    Sp12to4 I__1148 (
            .O(N__6462),
            .I(N__6449));
    Sp12to4 I__1147 (
            .O(N__6459),
            .I(N__6449));
    LocalMux I__1146 (
            .O(N__6456),
            .I(N__6449));
    Span12Mux_h I__1145 (
            .O(N__6449),
            .I(N__6446));
    Span12Mux_v I__1144 (
            .O(N__6446),
            .I(N__6443));
    Odrv12 I__1143 (
            .O(N__6443),
            .I(PORTSIZE_c));
    InMux I__1142 (
            .O(N__6440),
            .I(N__6437));
    LocalMux I__1141 (
            .O(N__6437),
            .I(N__6429));
    InMux I__1140 (
            .O(N__6436),
            .I(N__6424));
    InMux I__1139 (
            .O(N__6435),
            .I(N__6424));
    InMux I__1138 (
            .O(N__6434),
            .I(N__6419));
    InMux I__1137 (
            .O(N__6433),
            .I(N__6419));
    InMux I__1136 (
            .O(N__6432),
            .I(N__6416));
    Odrv4 I__1135 (
            .O(N__6429),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1134 (
            .O(N__6424),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1133 (
            .O(N__6419),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1132 (
            .O(N__6416),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    CascadeMux I__1131 (
            .O(N__6407),
            .I(\U111_CYCLE_SM.N_60_cascade_ ));
    InMux I__1130 (
            .O(N__6404),
            .I(N__6401));
    LocalMux I__1129 (
            .O(N__6401),
            .I(N__6398));
    Span4Mux_v I__1128 (
            .O(N__6398),
            .I(N__6395));
    Odrv4 I__1127 (
            .O(N__6395),
            .I(READ_CYCLE_ACTIVE_rep6_i_ess));
    IoInMux I__1126 (
            .O(N__6392),
            .I(N__6389));
    LocalMux I__1125 (
            .O(N__6389),
            .I(N__6386));
    Span4Mux_s1_v I__1124 (
            .O(N__6386),
            .I(N__6383));
    Span4Mux_v I__1123 (
            .O(N__6383),
            .I(N__6380));
    Sp12to4 I__1122 (
            .O(N__6380),
            .I(N__6377));
    Span12Mux_h I__1121 (
            .O(N__6377),
            .I(N__6374));
    Odrv12 I__1120 (
            .O(N__6374),
            .I(N_211_i));
    CascadeMux I__1119 (
            .O(N__6371),
            .I(\U111_CYCLE_SM.N_75_cascade_ ));
    InMux I__1118 (
            .O(N__6368),
            .I(N__6365));
    LocalMux I__1117 (
            .O(N__6365),
            .I(\U111_CYCLE_SM.LATCH_EN_5 ));
    CascadeMux I__1116 (
            .O(N__6362),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa_cascade_ ));
    InMux I__1115 (
            .O(N__6359),
            .I(N__6352));
    InMux I__1114 (
            .O(N__6358),
            .I(N__6349));
    InMux I__1113 (
            .O(N__6357),
            .I(N__6342));
    InMux I__1112 (
            .O(N__6356),
            .I(N__6342));
    InMux I__1111 (
            .O(N__6355),
            .I(N__6342));
    LocalMux I__1110 (
            .O(N__6352),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    LocalMux I__1109 (
            .O(N__6349),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    LocalMux I__1108 (
            .O(N__6342),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    InMux I__1107 (
            .O(N__6335),
            .I(N__6329));
    InMux I__1106 (
            .O(N__6334),
            .I(N__6329));
    LocalMux I__1105 (
            .O(N__6329),
            .I(N__6326));
    Span4Mux_h I__1104 (
            .O(N__6326),
            .I(N__6323));
    Sp12to4 I__1103 (
            .O(N__6323),
            .I(N__6320));
    Span12Mux_v I__1102 (
            .O(N__6320),
            .I(N__6317));
    Span12Mux_h I__1101 (
            .O(N__6317),
            .I(N__6314));
    Odrv12 I__1100 (
            .O(N__6314),
            .I(SIZ_c_1));
    CascadeMux I__1099 (
            .O(N__6311),
            .I(N__6307));
    CascadeMux I__1098 (
            .O(N__6310),
            .I(N__6304));
    InMux I__1097 (
            .O(N__6307),
            .I(N__6301));
    InMux I__1096 (
            .O(N__6304),
            .I(N__6298));
    LocalMux I__1095 (
            .O(N__6301),
            .I(N__6293));
    LocalMux I__1094 (
            .O(N__6298),
            .I(N__6293));
    Span4Mux_v I__1093 (
            .O(N__6293),
            .I(N__6290));
    Span4Mux_v I__1092 (
            .O(N__6290),
            .I(N__6287));
    Sp12to4 I__1091 (
            .O(N__6287),
            .I(N__6284));
    Span12Mux_h I__1090 (
            .O(N__6284),
            .I(N__6281));
    Odrv12 I__1089 (
            .O(N__6281),
            .I(SIZ_c_0));
    InMux I__1088 (
            .O(N__6278),
            .I(N__6275));
    LocalMux I__1087 (
            .O(N__6275),
            .I(N__6272));
    Odrv12 I__1086 (
            .O(N__6272),
            .I(WRITE_CYCLE_ACTIVE_rep9_i_ess));
    InMux I__1085 (
            .O(N__6269),
            .I(N__6266));
    LocalMux I__1084 (
            .O(N__6266),
            .I(N__6263));
    Odrv12 I__1083 (
            .O(N__6263),
            .I(WRITE_CYCLE_ACTIVE_rep13_i_ess));
    InMux I__1082 (
            .O(N__6260),
            .I(N__6257));
    LocalMux I__1081 (
            .O(N__6257),
            .I(N__6254));
    Span4Mux_v I__1080 (
            .O(N__6254),
            .I(N__6251));
    Odrv4 I__1079 (
            .O(N__6251),
            .I(WRITE_CYCLE_ACTIVE_rep6_i_ess));
    IoInMux I__1078 (
            .O(N__6248),
            .I(N__6245));
    LocalMux I__1077 (
            .O(N__6245),
            .I(N__6242));
    Span4Mux_s3_v I__1076 (
            .O(N__6242),
            .I(N__6239));
    Odrv4 I__1075 (
            .O(N__6239),
            .I(LBENn_c_i_0));
    InMux I__1074 (
            .O(N__6236),
            .I(N__6233));
    LocalMux I__1073 (
            .O(N__6233),
            .I(\U111_CYCLE_SM.N_33 ));
    InMux I__1072 (
            .O(N__6230),
            .I(N__6227));
    LocalMux I__1071 (
            .O(N__6227),
            .I(\U111_CYCLE_SM.N_49 ));
    InMux I__1070 (
            .O(N__6224),
            .I(N__6221));
    LocalMux I__1069 (
            .O(N__6221),
            .I(\U111_CYCLE_SM.N_75 ));
    InMux I__1068 (
            .O(N__6218),
            .I(N__6215));
    LocalMux I__1067 (
            .O(N__6215),
            .I(N__6212));
    Span12Mux_h I__1066 (
            .O(N__6212),
            .I(N__6209));
    Span12Mux_v I__1065 (
            .O(N__6209),
            .I(N__6206));
    Odrv12 I__1064 (
            .O(N__6206),
            .I(TS_CPUn_c));
    InMux I__1063 (
            .O(N__6203),
            .I(N__6200));
    LocalMux I__1062 (
            .O(N__6200),
            .I(N__6197));
    Span4Mux_h I__1061 (
            .O(N__6197),
            .I(N__6194));
    Sp12to4 I__1060 (
            .O(N__6194),
            .I(N__6191));
    Span12Mux_h I__1059 (
            .O(N__6191),
            .I(N__6188));
    Odrv12 I__1058 (
            .O(N__6188),
            .I(BGn_c));
    InMux I__1057 (
            .O(N__6185),
            .I(N__6181));
    InMux I__1056 (
            .O(N__6184),
            .I(N__6178));
    LocalMux I__1055 (
            .O(N__6181),
            .I(\U111_CYCLE_SM.TS_DELAYZ0 ));
    LocalMux I__1054 (
            .O(N__6178),
            .I(\U111_CYCLE_SM.TS_DELAYZ0 ));
    InMux I__1053 (
            .O(N__6173),
            .I(N__6170));
    LocalMux I__1052 (
            .O(N__6170),
            .I(N__6167));
    Span4Mux_v I__1051 (
            .O(N__6167),
            .I(N__6164));
    Span4Mux_h I__1050 (
            .O(N__6164),
            .I(N__6161));
    Odrv4 I__1049 (
            .O(N__6161),
            .I(WRITE_CYCLE_ACTIVE_rep11_i_ess));
    InMux I__1048 (
            .O(N__6158),
            .I(N__6155));
    LocalMux I__1047 (
            .O(N__6155),
            .I(N__6152));
    Span4Mux_v I__1046 (
            .O(N__6152),
            .I(N__6149));
    Span4Mux_h I__1045 (
            .O(N__6149),
            .I(N__6146));
    Odrv4 I__1044 (
            .O(N__6146),
            .I(WRITE_CYCLE_ACTIVE_rep5_i_ess));
    InMux I__1043 (
            .O(N__6143),
            .I(N__6140));
    LocalMux I__1042 (
            .O(N__6140),
            .I(N__6137));
    Odrv12 I__1041 (
            .O(N__6137),
            .I(WRITE_CYCLE_ACTIVE_rep15_i_ess));
    IoInMux I__1040 (
            .O(N__6134),
            .I(N__6130));
    IoInMux I__1039 (
            .O(N__6133),
            .I(N__6127));
    LocalMux I__1038 (
            .O(N__6130),
            .I(N__6124));
    LocalMux I__1037 (
            .O(N__6127),
            .I(N__6119));
    Span4Mux_s2_v I__1036 (
            .O(N__6124),
            .I(N__6116));
    IoInMux I__1035 (
            .O(N__6123),
            .I(N__6113));
    IoInMux I__1034 (
            .O(N__6122),
            .I(N__6110));
    IoSpan4Mux I__1033 (
            .O(N__6119),
            .I(N__6107));
    Span4Mux_h I__1032 (
            .O(N__6116),
            .I(N__6104));
    LocalMux I__1031 (
            .O(N__6113),
            .I(N__6101));
    LocalMux I__1030 (
            .O(N__6110),
            .I(N__6098));
    Span4Mux_s3_h I__1029 (
            .O(N__6107),
            .I(N__6095));
    Span4Mux_h I__1028 (
            .O(N__6104),
            .I(N__6090));
    Span4Mux_s2_v I__1027 (
            .O(N__6101),
            .I(N__6090));
    IoSpan4Mux I__1026 (
            .O(N__6098),
            .I(N__6087));
    Span4Mux_h I__1025 (
            .O(N__6095),
            .I(N__6084));
    Span4Mux_v I__1024 (
            .O(N__6090),
            .I(N__6081));
    Span4Mux_s3_h I__1023 (
            .O(N__6087),
            .I(N__6078));
    Span4Mux_h I__1022 (
            .O(N__6084),
            .I(N__6075));
    Span4Mux_v I__1021 (
            .O(N__6081),
            .I(N__6072));
    Span4Mux_h I__1020 (
            .O(N__6078),
            .I(N__6069));
    Span4Mux_h I__1019 (
            .O(N__6075),
            .I(N__6066));
    Span4Mux_v I__1018 (
            .O(N__6072),
            .I(N__6061));
    Span4Mux_h I__1017 (
            .O(N__6069),
            .I(N__6061));
    Odrv4 I__1016 (
            .O(N__6066),
            .I(GB_BUFFER_CLK40_THRU_CO));
    Odrv4 I__1015 (
            .O(N__6061),
            .I(GB_BUFFER_CLK40_THRU_CO));
    InMux I__1014 (
            .O(N__6056),
            .I(N__6053));
    LocalMux I__1013 (
            .O(N__6053),
            .I(N__6050));
    Span4Mux_v I__1012 (
            .O(N__6050),
            .I(N__6047));
    Odrv4 I__1011 (
            .O(N__6047),
            .I(WRITE_CYCLE_ACTIVE_rep24_i_ess));
    InMux I__1010 (
            .O(N__6044),
            .I(N__6038));
    InMux I__1009 (
            .O(N__6043),
            .I(N__6038));
    LocalMux I__1008 (
            .O(N__6038),
            .I(N__6035));
    Span12Mux_h I__1007 (
            .O(N__6035),
            .I(N__6031));
    InMux I__1006 (
            .O(N__6034),
            .I(N__6028));
    Odrv12 I__1005 (
            .O(N__6031),
            .I(\U111_CYCLE_SM.A2_ENZ0 ));
    LocalMux I__1004 (
            .O(N__6028),
            .I(\U111_CYCLE_SM.A2_ENZ0 ));
    InMux I__1003 (
            .O(N__6023),
            .I(N__6020));
    LocalMux I__1002 (
            .O(N__6020),
            .I(N__6017));
    Span4Mux_v I__1001 (
            .O(N__6017),
            .I(N__6014));
    Span4Mux_h I__1000 (
            .O(N__6014),
            .I(N__6011));
    Odrv4 I__999 (
            .O(N__6011),
            .I(\U111_CYCLE_SM.N_67 ));
    InMux I__998 (
            .O(N__6008),
            .I(N__6004));
    InMux I__997 (
            .O(N__6007),
            .I(N__6001));
    LocalMux I__996 (
            .O(N__6004),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    LocalMux I__995 (
            .O(N__6001),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    IoInMux I__994 (
            .O(N__5996),
            .I(N__5993));
    LocalMux I__993 (
            .O(N__5993),
            .I(N__5990));
    IoSpan4Mux I__992 (
            .O(N__5990),
            .I(N__5987));
    Span4Mux_s2_h I__991 (
            .O(N__5987),
            .I(N__5983));
    InMux I__990 (
            .O(N__5986),
            .I(N__5980));
    Span4Mux_v I__989 (
            .O(N__5983),
            .I(N__5977));
    LocalMux I__988 (
            .O(N__5980),
            .I(N__5974));
    Sp12to4 I__987 (
            .O(N__5977),
            .I(N__5971));
    Sp12to4 I__986 (
            .O(N__5974),
            .I(N__5968));
    Span12Mux_s9_h I__985 (
            .O(N__5971),
            .I(N__5965));
    Span12Mux_v I__984 (
            .O(N__5968),
            .I(N__5962));
    Span12Mux_h I__983 (
            .O(N__5965),
            .I(N__5959));
    Span12Mux_h I__982 (
            .O(N__5962),
            .I(N__5956));
    Odrv12 I__981 (
            .O(N__5959),
            .I(D_LM_040_in_5));
    Odrv12 I__980 (
            .O(N__5956),
            .I(D_LM_040_in_5));
    InMux I__979 (
            .O(N__5951),
            .I(N__5948));
    LocalMux I__978 (
            .O(N__5948),
            .I(N__5945));
    Span4Mux_v I__977 (
            .O(N__5945),
            .I(N__5942));
    Span4Mux_h I__976 (
            .O(N__5942),
            .I(N__5939));
    Sp12to4 I__975 (
            .O(N__5939),
            .I(N__5936));
    Span12Mux_h I__974 (
            .O(N__5936),
            .I(N__5933));
    Odrv12 I__973 (
            .O(N__5933),
            .I(D_UU_040_in_5));
    IoInMux I__972 (
            .O(N__5930),
            .I(N__5927));
    LocalMux I__971 (
            .O(N__5927),
            .I(N__5924));
    Span4Mux_s3_h I__970 (
            .O(N__5924),
            .I(N__5921));
    Span4Mux_h I__969 (
            .O(N__5921),
            .I(N__5918));
    Span4Mux_h I__968 (
            .O(N__5918),
            .I(N__5915));
    Span4Mux_v I__967 (
            .O(N__5915),
            .I(N__5912));
    Odrv4 I__966 (
            .O(N__5912),
            .I(un1_D_UU_040_5));
    IoInMux I__965 (
            .O(N__5909),
            .I(N__5906));
    LocalMux I__964 (
            .O(N__5906),
            .I(N__5903));
    IoSpan4Mux I__963 (
            .O(N__5903),
            .I(N__5899));
    InMux I__962 (
            .O(N__5902),
            .I(N__5896));
    IoSpan4Mux I__961 (
            .O(N__5899),
            .I(N__5893));
    LocalMux I__960 (
            .O(N__5896),
            .I(N__5890));
    Span4Mux_s2_h I__959 (
            .O(N__5893),
            .I(N__5887));
    Span4Mux_v I__958 (
            .O(N__5890),
            .I(N__5884));
    Sp12to4 I__957 (
            .O(N__5887),
            .I(N__5881));
    Sp12to4 I__956 (
            .O(N__5884),
            .I(N__5878));
    Span12Mux_h I__955 (
            .O(N__5881),
            .I(N__5873));
    Span12Mux_v I__954 (
            .O(N__5878),
            .I(N__5873));
    Span12Mux_h I__953 (
            .O(N__5873),
            .I(N__5870));
    Odrv12 I__952 (
            .O(N__5870),
            .I(D_LM_040_in_3));
    InMux I__951 (
            .O(N__5867),
            .I(N__5864));
    LocalMux I__950 (
            .O(N__5864),
            .I(N__5861));
    Span4Mux_v I__949 (
            .O(N__5861),
            .I(N__5858));
    Span4Mux_h I__948 (
            .O(N__5858),
            .I(N__5855));
    Sp12to4 I__947 (
            .O(N__5855),
            .I(N__5852));
    Span12Mux_h I__946 (
            .O(N__5852),
            .I(N__5849));
    Odrv12 I__945 (
            .O(N__5849),
            .I(D_UU_040_in_3));
    IoInMux I__944 (
            .O(N__5846),
            .I(N__5843));
    LocalMux I__943 (
            .O(N__5843),
            .I(N__5840));
    IoSpan4Mux I__942 (
            .O(N__5840),
            .I(N__5837));
    Sp12to4 I__941 (
            .O(N__5837),
            .I(N__5834));
    Span12Mux_s6_v I__940 (
            .O(N__5834),
            .I(N__5831));
    Odrv12 I__939 (
            .O(N__5831),
            .I(un1_D_UU_040_3));
    InMux I__938 (
            .O(N__5828),
            .I(N__5825));
    LocalMux I__937 (
            .O(N__5825),
            .I(N__5822));
    Span4Mux_v I__936 (
            .O(N__5822),
            .I(N__5819));
    Sp12to4 I__935 (
            .O(N__5819),
            .I(N__5816));
    Span12Mux_h I__934 (
            .O(N__5816),
            .I(N__5813));
    Odrv12 I__933 (
            .O(N__5813),
            .I(D_LL_AMIGA_in_3));
    IoInMux I__932 (
            .O(N__5810),
            .I(N__5807));
    LocalMux I__931 (
            .O(N__5807),
            .I(N__5804));
    IoSpan4Mux I__930 (
            .O(N__5804),
            .I(N__5801));
    Span4Mux_s1_h I__929 (
            .O(N__5801),
            .I(N__5798));
    Span4Mux_v I__928 (
            .O(N__5798),
            .I(N__5795));
    Sp12to4 I__927 (
            .O(N__5795),
            .I(N__5792));
    Span12Mux_s10_h I__926 (
            .O(N__5792),
            .I(N__5789));
    Odrv12 I__925 (
            .O(N__5789),
            .I(un2_D_LL_AMIGA_3));
    InMux I__924 (
            .O(N__5786),
            .I(N__5783));
    LocalMux I__923 (
            .O(N__5783),
            .I(N__5780));
    Span4Mux_v I__922 (
            .O(N__5780),
            .I(N__5777));
    Sp12to4 I__921 (
            .O(N__5777),
            .I(N__5774));
    Odrv12 I__920 (
            .O(N__5774),
            .I(WRITE_CYCLE_ACTIVE_rep30_i_ess));
    InMux I__919 (
            .O(N__5771),
            .I(N__5768));
    LocalMux I__918 (
            .O(N__5768),
            .I(N__5765));
    Span4Mux_v I__917 (
            .O(N__5765),
            .I(N__5762));
    Span4Mux_h I__916 (
            .O(N__5762),
            .I(N__5759));
    Odrv4 I__915 (
            .O(N__5759),
            .I(WRITE_CYCLE_ACTIVE_rep14_i_ess));
    InMux I__914 (
            .O(N__5756),
            .I(N__5753));
    LocalMux I__913 (
            .O(N__5753),
            .I(N__5750));
    Span4Mux_v I__912 (
            .O(N__5750),
            .I(N__5747));
    Odrv4 I__911 (
            .O(N__5747),
            .I(WRITE_CYCLE_ACTIVE_rep1_i_ess));
    InMux I__910 (
            .O(N__5744),
            .I(N__5741));
    LocalMux I__909 (
            .O(N__5741),
            .I(N__5738));
    Span4Mux_v I__908 (
            .O(N__5738),
            .I(N__5735));
    Odrv4 I__907 (
            .O(N__5735),
            .I(WRITE_CYCLE_ACTIVE_rep23_i_ess));
    InMux I__906 (
            .O(N__5732),
            .I(N__5729));
    LocalMux I__905 (
            .O(N__5729),
            .I(N__5726));
    Span4Mux_h I__904 (
            .O(N__5726),
            .I(N__5723));
    Span4Mux_v I__903 (
            .O(N__5723),
            .I(N__5720));
    Span4Mux_h I__902 (
            .O(N__5720),
            .I(N__5717));
    Odrv4 I__901 (
            .O(N__5717),
            .I(WRITE_CYCLE_ACTIVE_rep29_i_ess));
    InMux I__900 (
            .O(N__5714),
            .I(N__5711));
    LocalMux I__899 (
            .O(N__5711),
            .I(N__5708));
    Span4Mux_v I__898 (
            .O(N__5708),
            .I(N__5705));
    Odrv4 I__897 (
            .O(N__5705),
            .I(WRITE_CYCLE_ACTIVE_rep3_i_ess));
    InMux I__896 (
            .O(N__5702),
            .I(N__5699));
    LocalMux I__895 (
            .O(N__5699),
            .I(N__5696));
    Span4Mux_h I__894 (
            .O(N__5696),
            .I(N__5693));
    Odrv4 I__893 (
            .O(N__5693),
            .I(WRITE_CYCLE_ACTIVE_rep4_i_ess));
    InMux I__892 (
            .O(N__5690),
            .I(N__5687));
    LocalMux I__891 (
            .O(N__5687),
            .I(N__5684));
    Odrv12 I__890 (
            .O(N__5684),
            .I(WRITE_CYCLE_ACTIVE_rep12_i_ess));
    InMux I__889 (
            .O(N__5681),
            .I(N__5678));
    LocalMux I__888 (
            .O(N__5678),
            .I(WRITE_CYCLE_ACTIVE_rep7_i_ess));
    IoInMux I__887 (
            .O(N__5675),
            .I(N__5672));
    LocalMux I__886 (
            .O(N__5672),
            .I(N__5669));
    IoSpan4Mux I__885 (
            .O(N__5669),
            .I(N__5666));
    Span4Mux_s1_v I__884 (
            .O(N__5666),
            .I(N__5663));
    Sp12to4 I__883 (
            .O(N__5663),
            .I(N__5660));
    Span12Mux_s9_v I__882 (
            .O(N__5660),
            .I(N__5657));
    Odrv12 I__881 (
            .O(N__5657),
            .I(N_244_i));
    InMux I__880 (
            .O(N__5654),
            .I(N__5651));
    LocalMux I__879 (
            .O(N__5651),
            .I(N__5648));
    Span4Mux_h I__878 (
            .O(N__5648),
            .I(N__5645));
    Span4Mux_v I__877 (
            .O(N__5645),
            .I(N__5642));
    Odrv4 I__876 (
            .O(N__5642),
            .I(WRITE_CYCLE_ACTIVE_rep28_i_ess));
    InMux I__875 (
            .O(N__5639),
            .I(N__5636));
    LocalMux I__874 (
            .O(N__5636),
            .I(N__5633));
    Odrv12 I__873 (
            .O(N__5633),
            .I(WRITE_CYCLE_ACTIVE_i_ess));
    InMux I__872 (
            .O(N__5630),
            .I(N__5627));
    LocalMux I__871 (
            .O(N__5627),
            .I(N__5624));
    Odrv4 I__870 (
            .O(N__5624),
            .I(WRITE_CYCLE_ACTIVE_rep18_i_ess));
    InMux I__869 (
            .O(N__5621),
            .I(N__5618));
    LocalMux I__868 (
            .O(N__5618),
            .I(N__5615));
    Span12Mux_s6_h I__867 (
            .O(N__5615),
            .I(N__5612));
    Odrv12 I__866 (
            .O(N__5612),
            .I(WRITE_CYCLE_ACTIVE_rep10_i_ess));
    InMux I__865 (
            .O(N__5609),
            .I(N__5606));
    LocalMux I__864 (
            .O(N__5606),
            .I(N__5603));
    Span4Mux_h I__863 (
            .O(N__5603),
            .I(N__5600));
    Sp12to4 I__862 (
            .O(N__5600),
            .I(N__5597));
    Odrv12 I__861 (
            .O(N__5597),
            .I(WRITE_CYCLE_ACTIVE_rep26_i_ess));
    InMux I__860 (
            .O(N__5594),
            .I(N__5591));
    LocalMux I__859 (
            .O(N__5591),
            .I(N__5588));
    Span4Mux_v I__858 (
            .O(N__5588),
            .I(N__5585));
    Odrv4 I__857 (
            .O(N__5585),
            .I(WRITE_CYCLE_ACTIVE_rep22_i_ess));
    InMux I__856 (
            .O(N__5582),
            .I(N__5579));
    LocalMux I__855 (
            .O(N__5579),
            .I(N__5576));
    Sp12to4 I__854 (
            .O(N__5576),
            .I(N__5573));
    Span12Mux_v I__853 (
            .O(N__5573),
            .I(N__5570));
    Odrv12 I__852 (
            .O(N__5570),
            .I(WRITE_CYCLE_ACTIVE_rep0_i_ess));
    InMux I__851 (
            .O(N__5567),
            .I(N__5564));
    LocalMux I__850 (
            .O(N__5564),
            .I(N__5561));
    Span4Mux_v I__849 (
            .O(N__5561),
            .I(N__5558));
    Span4Mux_h I__848 (
            .O(N__5558),
            .I(N__5555));
    Odrv4 I__847 (
            .O(N__5555),
            .I(WRITE_CYCLE_ACTIVE_rep21_i_ess));
    InMux I__846 (
            .O(N__5552),
            .I(N__5549));
    LocalMux I__845 (
            .O(N__5549),
            .I(N__5546));
    Span4Mux_h I__844 (
            .O(N__5546),
            .I(N__5543));
    Span4Mux_v I__843 (
            .O(N__5543),
            .I(N__5540));
    Odrv4 I__842 (
            .O(N__5540),
            .I(WRITE_CYCLE_ACTIVE_rep2_i_ess));
    IoInMux I__841 (
            .O(N__5537),
            .I(N__5534));
    LocalMux I__840 (
            .O(N__5534),
            .I(N__5531));
    IoSpan4Mux I__839 (
            .O(N__5531),
            .I(N__5528));
    Sp12to4 I__838 (
            .O(N__5528),
            .I(N__5525));
    Span12Mux_s7_h I__837 (
            .O(N__5525),
            .I(N__5522));
    Span12Mux_h I__836 (
            .O(N__5522),
            .I(N__5519));
    Odrv12 I__835 (
            .O(N__5519),
            .I(un2_D_LM_AMIGA_0));
    IoInMux I__834 (
            .O(N__5516),
            .I(N__5513));
    LocalMux I__833 (
            .O(N__5513),
            .I(N__5510));
    Span4Mux_s3_h I__832 (
            .O(N__5510),
            .I(N__5507));
    Span4Mux_v I__831 (
            .O(N__5507),
            .I(N__5504));
    Span4Mux_h I__830 (
            .O(N__5504),
            .I(N__5501));
    Span4Mux_h I__829 (
            .O(N__5501),
            .I(N__5498));
    Odrv4 I__828 (
            .O(N__5498),
            .I(N_268_i));
    IoInMux I__827 (
            .O(N__5495),
            .I(N__5492));
    LocalMux I__826 (
            .O(N__5492),
            .I(N__5489));
    Span12Mux_s11_h I__825 (
            .O(N__5489),
            .I(N__5486));
    Odrv12 I__824 (
            .O(N__5486),
            .I(N_255_i));
    IoInMux I__823 (
            .O(N__5483),
            .I(N__5480));
    LocalMux I__822 (
            .O(N__5480),
            .I(N__5477));
    IoSpan4Mux I__821 (
            .O(N__5477),
            .I(N__5474));
    Span4Mux_s1_v I__820 (
            .O(N__5474),
            .I(N__5471));
    Sp12to4 I__819 (
            .O(N__5471),
            .I(N__5468));
    Span12Mux_v I__818 (
            .O(N__5468),
            .I(N__5465));
    Odrv12 I__817 (
            .O(N__5465),
            .I(TSn_c));
    InMux I__816 (
            .O(N__5462),
            .I(N__5459));
    LocalMux I__815 (
            .O(N__5459),
            .I(N__5456));
    Span12Mux_s8_h I__814 (
            .O(N__5456),
            .I(N__5453));
    Odrv12 I__813 (
            .O(N__5453),
            .I(WRITE_CYCLE_ACTIVE_rep17_i_ess));
    InMux I__812 (
            .O(N__5450),
            .I(N__5447));
    LocalMux I__811 (
            .O(N__5447),
            .I(N__5444));
    Span4Mux_v I__810 (
            .O(N__5444),
            .I(N__5441));
    Odrv4 I__809 (
            .O(N__5441),
            .I(WRITE_CYCLE_ACTIVE_rep19_i_ess));
    InMux I__808 (
            .O(N__5438),
            .I(N__5435));
    LocalMux I__807 (
            .O(N__5435),
            .I(N__5432));
    Span4Mux_v I__806 (
            .O(N__5432),
            .I(N__5429));
    Odrv4 I__805 (
            .O(N__5429),
            .I(WRITE_CYCLE_ACTIVE_rep8_i_ess));
    InMux I__804 (
            .O(N__5426),
            .I(N__5423));
    LocalMux I__803 (
            .O(N__5423),
            .I(N__5420));
    Span4Mux_v I__802 (
            .O(N__5420),
            .I(N__5417));
    Span4Mux_h I__801 (
            .O(N__5417),
            .I(N__5414));
    Odrv4 I__800 (
            .O(N__5414),
            .I(WRITE_CYCLE_ACTIVE_rep25_i_ess));
    InMux I__799 (
            .O(N__5411),
            .I(N__5408));
    LocalMux I__798 (
            .O(N__5408),
            .I(N__5405));
    Span12Mux_h I__797 (
            .O(N__5405),
            .I(N__5402));
    Odrv12 I__796 (
            .O(N__5402),
            .I(WRITE_CYCLE_ACTIVE_rep27_i_ess));
    IoInMux I__795 (
            .O(N__5399),
            .I(N__5396));
    LocalMux I__794 (
            .O(N__5396),
            .I(N__5393));
    Span4Mux_s2_v I__793 (
            .O(N__5393),
            .I(N__5390));
    Span4Mux_h I__792 (
            .O(N__5390),
            .I(N__5387));
    Span4Mux_v I__791 (
            .O(N__5387),
            .I(N__5384));
    Odrv4 I__790 (
            .O(N__5384),
            .I(N_237_i));
    IoInMux I__789 (
            .O(N__5381),
            .I(N__5377));
    InMux I__788 (
            .O(N__5380),
            .I(N__5374));
    LocalMux I__787 (
            .O(N__5377),
            .I(N__5371));
    LocalMux I__786 (
            .O(N__5374),
            .I(N__5368));
    IoSpan4Mux I__785 (
            .O(N__5371),
            .I(N__5365));
    Span4Mux_v I__784 (
            .O(N__5368),
            .I(N__5362));
    IoSpan4Mux I__783 (
            .O(N__5365),
            .I(N__5359));
    Sp12to4 I__782 (
            .O(N__5362),
            .I(N__5356));
    Span4Mux_s2_h I__781 (
            .O(N__5359),
            .I(N__5353));
    Span12Mux_h I__780 (
            .O(N__5356),
            .I(N__5350));
    Sp12to4 I__779 (
            .O(N__5353),
            .I(N__5347));
    Span12Mux_v I__778 (
            .O(N__5350),
            .I(N__5344));
    Span12Mux_h I__777 (
            .O(N__5347),
            .I(N__5341));
    Span12Mux_v I__776 (
            .O(N__5344),
            .I(N__5338));
    Span12Mux_h I__775 (
            .O(N__5341),
            .I(N__5335));
    Odrv12 I__774 (
            .O(N__5338),
            .I(D_LM_040_in_0));
    Odrv12 I__773 (
            .O(N__5335),
            .I(D_LM_040_in_0));
    InMux I__772 (
            .O(N__5330),
            .I(N__5327));
    LocalMux I__771 (
            .O(N__5327),
            .I(N__5324));
    Span4Mux_v I__770 (
            .O(N__5324),
            .I(N__5321));
    Span4Mux_h I__769 (
            .O(N__5321),
            .I(N__5318));
    Sp12to4 I__768 (
            .O(N__5318),
            .I(N__5315));
    Span12Mux_h I__767 (
            .O(N__5315),
            .I(N__5312));
    Odrv12 I__766 (
            .O(N__5312),
            .I(D_UU_040_in_0));
    IoInMux I__765 (
            .O(N__5309),
            .I(N__5306));
    LocalMux I__764 (
            .O(N__5306),
            .I(N__5303));
    Span4Mux_s2_v I__763 (
            .O(N__5303),
            .I(N__5300));
    Span4Mux_h I__762 (
            .O(N__5300),
            .I(N__5297));
    Span4Mux_v I__761 (
            .O(N__5297),
            .I(N__5294));
    Odrv4 I__760 (
            .O(N__5294),
            .I(un1_D_UU_040_0));
    IoInMux I__759 (
            .O(N__5291),
            .I(N__5288));
    LocalMux I__758 (
            .O(N__5288),
            .I(N__5285));
    IoSpan4Mux I__757 (
            .O(N__5285),
            .I(N__5281));
    IoInMux I__756 (
            .O(N__5284),
            .I(N__5278));
    IoSpan4Mux I__755 (
            .O(N__5281),
            .I(N__5275));
    LocalMux I__754 (
            .O(N__5278),
            .I(N__5272));
    IoSpan4Mux I__753 (
            .O(N__5275),
            .I(N__5267));
    IoSpan4Mux I__752 (
            .O(N__5272),
            .I(N__5267));
    Span4Mux_s3_v I__751 (
            .O(N__5267),
            .I(N__5264));
    Odrv4 I__750 (
            .O(N__5264),
            .I(CONSTANT_ONE_NET));
    InMux I__749 (
            .O(N__5261),
            .I(N__5258));
    LocalMux I__748 (
            .O(N__5258),
            .I(N__5255));
    Span12Mux_v I__747 (
            .O(N__5255),
            .I(N__5252));
    Odrv12 I__746 (
            .O(N__5252),
            .I(D_LL_AMIGA_in_6));
    IoInMux I__745 (
            .O(N__5249),
            .I(N__5246));
    LocalMux I__744 (
            .O(N__5246),
            .I(N__5243));
    Span4Mux_s0_h I__743 (
            .O(N__5243),
            .I(N__5240));
    Sp12to4 I__742 (
            .O(N__5240),
            .I(N__5237));
    Span12Mux_s11_v I__741 (
            .O(N__5237),
            .I(N__5234));
    Span12Mux_h I__740 (
            .O(N__5234),
            .I(N__5231));
    Odrv12 I__739 (
            .O(N__5231),
            .I(un2_D_LL_AMIGA_6));
    InMux I__738 (
            .O(N__5228),
            .I(N__5225));
    LocalMux I__737 (
            .O(N__5225),
            .I(N__5222));
    Span12Mux_h I__736 (
            .O(N__5222),
            .I(N__5219));
    Odrv12 I__735 (
            .O(N__5219),
            .I(D_LM_AMIGA_in_1));
    IoInMux I__734 (
            .O(N__5216),
            .I(N__5213));
    LocalMux I__733 (
            .O(N__5213),
            .I(N__5210));
    Span12Mux_s8_h I__732 (
            .O(N__5210),
            .I(N__5207));
    Span12Mux_h I__731 (
            .O(N__5207),
            .I(N__5204));
    Odrv12 I__730 (
            .O(N__5204),
            .I(un2_D_LM_AMIGA_1));
    InMux I__729 (
            .O(N__5201),
            .I(N__5198));
    LocalMux I__728 (
            .O(N__5198),
            .I(N__5195));
    Span4Mux_v I__727 (
            .O(N__5195),
            .I(N__5192));
    Sp12to4 I__726 (
            .O(N__5192),
            .I(N__5189));
    Span12Mux_h I__725 (
            .O(N__5189),
            .I(N__5186));
    Odrv12 I__724 (
            .O(N__5186),
            .I(D_LM_AMIGA_in_3));
    IoInMux I__723 (
            .O(N__5183),
            .I(N__5180));
    LocalMux I__722 (
            .O(N__5180),
            .I(N__5177));
    IoSpan4Mux I__721 (
            .O(N__5177),
            .I(N__5174));
    Span4Mux_s3_h I__720 (
            .O(N__5174),
            .I(N__5171));
    Span4Mux_v I__719 (
            .O(N__5171),
            .I(N__5168));
    Span4Mux_h I__718 (
            .O(N__5168),
            .I(N__5165));
    Sp12to4 I__717 (
            .O(N__5165),
            .I(N__5162));
    Odrv12 I__716 (
            .O(N__5162),
            .I(un2_D_LM_AMIGA_3));
    IoInMux I__715 (
            .O(N__5159),
            .I(N__5156));
    LocalMux I__714 (
            .O(N__5156),
            .I(N__5153));
    IoSpan4Mux I__713 (
            .O(N__5153),
            .I(N__5150));
    Span4Mux_s3_v I__712 (
            .O(N__5150),
            .I(N__5147));
    Span4Mux_v I__711 (
            .O(N__5147),
            .I(N__5144));
    Odrv4 I__710 (
            .O(N__5144),
            .I(LBENn_c_i));
    InMux I__709 (
            .O(N__5141),
            .I(N__5138));
    LocalMux I__708 (
            .O(N__5138),
            .I(N__5134));
    IoInMux I__707 (
            .O(N__5137),
            .I(N__5131));
    Span4Mux_v I__706 (
            .O(N__5134),
            .I(N__5128));
    LocalMux I__705 (
            .O(N__5131),
            .I(N__5125));
    Span4Mux_h I__704 (
            .O(N__5128),
            .I(N__5122));
    Span12Mux_s5_h I__703 (
            .O(N__5125),
            .I(N__5119));
    Span4Mux_v I__702 (
            .O(N__5122),
            .I(N__5116));
    Span12Mux_h I__701 (
            .O(N__5119),
            .I(N__5113));
    Sp12to4 I__700 (
            .O(N__5116),
            .I(N__5110));
    Span12Mux_v I__699 (
            .O(N__5113),
            .I(N__5107));
    Span12Mux_h I__698 (
            .O(N__5110),
            .I(N__5104));
    Span12Mux_h I__697 (
            .O(N__5107),
            .I(N__5099));
    Span12Mux_v I__696 (
            .O(N__5104),
            .I(N__5099));
    Odrv12 I__695 (
            .O(N__5099),
            .I(D_LM_040_in_2));
    InMux I__694 (
            .O(N__5096),
            .I(N__5093));
    LocalMux I__693 (
            .O(N__5093),
            .I(N__5090));
    Span4Mux_v I__692 (
            .O(N__5090),
            .I(N__5087));
    Span4Mux_h I__691 (
            .O(N__5087),
            .I(N__5084));
    Sp12to4 I__690 (
            .O(N__5084),
            .I(N__5081));
    Span12Mux_h I__689 (
            .O(N__5081),
            .I(N__5078));
    Odrv12 I__688 (
            .O(N__5078),
            .I(D_UU_040_in_2));
    IoInMux I__687 (
            .O(N__5075),
            .I(N__5072));
    LocalMux I__686 (
            .O(N__5072),
            .I(N__5069));
    IoSpan4Mux I__685 (
            .O(N__5069),
            .I(N__5066));
    Span4Mux_s2_v I__684 (
            .O(N__5066),
            .I(N__5063));
    Span4Mux_v I__683 (
            .O(N__5063),
            .I(N__5060));
    Odrv4 I__682 (
            .O(N__5060),
            .I(un1_D_UU_040_2));
    InMux I__681 (
            .O(N__5057),
            .I(N__5054));
    LocalMux I__680 (
            .O(N__5054),
            .I(N__5051));
    Span4Mux_v I__679 (
            .O(N__5051),
            .I(N__5048));
    Sp12to4 I__678 (
            .O(N__5048),
            .I(N__5045));
    Span12Mux_h I__677 (
            .O(N__5045),
            .I(N__5042));
    Odrv12 I__676 (
            .O(N__5042),
            .I(D_LM_AMIGA_in_0));
    IoInMux I__675 (
            .O(N__5039),
            .I(N__5036));
    LocalMux I__674 (
            .O(N__5036),
            .I(N__5033));
    Span12Mux_s5_h I__673 (
            .O(N__5033),
            .I(N__5030));
    Odrv12 I__672 (
            .O(N__5030),
            .I(N_256_i));
    InMux I__671 (
            .O(N__5027),
            .I(N__5024));
    LocalMux I__670 (
            .O(N__5024),
            .I(N__5021));
    Odrv12 I__669 (
            .O(N__5021),
            .I(D_LM_AMIGA_in_2));
    IoInMux I__668 (
            .O(N__5018),
            .I(N__5015));
    LocalMux I__667 (
            .O(N__5015),
            .I(N__5012));
    Sp12to4 I__666 (
            .O(N__5012),
            .I(N__5009));
    Span12Mux_s5_h I__665 (
            .O(N__5009),
            .I(N__5006));
    Span12Mux_h I__664 (
            .O(N__5006),
            .I(N__5003));
    Span12Mux_v I__663 (
            .O(N__5003),
            .I(N__5000));
    Odrv12 I__662 (
            .O(N__5000),
            .I(un2_D_LM_AMIGA_2));
    IoInMux I__661 (
            .O(N__4997),
            .I(N__4994));
    LocalMux I__660 (
            .O(N__4994),
            .I(N__4991));
    Span12Mux_s8_h I__659 (
            .O(N__4991),
            .I(N__4988));
    Odrv12 I__658 (
            .O(N__4988),
            .I(N_245_i));
    InMux I__657 (
            .O(N__4985),
            .I(N__4982));
    LocalMux I__656 (
            .O(N__4982),
            .I(N__4979));
    Span4Mux_v I__655 (
            .O(N__4979),
            .I(N__4976));
    Sp12to4 I__654 (
            .O(N__4976),
            .I(N__4973));
    Odrv12 I__653 (
            .O(N__4973),
            .I(D_LM_AMIGA_in_4));
    IoInMux I__652 (
            .O(N__4970),
            .I(N__4967));
    LocalMux I__651 (
            .O(N__4967),
            .I(N__4964));
    IoSpan4Mux I__650 (
            .O(N__4964),
            .I(N__4961));
    Sp12to4 I__649 (
            .O(N__4961),
            .I(N__4958));
    Span12Mux_s9_h I__648 (
            .O(N__4958),
            .I(N__4955));
    Span12Mux_h I__647 (
            .O(N__4955),
            .I(N__4952));
    Odrv12 I__646 (
            .O(N__4952),
            .I(un2_D_LM_AMIGA_4));
    InMux I__645 (
            .O(N__4949),
            .I(N__4946));
    LocalMux I__644 (
            .O(N__4946),
            .I(N__4943));
    Span4Mux_v I__643 (
            .O(N__4943),
            .I(N__4940));
    Span4Mux_h I__642 (
            .O(N__4940),
            .I(N__4937));
    Odrv4 I__641 (
            .O(N__4937),
            .I(WRITE_CYCLE_ACTIVE_rep16_i_ess));
    InMux I__640 (
            .O(N__4934),
            .I(N__4931));
    LocalMux I__639 (
            .O(N__4931),
            .I(WRITE_CYCLE_ACTIVE_rep20_i_ess));
    IoInMux I__638 (
            .O(N__4928),
            .I(N__4925));
    LocalMux I__637 (
            .O(N__4925),
            .I(N__4922));
    IoSpan4Mux I__636 (
            .O(N__4922),
            .I(N__4919));
    Span4Mux_s2_h I__635 (
            .O(N__4919),
            .I(N__4916));
    Span4Mux_h I__634 (
            .O(N__4916),
            .I(N__4913));
    Span4Mux_h I__633 (
            .O(N__4913),
            .I(N__4910));
    Odrv4 I__632 (
            .O(N__4910),
            .I(N_259_i));
    IoInMux I__631 (
            .O(N__4907),
            .I(N__4904));
    LocalMux I__630 (
            .O(N__4904),
            .I(N__4901));
    IoSpan4Mux I__629 (
            .O(N__4901),
            .I(N__4898));
    IoSpan4Mux I__628 (
            .O(N__4898),
            .I(N__4895));
    Span4Mux_s2_v I__627 (
            .O(N__4895),
            .I(N__4892));
    Span4Mux_v I__626 (
            .O(N__4892),
            .I(N__4889));
    Odrv4 I__625 (
            .O(N__4889),
            .I(N_240_i));
    IoInMux I__624 (
            .O(N__4886),
            .I(N__4883));
    LocalMux I__623 (
            .O(N__4883),
            .I(N__4880));
    Span12Mux_s7_v I__622 (
            .O(N__4880),
            .I(N__4877));
    Odrv12 I__621 (
            .O(N__4877),
            .I(N_243_i));
    IoInMux I__620 (
            .O(N__4874),
            .I(N__4871));
    LocalMux I__619 (
            .O(N__4871),
            .I(N__4868));
    Span4Mux_s2_h I__618 (
            .O(N__4868),
            .I(N__4865));
    Sp12to4 I__617 (
            .O(N__4865),
            .I(N__4862));
    Span12Mux_s9_v I__616 (
            .O(N__4862),
            .I(N__4859));
    Odrv12 I__615 (
            .O(N__4859),
            .I(N_263_i));
    IoInMux I__614 (
            .O(N__4856),
            .I(N__4853));
    LocalMux I__613 (
            .O(N__4853),
            .I(N__4850));
    Span4Mux_s2_h I__612 (
            .O(N__4850),
            .I(N__4847));
    Span4Mux_v I__611 (
            .O(N__4847),
            .I(N__4844));
    Span4Mux_v I__610 (
            .O(N__4844),
            .I(N__4841));
    Span4Mux_h I__609 (
            .O(N__4841),
            .I(N__4838));
    Odrv4 I__608 (
            .O(N__4838),
            .I(N_265_i));
    IoInMux I__607 (
            .O(N__4835),
            .I(N__4832));
    LocalMux I__606 (
            .O(N__4832),
            .I(N__4829));
    Span12Mux_s9_h I__605 (
            .O(N__4829),
            .I(N__4826));
    Odrv12 I__604 (
            .O(N__4826),
            .I(N_257_i));
    InMux I__603 (
            .O(N__4823),
            .I(N__4820));
    LocalMux I__602 (
            .O(N__4820),
            .I(N__4817));
    Span4Mux_v I__601 (
            .O(N__4817),
            .I(N__4814));
    Sp12to4 I__600 (
            .O(N__4814),
            .I(N__4811));
    Odrv12 I__599 (
            .O(N__4811),
            .I(D_LM_AMIGA_in_5));
    IoInMux I__598 (
            .O(N__4808),
            .I(N__4805));
    LocalMux I__597 (
            .O(N__4805),
            .I(N__4802));
    Span12Mux_s10_h I__596 (
            .O(N__4802),
            .I(N__4799));
    Span12Mux_h I__595 (
            .O(N__4799),
            .I(N__4796));
    Odrv12 I__594 (
            .O(N__4796),
            .I(un2_D_LM_AMIGA_5));
    IoInMux I__593 (
            .O(N__4793),
            .I(N__4790));
    LocalMux I__592 (
            .O(N__4790),
            .I(N__4787));
    Span12Mux_s10_v I__591 (
            .O(N__4787),
            .I(N__4784));
    Odrv12 I__590 (
            .O(N__4784),
            .I(N_250_i));
    InMux I__589 (
            .O(N__4781),
            .I(N__4778));
    LocalMux I__588 (
            .O(N__4778),
            .I(N__4775));
    Span4Mux_v I__587 (
            .O(N__4775),
            .I(N__4772));
    Span4Mux_h I__586 (
            .O(N__4772),
            .I(N__4769));
    Span4Mux_h I__585 (
            .O(N__4769),
            .I(N__4766));
    Odrv4 I__584 (
            .O(N__4766),
            .I(D_LM_AMIGA_in_7));
    IoInMux I__583 (
            .O(N__4763),
            .I(N__4760));
    LocalMux I__582 (
            .O(N__4760),
            .I(N__4757));
    IoSpan4Mux I__581 (
            .O(N__4757),
            .I(N__4754));
    Span4Mux_s3_h I__580 (
            .O(N__4754),
            .I(N__4751));
    Sp12to4 I__579 (
            .O(N__4751),
            .I(N__4748));
    Span12Mux_s11_h I__578 (
            .O(N__4748),
            .I(N__4745));
    Odrv12 I__577 (
            .O(N__4745),
            .I(un2_D_LM_AMIGA_7));
    IoInMux I__576 (
            .O(N__4742),
            .I(N__4739));
    LocalMux I__575 (
            .O(N__4739),
            .I(N__4736));
    IoSpan4Mux I__574 (
            .O(N__4736),
            .I(N__4733));
    Span4Mux_s3_h I__573 (
            .O(N__4733),
            .I(N__4730));
    Span4Mux_h I__572 (
            .O(N__4730),
            .I(N__4727));
    Odrv4 I__571 (
            .O(N__4727),
            .I(N_238_i));
    IoInMux I__570 (
            .O(N__4724),
            .I(N__4721));
    LocalMux I__569 (
            .O(N__4721),
            .I(N__4718));
    Span4Mux_s3_v I__568 (
            .O(N__4718),
            .I(N__4715));
    Span4Mux_v I__567 (
            .O(N__4715),
            .I(N__4712));
    Odrv4 I__566 (
            .O(N__4712),
            .I(N_241_i));
    IoInMux I__565 (
            .O(N__4709),
            .I(N__4706));
    LocalMux I__564 (
            .O(N__4706),
            .I(N__4703));
    Span12Mux_s10_h I__563 (
            .O(N__4703),
            .I(N__4700));
    Odrv12 I__562 (
            .O(N__4700),
            .I(N_261_i));
    IoInMux I__561 (
            .O(N__4697),
            .I(N__4694));
    LocalMux I__560 (
            .O(N__4694),
            .I(N__4691));
    IoSpan4Mux I__559 (
            .O(N__4691),
            .I(N__4688));
    Span4Mux_s1_h I__558 (
            .O(N__4688),
            .I(N__4685));
    Span4Mux_h I__557 (
            .O(N__4685),
            .I(N__4682));
    Odrv4 I__556 (
            .O(N__4682),
            .I(N_248_i));
    InMux I__555 (
            .O(N__4679),
            .I(N__4676));
    LocalMux I__554 (
            .O(N__4676),
            .I(N__4673));
    Span4Mux_v I__553 (
            .O(N__4673),
            .I(N__4670));
    Sp12to4 I__552 (
            .O(N__4670),
            .I(N__4667));
    Odrv12 I__551 (
            .O(N__4667),
            .I(D_LL_AMIGA_in_5));
    IoInMux I__550 (
            .O(N__4664),
            .I(N__4661));
    LocalMux I__549 (
            .O(N__4661),
            .I(N__4658));
    Span4Mux_s2_h I__548 (
            .O(N__4658),
            .I(N__4655));
    Span4Mux_v I__547 (
            .O(N__4655),
            .I(N__4652));
    Sp12to4 I__546 (
            .O(N__4652),
            .I(N__4649));
    Span12Mux_s11_h I__545 (
            .O(N__4649),
            .I(N__4646));
    Span12Mux_h I__544 (
            .O(N__4646),
            .I(N__4643));
    Odrv12 I__543 (
            .O(N__4643),
            .I(un2_D_LL_AMIGA_5));
    InMux I__542 (
            .O(N__4640),
            .I(N__4637));
    LocalMux I__541 (
            .O(N__4637),
            .I(N__4634));
    Span4Mux_h I__540 (
            .O(N__4634),
            .I(N__4631));
    Span4Mux_h I__539 (
            .O(N__4631),
            .I(N__4627));
    InMux I__538 (
            .O(N__4630),
            .I(N__4624));
    Sp12to4 I__537 (
            .O(N__4627),
            .I(N__4621));
    LocalMux I__536 (
            .O(N__4624),
            .I(N__4618));
    Span12Mux_v I__535 (
            .O(N__4621),
            .I(N__4613));
    Span12Mux_h I__534 (
            .O(N__4618),
            .I(N__4613));
    Odrv12 I__533 (
            .O(N__4613),
            .I(A_040_c_1));
    InMux I__532 (
            .O(N__4610),
            .I(N__4607));
    LocalMux I__531 (
            .O(N__4607),
            .I(N__4604));
    Span4Mux_v I__530 (
            .O(N__4604),
            .I(N__4601));
    Sp12to4 I__529 (
            .O(N__4601),
            .I(N__4598));
    Odrv12 I__528 (
            .O(N__4598),
            .I(D_LM_AMIGA_in_6));
    IoInMux I__527 (
            .O(N__4595),
            .I(N__4592));
    LocalMux I__526 (
            .O(N__4592),
            .I(N__4589));
    IoSpan4Mux I__525 (
            .O(N__4589),
            .I(N__4586));
    Span4Mux_s0_h I__524 (
            .O(N__4586),
            .I(N__4583));
    Sp12to4 I__523 (
            .O(N__4583),
            .I(N__4580));
    Span12Mux_h I__522 (
            .O(N__4580),
            .I(N__4577));
    Odrv12 I__521 (
            .O(N__4577),
            .I(un2_D_LM_AMIGA_6));
    IoInMux I__520 (
            .O(N__4574),
            .I(N__4571));
    LocalMux I__519 (
            .O(N__4571),
            .I(N__4568));
    IoSpan4Mux I__518 (
            .O(N__4568),
            .I(N__4565));
    IoSpan4Mux I__517 (
            .O(N__4565),
            .I(N__4562));
    Span4Mux_s3_h I__516 (
            .O(N__4562),
            .I(N__4559));
    Span4Mux_h I__515 (
            .O(N__4559),
            .I(N__4556));
    Odrv4 I__514 (
            .O(N__4556),
            .I(N_242_i));
    IoInMux I__513 (
            .O(N__4553),
            .I(N__4550));
    LocalMux I__512 (
            .O(N__4550),
            .I(N__4547));
    IoSpan4Mux I__511 (
            .O(N__4547),
            .I(N__4544));
    Span4Mux_s3_h I__510 (
            .O(N__4544),
            .I(N__4541));
    Span4Mux_h I__509 (
            .O(N__4541),
            .I(N__4538));
    Odrv4 I__508 (
            .O(N__4538),
            .I(N_260_i));
    InMux I__507 (
            .O(N__4535),
            .I(N__4532));
    LocalMux I__506 (
            .O(N__4532),
            .I(N__4528));
    IoInMux I__505 (
            .O(N__4531),
            .I(N__4525));
    Span4Mux_v I__504 (
            .O(N__4528),
            .I(N__4522));
    LocalMux I__503 (
            .O(N__4525),
            .I(N__4519));
    Sp12to4 I__502 (
            .O(N__4522),
            .I(N__4516));
    Span4Mux_s2_h I__501 (
            .O(N__4519),
            .I(N__4513));
    Span12Mux_h I__500 (
            .O(N__4516),
            .I(N__4510));
    Span4Mux_v I__499 (
            .O(N__4513),
            .I(N__4507));
    Span12Mux_h I__498 (
            .O(N__4510),
            .I(N__4504));
    Sp12to4 I__497 (
            .O(N__4507),
            .I(N__4501));
    Span12Mux_v I__496 (
            .O(N__4504),
            .I(N__4498));
    Span12Mux_s11_h I__495 (
            .O(N__4501),
            .I(N__4495));
    Span12Mux_v I__494 (
            .O(N__4498),
            .I(N__4492));
    Span12Mux_h I__493 (
            .O(N__4495),
            .I(N__4489));
    Odrv12 I__492 (
            .O(N__4492),
            .I(D_LL_040_in_3));
    Odrv12 I__491 (
            .O(N__4489),
            .I(D_LL_040_in_3));
    InMux I__490 (
            .O(N__4484),
            .I(N__4481));
    LocalMux I__489 (
            .O(N__4481),
            .I(N__4478));
    Span4Mux_v I__488 (
            .O(N__4478),
            .I(N__4475));
    Span4Mux_v I__487 (
            .O(N__4475),
            .I(N__4472));
    Sp12to4 I__486 (
            .O(N__4472),
            .I(N__4469));
    Span12Mux_h I__485 (
            .O(N__4469),
            .I(N__4466));
    Odrv12 I__484 (
            .O(N__4466),
            .I(D_UM_040_in_3));
    IoInMux I__483 (
            .O(N__4463),
            .I(N__4460));
    LocalMux I__482 (
            .O(N__4460),
            .I(N__4457));
    IoSpan4Mux I__481 (
            .O(N__4457),
            .I(N__4454));
    Span4Mux_s2_h I__480 (
            .O(N__4454),
            .I(N__4451));
    Span4Mux_h I__479 (
            .O(N__4451),
            .I(N__4448));
    Odrv4 I__478 (
            .O(N__4448),
            .I(un1_D_UM_040_3));
    IoInMux I__477 (
            .O(N__4445),
            .I(N__4442));
    LocalMux I__476 (
            .O(N__4442),
            .I(N__4439));
    Span4Mux_s3_v I__475 (
            .O(N__4439),
            .I(N__4436));
    Span4Mux_v I__474 (
            .O(N__4436),
            .I(N__4433));
    Odrv4 I__473 (
            .O(N__4433),
            .I(N_239_i));
    InMux I__472 (
            .O(N__4430),
            .I(N__4427));
    LocalMux I__471 (
            .O(N__4427),
            .I(N__4424));
    Span4Mux_v I__470 (
            .O(N__4424),
            .I(N__4421));
    Sp12to4 I__469 (
            .O(N__4421),
            .I(N__4418));
    Span12Mux_h I__468 (
            .O(N__4418),
            .I(N__4415));
    Span12Mux_h I__467 (
            .O(N__4415),
            .I(N__4412));
    Odrv12 I__466 (
            .O(N__4412),
            .I(D_UU_040_in_6));
    IoInMux I__465 (
            .O(N__4409),
            .I(N__4406));
    LocalMux I__464 (
            .O(N__4406),
            .I(N__4403));
    Span4Mux_s2_h I__463 (
            .O(N__4403),
            .I(N__4399));
    InMux I__462 (
            .O(N__4402),
            .I(N__4396));
    Span4Mux_v I__461 (
            .O(N__4399),
            .I(N__4393));
    LocalMux I__460 (
            .O(N__4396),
            .I(N__4390));
    Sp12to4 I__459 (
            .O(N__4393),
            .I(N__4387));
    Sp12to4 I__458 (
            .O(N__4390),
            .I(N__4384));
    Span12Mux_h I__457 (
            .O(N__4387),
            .I(N__4381));
    Span12Mux_s11_v I__456 (
            .O(N__4384),
            .I(N__4378));
    Span12Mux_h I__455 (
            .O(N__4381),
            .I(N__4375));
    Span12Mux_h I__454 (
            .O(N__4378),
            .I(N__4372));
    Odrv12 I__453 (
            .O(N__4375),
            .I(D_LM_040_in_6));
    Odrv12 I__452 (
            .O(N__4372),
            .I(D_LM_040_in_6));
    IoInMux I__451 (
            .O(N__4367),
            .I(N__4364));
    LocalMux I__450 (
            .O(N__4364),
            .I(N__4361));
    Span4Mux_s2_v I__449 (
            .O(N__4361),
            .I(N__4358));
    Span4Mux_h I__448 (
            .O(N__4358),
            .I(N__4355));
    Span4Mux_v I__447 (
            .O(N__4355),
            .I(N__4352));
    Odrv4 I__446 (
            .O(N__4352),
            .I(un1_D_UU_040_6));
    IoInMux I__445 (
            .O(N__4349),
            .I(N__4346));
    LocalMux I__444 (
            .O(N__4346),
            .I(N__4343));
    IoSpan4Mux I__443 (
            .O(N__4343),
            .I(N__4340));
    IoSpan4Mux I__442 (
            .O(N__4340),
            .I(N__4337));
    Span4Mux_s3_h I__441 (
            .O(N__4337),
            .I(N__4334));
    Odrv4 I__440 (
            .O(N__4334),
            .I(N_253_i));
    IoInMux I__439 (
            .O(N__4331),
            .I(N__4328));
    LocalMux I__438 (
            .O(N__4328),
            .I(N__4325));
    IoSpan4Mux I__437 (
            .O(N__4325),
            .I(N__4322));
    Span4Mux_s3_h I__436 (
            .O(N__4322),
            .I(N__4319));
    Span4Mux_v I__435 (
            .O(N__4319),
            .I(N__4316));
    Odrv4 I__434 (
            .O(N__4316),
            .I(N_254_i));
    IoInMux I__433 (
            .O(N__4313),
            .I(N__4310));
    LocalMux I__432 (
            .O(N__4310),
            .I(N__4307));
    IoSpan4Mux I__431 (
            .O(N__4307),
            .I(N__4304));
    Span4Mux_s3_h I__430 (
            .O(N__4304),
            .I(N__4301));
    Span4Mux_v I__429 (
            .O(N__4301),
            .I(N__4298));
    Odrv4 I__428 (
            .O(N__4298),
            .I(N_252_i));
    IoInMux I__427 (
            .O(N__4295),
            .I(N__4292));
    LocalMux I__426 (
            .O(N__4292),
            .I(N__4289));
    Odrv12 I__425 (
            .O(N__4289),
            .I(U111_CYCLE_SM_A_AMIGA_0_i_1));
    InMux I__424 (
            .O(N__4286),
            .I(N__4283));
    LocalMux I__423 (
            .O(N__4283),
            .I(N__4280));
    Span4Mux_h I__422 (
            .O(N__4280),
            .I(N__4277));
    Span4Mux_v I__421 (
            .O(N__4277),
            .I(N__4274));
    Odrv4 I__420 (
            .O(N__4274),
            .I(A_040_c_0));
    IoInMux I__419 (
            .O(N__4271),
            .I(N__4268));
    LocalMux I__418 (
            .O(N__4268),
            .I(N__4265));
    Span4Mux_s2_v I__417 (
            .O(N__4265),
            .I(N__4262));
    Span4Mux_v I__416 (
            .O(N__4262),
            .I(N__4259));
    Odrv4 I__415 (
            .O(N__4259),
            .I(A_AMIGA_c_0));
    IoInMux I__414 (
            .O(N__4256),
            .I(N__4253));
    LocalMux I__413 (
            .O(N__4253),
            .I(N__4250));
    Span4Mux_s2_h I__412 (
            .O(N__4250),
            .I(N__4247));
    Span4Mux_v I__411 (
            .O(N__4247),
            .I(N__4244));
    Span4Mux_h I__410 (
            .O(N__4244),
            .I(N__4241));
    Odrv4 I__409 (
            .O(N__4241),
            .I(N_264_i));
    IoInMux I__408 (
            .O(N__4238),
            .I(N__4235));
    LocalMux I__407 (
            .O(N__4235),
            .I(N__4232));
    IoSpan4Mux I__406 (
            .O(N__4232),
            .I(N__4229));
    IoSpan4Mux I__405 (
            .O(N__4229),
            .I(N__4226));
    Span4Mux_s2_h I__404 (
            .O(N__4226),
            .I(N__4223));
    Span4Mux_h I__403 (
            .O(N__4223),
            .I(N__4220));
    Odrv4 I__402 (
            .O(N__4220),
            .I(N_262_i));
    IoInMux I__401 (
            .O(N__4217),
            .I(N__4214));
    LocalMux I__400 (
            .O(N__4214),
            .I(N__4211));
    Span4Mux_s2_h I__399 (
            .O(N__4211),
            .I(N__4208));
    Span4Mux_h I__398 (
            .O(N__4208),
            .I(N__4205));
    Odrv4 I__397 (
            .O(N__4205),
            .I(N_258_i));
    IoInMux I__396 (
            .O(N__4202),
            .I(N__4199));
    LocalMux I__395 (
            .O(N__4199),
            .I(N__4196));
    IoSpan4Mux I__394 (
            .O(N__4196),
            .I(N__4193));
    Span4Mux_s3_h I__393 (
            .O(N__4193),
            .I(N__4190));
    Odrv4 I__392 (
            .O(N__4190),
            .I(N_246_i));
    IoInMux I__391 (
            .O(N__4187),
            .I(N__4184));
    LocalMux I__390 (
            .O(N__4184),
            .I(N__4181));
    Span4Mux_s0_v I__389 (
            .O(N__4181),
            .I(N__4178));
    Sp12to4 I__388 (
            .O(N__4178),
            .I(N__4175));
    Span12Mux_h I__387 (
            .O(N__4175),
            .I(N__4172));
    Span12Mux_v I__386 (
            .O(N__4172),
            .I(N__4169));
    Span12Mux_v I__385 (
            .O(N__4169),
            .I(N__4166));
    Odrv12 I__384 (
            .O(N__4166),
            .I(TAn_in));
    IoInMux I__383 (
            .O(N__4163),
            .I(N__4160));
    LocalMux I__382 (
            .O(N__4160),
            .I(N__4157));
    Span4Mux_s0_h I__381 (
            .O(N__4157),
            .I(N__4154));
    Span4Mux_h I__380 (
            .O(N__4154),
            .I(N__4151));
    Odrv4 I__379 (
            .O(N__4151),
            .I(N_267_i));
    IoInMux I__378 (
            .O(N__4148),
            .I(N__4145));
    LocalMux I__377 (
            .O(N__4145),
            .I(N__4142));
    Odrv12 I__376 (
            .O(N__4142),
            .I(RESETn_c_i));
    IoInMux I__375 (
            .O(N__4139),
            .I(N__4136));
    LocalMux I__374 (
            .O(N__4136),
            .I(N__4133));
    Span4Mux_s1_h I__373 (
            .O(N__4133),
            .I(N__4130));
    Span4Mux_v I__372 (
            .O(N__4130),
            .I(N__4127));
    Span4Mux_h I__371 (
            .O(N__4127),
            .I(N__4124));
    Odrv4 I__370 (
            .O(N__4124),
            .I(N_266_i));
    IoInMux I__369 (
            .O(N__4121),
            .I(N__4118));
    LocalMux I__368 (
            .O(N__4118),
            .I(N__4115));
    Odrv12 I__367 (
            .O(N__4115),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_0 ));
    IoInMux I__366 (
            .O(N__4112),
            .I(N__4109));
    LocalMux I__365 (
            .O(N__4109),
            .I(N__4106));
    Span4Mux_s3_h I__364 (
            .O(N__4106),
            .I(N__4103));
    Odrv4 I__363 (
            .O(N__4103),
            .I(N_247_i));
    IoInMux I__362 (
            .O(N__4100),
            .I(N__4097));
    LocalMux I__361 (
            .O(N__4097),
            .I(N__4094));
    IoSpan4Mux I__360 (
            .O(N__4094),
            .I(N__4091));
    Span4Mux_s0_h I__359 (
            .O(N__4091),
            .I(N__4088));
    Span4Mux_h I__358 (
            .O(N__4088),
            .I(N__4085));
    Odrv4 I__357 (
            .O(N__4085),
            .I(N_249_i));
    IoInMux I__356 (
            .O(N__4082),
            .I(N__4079));
    LocalMux I__355 (
            .O(N__4079),
            .I(N__4076));
    IoSpan4Mux I__354 (
            .O(N__4076),
            .I(N__4073));
    Span4Mux_s3_v I__353 (
            .O(N__4073),
            .I(N__4070));
    Span4Mux_v I__352 (
            .O(N__4070),
            .I(N__4067));
    Odrv4 I__351 (
            .O(N__4067),
            .I(N_251_i));
    IoInMux I__350 (
            .O(N__4064),
            .I(N__4061));
    LocalMux I__349 (
            .O(N__4061),
            .I(N__4058));
    Span4Mux_s0_h I__348 (
            .O(N__4058),
            .I(N__4055));
    Span4Mux_h I__347 (
            .O(N__4055),
            .I(N__4052));
    Span4Mux_h I__346 (
            .O(N__4052),
            .I(N__4049));
    Sp12to4 I__345 (
            .O(N__4049),
            .I(N__4046));
    Span12Mux_v I__344 (
            .O(N__4046),
            .I(N__4043));
    Span12Mux_v I__343 (
            .O(N__4043),
            .I(N__4040));
    Span12Mux_h I__342 (
            .O(N__4040),
            .I(N__4037));
    Odrv12 I__341 (
            .O(N__4037),
            .I(TCIn_c));
    INV \INVU111_CYCLE_SM.TSnC  (
            .O(\INVU111_CYCLE_SM.TSnC_net ),
            .I(N__9410));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__4148),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__4121),
            .GLOBALBUFFEROUTPUT(\U111_CYCLE_SM.CYCLE_STATE_0_g_0 ));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_6_LC_1_6_5.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_6_LC_1_6_5.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_6_LC_1_6_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_6_LC_1_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5786),
            .lcout(N_267_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_1_10_1.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_1_10_1.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_1_10_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_1_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6709),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_5_LC_1_11_1.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_5_LC_1_11_1.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_5_LC_1_11_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_5_LC_1_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5732),
            .lcout(N_266_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_LC_1_11_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_LC_1_11_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__9251),
            .in2(_gnd_net_),
            .in3(N__7094),
            .lcout(\U111_CYCLE_SM.CYCLE_STATE_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_2_LC_1_14_6.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_2_LC_1_14_6.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_2_LC_1_14_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_2_LC_1_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5621),
            .lcout(N_247_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_4_LC_1_16_7.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_4_LC_1_16_7.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_4_LC_1_16_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_4_LC_1_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5690),
            .lcout(N_249_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_6_LC_1_19_3.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_6_LC_1_19_3.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_6_LC_1_19_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_6_LC_1_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5771),
            .lcout(N_251_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_AMIGA_iobuf_RNO_0_LC_2_12_1.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_0_LC_2_12_1.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_0_LC_2_12_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_0_LC_2_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4949),
            .lcout(N_253_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_AMIGA_iobuf_RNO_1_LC_2_13_5.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_1_LC_2_13_5.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_1_LC_2_13_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_1_LC_2_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5462),
            .lcout(N_254_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_7_LC_2_15_0.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_7_LC_2_15_0.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_7_LC_2_15_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_7_LC_2_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6143),
            .lcout(N_252_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_1  (
            .in0(_gnd_net_),
            .in1(N__4630),
            .in2(_gnd_net_),
            .in3(N__6044),
            .lcout(U111_CYCLE_SM_A_AMIGA_0_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_2  (
            .in0(N__6043),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4286),
            .lcout(A_AMIGA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_3_LC_3_6_6.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_3_LC_3_6_6.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_3_LC_3_6_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_3_LC_3_6_6 (
            .in0(N__5411),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_264_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_1_LC_3_11_5.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_1_LC_3_11_5.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_1_LC_3_11_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_1_LC_3_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5426),
            .lcout(N_262_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_AMIGA_iobuf_RNO_5_LC_3_15_3.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_5_LC_3_15_3.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_5_LC_3_15_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_5_LC_3_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5567),
            .lcout(N_258_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_1_LC_3_15_5.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_1_LC_3_15_5.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_1_LC_3_15_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_1_LC_3_15_5 (
            .in0(N__6278),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_246_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_3_LC_3_18_1.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_3_LC_3_18_1.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_3_LC_3_18_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_3_LC_3_18_1 (
            .in0(N__6173),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_248_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_5_6_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_5_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_5_6_0  (
            .in0(N__11163),
            .in1(N__7409),
            .in2(_gnd_net_),
            .in3(N__4679),
            .lcout(un2_D_LL_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_5_11_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_5_11_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_5_11_2  (
            .in0(N__6465),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4640),
            .lcout(\U111_CYCLE_SM.N_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_5_16_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_5_16_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_5_16_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_5_16_7  (
            .in0(N__11118),
            .in1(N__8823),
            .in2(_gnd_net_),
            .in3(N__4610),
            .lcout(un2_D_LM_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_AMIGA_iobuf_RNO_5_LC_5_17_2.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_5_LC_5_17_2.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_5_LC_5_17_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_5_LC_5_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6158),
            .lcout(N_242_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_AMIGA_iobuf_RNO_7_LC_5_17_6.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_7_LC_5_17_6.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_7_LC_5_17_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_7_LC_5_17_6 (
            .in0(N__5744),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_260_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_5_18_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_5_18_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_5_18_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_5_18_1  (
            .in0(N__11139),
            .in1(N__4535),
            .in2(_gnd_net_),
            .in3(N__4484),
            .lcout(un1_D_UM_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_AMIGA_iobuf_RNO_2_LC_5_19_5.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_2_LC_5_19_5.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_2_LC_5_19_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_2_LC_5_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5552),
            .lcout(N_239_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_5_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_5_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_5_20_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_5_20_3  (
            .in0(N__4430),
            .in1(N__4402),
            .in2(_gnd_net_),
            .in3(N__11166),
            .lcout(un1_D_UU_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_2_LC_6_4_3.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_2_LC_6_4_3.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_2_LC_6_4_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_2_LC_6_4_3 (
            .in0(N__5609),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_263_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_4_LC_6_8_3.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_4_LC_6_8_3.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_4_LC_6_8_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_4_LC_6_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5654),
            .lcout(N_265_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_AMIGA_iobuf_RNO_4_LC_6_14_4.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_4_LC_6_14_4.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_4_LC_6_14_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_4_LC_6_14_4 (
            .in0(N__4934),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_257_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_6_14_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_6_14_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_6_14_7  (
            .in0(N__8352),
            .in1(N__4823),
            .in2(_gnd_net_),
            .in3(N__11086),
            .lcout(un2_D_LM_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_5_LC_6_16_1.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_5_LC_6_16_1.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_5_LC_6_16_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_5_LC_6_16_1 (
            .in0(N__6269),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_250_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_6_16_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_6_16_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_6_16_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_6_16_5  (
            .in0(N__4781),
            .in1(N__10471),
            .in2(_gnd_net_),
            .in3(N__11117),
            .lcout(un2_D_LM_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_AMIGA_iobuf_RNO_1_LC_6_18_5.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_1_LC_6_18_5.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_1_LC_6_18_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_1_LC_6_18_5 (
            .in0(N__5756),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_238_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_AMIGA_iobuf_RNO_4_LC_6_19_6.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_4_LC_6_19_6.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_4_LC_6_19_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_4_LC_6_19_6 (
            .in0(N__5702),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_241_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_0_LC_7_9_1.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_0_LC_7_9_1.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_0_LC_7_9_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_0_LC_7_9_1 (
            .in0(N__6056),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_261_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_AMIGA_iobuf_RNO_3_LC_7_11_1.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_3_LC_7_11_1.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_3_LC_7_11_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_3_LC_7_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5450),
            .lcout(N_256_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_7_12_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_7_12_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_7_12_4  (
            .in0(N__10971),
            .in1(N__7319),
            .in2(_gnd_net_),
            .in3(N__5027),
            .lcout(un2_D_LM_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_0_LC_7_12_6.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_0_LC_7_12_6.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_0_LC_7_12_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_0_LC_7_12_6 (
            .in0(N__5438),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_245_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_7_13_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_7_13_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_7_13_5  (
            .in0(N__11048),
            .in1(N__8452),
            .in2(_gnd_net_),
            .in3(N__4985),
            .lcout(un2_D_LM_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep16_i_ess_LC_7_14_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep16_i_ess_LC_7_14_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep16_i_ess_LC_7_14_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep16_i_ess_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(N__10077),
            .in2(_gnd_net_),
            .in3(N__9690),
            .lcout(WRITE_CYCLE_ACTIVE_rep16_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9409),
            .ce(N__9297),
            .sr(N__9225));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep20_i_ess_LC_7_14_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep20_i_ess_LC_7_14_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep20_i_ess_LC_7_14_4 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep20_i_ess_LC_7_14_4  (
            .in0(N__9691),
            .in1(_gnd_net_),
            .in2(N__10090),
            .in3(_gnd_net_),
            .lcout(WRITE_CYCLE_ACTIVE_rep20_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9409),
            .ce(N__9297),
            .sr(N__9225));
    defparam D_LM_AMIGA_iobuf_RNO_6_LC_7_16_1.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_6_LC_7_16_1.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_6_LC_7_16_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_6_LC_7_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5594),
            .lcout(N_259_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_AMIGA_iobuf_RNO_3_LC_7_18_1.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_3_LC_7_18_1.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_3_LC_7_18_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_3_LC_7_18_1 (
            .in0(N__5714),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_240_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_AMIGA_iobuf_RNO_6_LC_7_19_3.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_6_LC_7_19_3.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_6_LC_7_19_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_6_LC_7_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6260),
            .lcout(N_243_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_AMIGA_iobuf_RNO_0_LC_7_20_0.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_0_LC_7_20_0.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_0_LC_7_20_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_0_LC_7_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5582),
            .lcout(N_237_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_7_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_7_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_7_20_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_7_20_3  (
            .in0(N__5380),
            .in1(N__5330),
            .in2(_gnd_net_),
            .in3(N__11120),
            .lcout(un1_D_UU_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_7_20_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_7_20_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_7_20_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_7_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_8_6_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_8_6_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_8_6_0  (
            .in0(N__5261),
            .in1(N__9095),
            .in2(_gnd_net_),
            .in3(N__11130),
            .lcout(un2_D_LL_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_8_10_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_8_10_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_8_10_2  (
            .in0(N__7545),
            .in1(N__5228),
            .in2(_gnd_net_),
            .in3(N__11046),
            .lcout(un2_D_LM_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_8_10_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_8_10_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_8_10_4  (
            .in0(N__8761),
            .in1(N__5201),
            .in2(_gnd_net_),
            .in3(N__11047),
            .lcout(un2_D_LM_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam BUFENn_obuf_RNO_LC_8_19_3.C_ON=1'b0;
    defparam BUFENn_obuf_RNO_LC_8_19_3.SEQ_MODE=4'b0000;
    defparam BUFENn_obuf_RNO_LC_8_19_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 BUFENn_obuf_RNO_LC_8_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8051),
            .lcout(LBENn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_8_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_8_20_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_8_20_3  (
            .in0(N__5141),
            .in1(N__5096),
            .in2(_gnd_net_),
            .in3(N__11119),
            .lcout(un1_D_UU_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_9_7_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_9_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_9_7_6  (
            .in0(N__5057),
            .in1(N__8168),
            .in2(_gnd_net_),
            .in3(N__11076),
            .lcout(un2_D_LM_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_7_LC_9_10_3.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_7_LC_9_10_3.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_7_LC_9_10_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_7_LC_9_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5639),
            .lcout(N_268_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_AMIGA_iobuf_RNO_2_LC_9_12_5.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_2_LC_9_12_5.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_2_LC_9_12_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_2_LC_9_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5630),
            .lcout(N_255_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TSn_LC_9_12_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TSn_LC_9_12_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TSn_LC_9_12_7 .LUT_INIT=16'b0111011101010111;
    LogicCell40 \U111_CYCLE_SM.TSn_LC_9_12_7  (
            .in0(N__6742),
            .in1(N__6007),
            .in2(N__8050),
            .in3(N__6185),
            .lcout(TSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.TSnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep17_i_ess_LC_9_13_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep17_i_ess_LC_9_13_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep17_i_ess_LC_9_13_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep17_i_ess_LC_9_13_0  (
            .in0(N__9609),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10002),
            .lcout(WRITE_CYCLE_ACTIVE_rep17_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9404),
            .ce(N__9299),
            .sr(N__9227));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep19_i_ess_LC_9_13_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep19_i_ess_LC_9_13_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep19_i_ess_LC_9_13_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep19_i_ess_LC_9_13_1  (
            .in0(N__10003),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9610),
            .lcout(WRITE_CYCLE_ACTIVE_rep19_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9404),
            .ce(N__9299),
            .sr(N__9227));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep21_i_ess_LC_9_13_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep21_i_ess_LC_9_13_2 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep21_i_ess_LC_9_13_2 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep21_i_ess_LC_9_13_2  (
            .in0(N__9615),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10000),
            .lcout(READ_CYCLE_ACTIVE_rep21_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9404),
            .ce(N__9299),
            .sr(N__9227));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep8_i_ess_LC_9_13_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep8_i_ess_LC_9_13_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep8_i_ess_LC_9_13_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep8_i_ess_LC_9_13_3  (
            .in0(N__10007),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9614),
            .lcout(WRITE_CYCLE_ACTIVE_rep8_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9404),
            .ce(N__9299),
            .sr(N__9227));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep25_i_ess_LC_9_13_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep25_i_ess_LC_9_13_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep25_i_ess_LC_9_13_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep25_i_ess_LC_9_13_4  (
            .in0(N__9611),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10004),
            .lcout(WRITE_CYCLE_ACTIVE_rep25_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9404),
            .ce(N__9299),
            .sr(N__9227));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep27_i_ess_LC_9_13_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep27_i_ess_LC_9_13_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep27_i_ess_LC_9_13_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep27_i_ess_LC_9_13_5  (
            .in0(N__10005),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9612),
            .lcout(WRITE_CYCLE_ACTIVE_rep27_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9404),
            .ce(N__9299),
            .sr(N__9227));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep28_i_ess_LC_9_13_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep28_i_ess_LC_9_13_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep28_i_ess_LC_9_13_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep28_i_ess_LC_9_13_6  (
            .in0(N__9613),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10006),
            .lcout(WRITE_CYCLE_ACTIVE_rep28_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9404),
            .ce(N__9299),
            .sr(N__9227));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_i_ess_LC_9_13_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_i_ess_LC_9_13_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_i_ess_LC_9_13_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_i_ess_LC_9_13_7  (
            .in0(N__10001),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9608),
            .lcout(WRITE_CYCLE_ACTIVE_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9404),
            .ce(N__9299),
            .sr(N__9227));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep18_i_ess_LC_9_14_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep18_i_ess_LC_9_14_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep18_i_ess_LC_9_14_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep18_i_ess_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__9992),
            .in2(_gnd_net_),
            .in3(N__9571),
            .lcout(WRITE_CYCLE_ACTIVE_rep18_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9400),
            .ce(N__9301),
            .sr(N__9231));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep10_i_ess_LC_9_14_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep10_i_ess_LC_9_14_2 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep10_i_ess_LC_9_14_2 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep10_i_ess_LC_9_14_2  (
            .in0(N__9570),
            .in1(_gnd_net_),
            .in2(N__10047),
            .in3(_gnd_net_),
            .lcout(WRITE_CYCLE_ACTIVE_rep10_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9400),
            .ce(N__9301),
            .sr(N__9231));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep26_i_ess_LC_9_14_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep26_i_ess_LC_9_14_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep26_i_ess_LC_9_14_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep26_i_ess_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__9999),
            .in2(_gnd_net_),
            .in3(N__9574),
            .lcout(WRITE_CYCLE_ACTIVE_rep26_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9400),
            .ce(N__9301),
            .sr(N__9231));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep22_i_ess_LC_9_14_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep22_i_ess_LC_9_14_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep22_i_ess_LC_9_14_4 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep22_i_ess_LC_9_14_4  (
            .in0(N__9573),
            .in1(_gnd_net_),
            .in2(N__10049),
            .in3(_gnd_net_),
            .lcout(WRITE_CYCLE_ACTIVE_rep22_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9400),
            .ce(N__9301),
            .sr(N__9231));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep0_i_ess_LC_9_14_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep0_i_ess_LC_9_14_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep0_i_ess_LC_9_14_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep0_i_ess_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__9988),
            .in2(_gnd_net_),
            .in3(N__9569),
            .lcout(WRITE_CYCLE_ACTIVE_rep0_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9400),
            .ce(N__9301),
            .sr(N__9231));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep21_i_ess_LC_9_14_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep21_i_ess_LC_9_14_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep21_i_ess_LC_9_14_6 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep21_i_ess_LC_9_14_6  (
            .in0(N__9572),
            .in1(_gnd_net_),
            .in2(N__10048),
            .in3(_gnd_net_),
            .lcout(WRITE_CYCLE_ACTIVE_rep21_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9400),
            .ce(N__9301),
            .sr(N__9231));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep2_i_ess_LC_9_15_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep2_i_ess_LC_9_15_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep2_i_ess_LC_9_15_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep2_i_ess_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__9850),
            .in2(_gnd_net_),
            .in3(N__9620),
            .lcout(WRITE_CYCLE_ACTIVE_rep2_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9396),
            .ce(N__9302),
            .sr(N__9235));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep14_i_ess_LC_9_15_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep14_i_ess_LC_9_15_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep14_i_ess_LC_9_15_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep14_i_ess_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__9842),
            .in2(_gnd_net_),
            .in3(N__9616),
            .lcout(WRITE_CYCLE_ACTIVE_rep14_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9396),
            .ce(N__9302),
            .sr(N__9235));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep1_i_ess_LC_9_15_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep1_i_ess_LC_9_15_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep1_i_ess_LC_9_15_4 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep1_i_ess_LC_9_15_4  (
            .in0(N__9617),
            .in1(_gnd_net_),
            .in2(N__9899),
            .in3(_gnd_net_),
            .lcout(WRITE_CYCLE_ACTIVE_rep1_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9396),
            .ce(N__9302),
            .sr(N__9235));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep23_i_ess_LC_9_15_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep23_i_ess_LC_9_15_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep23_i_ess_LC_9_15_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep23_i_ess_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__9846),
            .in2(_gnd_net_),
            .in3(N__9618),
            .lcout(WRITE_CYCLE_ACTIVE_rep23_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9396),
            .ce(N__9302),
            .sr(N__9235));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep29_i_ess_LC_9_15_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep29_i_ess_LC_9_15_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep29_i_ess_LC_9_15_6 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep29_i_ess_LC_9_15_6  (
            .in0(N__9619),
            .in1(_gnd_net_),
            .in2(N__9900),
            .in3(_gnd_net_),
            .lcout(WRITE_CYCLE_ACTIVE_rep29_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9396),
            .ce(N__9302),
            .sr(N__9235));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep3_i_ess_LC_9_15_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep3_i_ess_LC_9_15_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep3_i_ess_LC_9_15_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep3_i_ess_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__9851),
            .in2(_gnd_net_),
            .in3(N__9621),
            .lcout(WRITE_CYCLE_ACTIVE_rep3_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9396),
            .ce(N__9302),
            .sr(N__9235));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep4_i_ess_LC_9_16_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep4_i_ess_LC_9_16_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep4_i_ess_LC_9_16_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep4_i_ess_LC_9_16_3  (
            .in0(N__9680),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10009),
            .lcout(WRITE_CYCLE_ACTIVE_rep4_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9391),
            .ce(N__9304),
            .sr(N__9238));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep7_i_ess_LC_9_16_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep7_i_ess_LC_9_16_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep7_i_ess_LC_9_16_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep7_i_ess_LC_9_16_6  (
            .in0(N__10010),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9681),
            .lcout(WRITE_CYCLE_ACTIVE_rep7_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9391),
            .ce(N__9304),
            .sr(N__9238));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep12_i_ess_LC_9_16_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep12_i_ess_LC_9_16_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep12_i_ess_LC_9_16_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep12_i_ess_LC_9_16_7  (
            .in0(N__9679),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10008),
            .lcout(WRITE_CYCLE_ACTIVE_rep12_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9391),
            .ce(N__9304),
            .sr(N__9238));
    defparam D_UU_AMIGA_iobuf_RNO_7_LC_9_17_2.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_7_LC_9_17_2.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_7_LC_9_17_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_7_LC_9_17_2 (
            .in0(N__5681),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_244_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_9_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_9_20_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_9_20_1  (
            .in0(N__5986),
            .in1(N__5951),
            .in2(_gnd_net_),
            .in3(N__11144),
            .lcout(un1_D_UU_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_9_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_9_20_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_9_20_7  (
            .in0(N__5902),
            .in1(N__5867),
            .in2(_gnd_net_),
            .in3(N__11143),
            .lcout(un1_D_UU_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_10_2_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_10_2_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_10_2_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_10_2_0  (
            .in0(N__5828),
            .in1(N__7485),
            .in2(_gnd_net_),
            .in3(N__11111),
            .lcout(un2_D_LL_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep18_i_ess_LC_10_6_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep18_i_ess_LC_10_6_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep18_i_ess_LC_10_6_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep18_i_ess_LC_10_6_0  (
            .in0(N__10084),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9717),
            .lcout(READ_CYCLE_ACTIVE_rep18_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9418),
            .ce(N__9307),
            .sr(N__9236));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep28_i_ess_LC_10_6_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep28_i_ess_LC_10_6_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep28_i_ess_LC_10_6_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep28_i_ess_LC_10_6_4  (
            .in0(N__10086),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9719),
            .lcout(READ_CYCLE_ACTIVE_rep28_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9418),
            .ce(N__9307),
            .sr(N__9236));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep26_i_ess_LC_10_6_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep26_i_ess_LC_10_6_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep26_i_ess_LC_10_6_5 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep26_i_ess_LC_10_6_5  (
            .in0(N__9718),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10085),
            .lcout(READ_CYCLE_ACTIVE_rep26_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9418),
            .ce(N__9307),
            .sr(N__9236));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep30_i_ess_LC_10_7_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep30_i_ess_LC_10_7_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep30_i_ess_LC_10_7_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep30_i_ess_LC_10_7_1  (
            .in0(N__10082),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9696),
            .lcout(READ_CYCLE_ACTIVE_rep30_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9417),
            .ce(N__9305),
            .sr(N__9232));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep27_i_ess_LC_10_7_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep27_i_ess_LC_10_7_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep27_i_ess_LC_10_7_6 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep27_i_ess_LC_10_7_6  (
            .in0(N__9695),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10081),
            .lcout(READ_CYCLE_ACTIVE_rep27_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9417),
            .ce(N__9305),
            .sr(N__9232));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep30_i_ess_LC_10_7_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep30_i_ess_LC_10_7_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep30_i_ess_LC_10_7_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep30_i_ess_LC_10_7_7  (
            .in0(N__10083),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9694),
            .lcout(WRITE_CYCLE_ACTIVE_rep30_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9417),
            .ce(N__9305),
            .sr(N__9232));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep17_i_ess_LC_10_8_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep17_i_ess_LC_10_8_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep17_i_ess_LC_10_8_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep17_i_ess_LC_10_8_3  (
            .in0(_gnd_net_),
            .in1(N__10058),
            .in2(_gnd_net_),
            .in3(N__9697),
            .lcout(READ_CYCLE_ACTIVE_rep17_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9416),
            .ce(N__9303),
            .sr(N__9228));
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_10_9_0.C_ON=1'b0;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_10_9_0.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_10_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK40_THRU_LUT4_0_LC_10_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9422),
            .lcout(GB_BUFFER_CLK40_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep25_i_ess_LC_10_10_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep25_i_ess_LC_10_10_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep25_i_ess_LC_10_10_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep25_i_ess_LC_10_10_7  (
            .in0(_gnd_net_),
            .in1(N__10057),
            .in2(_gnd_net_),
            .in3(N__9709),
            .lcout(READ_CYCLE_ACTIVE_rep25_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9412),
            .ce(N__9300),
            .sr(N__9224));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep14_i_ess_LC_10_11_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep14_i_ess_LC_10_11_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep14_i_ess_LC_10_11_1 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep14_i_ess_LC_10_11_1  (
            .in0(N__9693),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10050),
            .lcout(READ_CYCLE_ACTIVE_rep14_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9411),
            .ce(N__9296),
            .sr(N__9226));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep24_i_ess_LC_10_11_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep24_i_ess_LC_10_11_2 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep24_i_ess_LC_10_11_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep24_i_ess_LC_10_11_2  (
            .in0(N__10051),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9692),
            .lcout(WRITE_CYCLE_ACTIVE_rep24_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9411),
            .ce(N__9296),
            .sr(N__9226));
    defparam \U111_CYCLE_SM.A2_EN_LC_10_12_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A2_EN_LC_10_12_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.A2_EN_LC_10_12_1 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \U111_CYCLE_SM.A2_EN_LC_10_12_1  (
            .in0(N__6034),
            .in1(N__6224),
            .in2(_gnd_net_),
            .in3(N__6941),
            .lcout(\U111_CYCLE_SM.A2_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9405),
            .ce(),
            .sr(N__9229));
    defparam \U111_CYCLE_SM.TA_DIS_LC_10_12_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TA_DIS_LC_10_12_3 .LUT_INIT=16'b0011001101110010;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_LC_10_12_3  (
            .in0(N__6436),
            .in1(N__6236),
            .in2(N__8068),
            .in3(N__6943),
            .lcout(\U111_CYCLE_SM.TA_DISZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9405),
            .ce(),
            .sr(N__9229));
    defparam \U111_CYCLE_SM.FLIP_WORD_LC_10_12_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_LC_10_12_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.FLIP_WORD_LC_10_12_4 .LUT_INIT=16'b1100110011111010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_LC_10_12_4  (
            .in0(N__6942),
            .in1(N__6023),
            .in2(N__10970),
            .in3(N__6435),
            .lcout(\U111_CYCLE_SM.FLIP_WORDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9405),
            .ce(),
            .sr(N__9229));
    defparam \U111_CYCLE_SM.LATCH_EN_LC_10_12_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LATCH_EN_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LATCH_EN_LC_10_12_5 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \U111_CYCLE_SM.LATCH_EN_LC_10_12_5  (
            .in0(N__6368),
            .in1(N__6940),
            .in2(N__10326),
            .in3(N__6359),
            .lcout(\U111_CYCLE_SM.LATCH_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9405),
            .ce(),
            .sr(N__9229));
    defparam \U111_CYCLE_SM.TS_EN_LC_10_12_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_LC_10_12_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TS_EN_LC_10_12_6 .LUT_INIT=16'b0000010000001110;
    LogicCell40 \U111_CYCLE_SM.TS_EN_LC_10_12_6  (
            .in0(N__6230),
            .in1(N__6008),
            .in2(N__6917),
            .in3(N__7250),
            .lcout(\U111_CYCLE_SM.TS_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9405),
            .ce(),
            .sr(N__9229));
    defparam \U111_CYCLE_SM.TS_DELAY_LC_10_13_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_DELAY_LC_10_13_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.TS_DELAY_LC_10_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.TS_DELAY_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6218),
            .lcout(\U111_CYCLE_SM.TS_DELAYZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9401),
            .ce(),
            .sr(N__9233));
    defparam \U111_CYCLE_SM.TS_DELAY_RNI91BJ_LC_10_14_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_DELAY_RNI91BJ_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_DELAY_RNI91BJ_LC_10_14_4 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \U111_CYCLE_SM.TS_DELAY_RNI91BJ_LC_10_14_4  (
            .in0(N__6203),
            .in1(N__8049),
            .in2(_gnd_net_),
            .in3(N__6184),
            .lcout(\U111_CYCLE_SM.N_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep6_i_ess_LC_10_15_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep6_i_ess_LC_10_15_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep6_i_ess_LC_10_15_0 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep6_i_ess_LC_10_15_0  (
            .in0(N__9582),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9837),
            .lcout(READ_CYCLE_ACTIVE_rep6_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9392),
            .ce(N__9306),
            .sr(N__9239));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep11_i_ess_LC_10_15_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep11_i_ess_LC_10_15_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep11_i_ess_LC_10_15_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep11_i_ess_LC_10_15_1  (
            .in0(N__9838),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9575),
            .lcout(WRITE_CYCLE_ACTIVE_rep11_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9392),
            .ce(N__9306),
            .sr(N__9239));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep23_i_ess_LC_10_15_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep23_i_ess_LC_10_15_2 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep23_i_ess_LC_10_15_2 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep23_i_ess_LC_10_15_2  (
            .in0(N__9580),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9835),
            .lcout(READ_CYCLE_ACTIVE_rep23_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9392),
            .ce(N__9306),
            .sr(N__9239));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep13_i_ess_LC_10_15_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep13_i_ess_LC_10_15_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep13_i_ess_LC_10_15_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep13_i_ess_LC_10_15_3  (
            .in0(N__9834),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9579),
            .lcout(READ_CYCLE_ACTIVE_rep13_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9392),
            .ce(N__9306),
            .sr(N__9239));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep5_i_ess_LC_10_15_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep5_i_ess_LC_10_15_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep5_i_ess_LC_10_15_4 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep5_i_ess_LC_10_15_4  (
            .in0(N__9581),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9836),
            .lcout(READ_CYCLE_ACTIVE_rep5_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9392),
            .ce(N__9306),
            .sr(N__9239));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep5_i_ess_LC_10_15_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep5_i_ess_LC_10_15_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep5_i_ess_LC_10_15_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep5_i_ess_LC_10_15_5  (
            .in0(N__9840),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9577),
            .lcout(WRITE_CYCLE_ACTIVE_rep5_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9392),
            .ce(N__9306),
            .sr(N__9239));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep15_i_ess_LC_10_15_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep15_i_ess_LC_10_15_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep15_i_ess_LC_10_15_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep15_i_ess_LC_10_15_6  (
            .in0(N__9576),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9839),
            .lcout(WRITE_CYCLE_ACTIVE_rep15_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9392),
            .ce(N__9306),
            .sr(N__9239));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep9_i_ess_LC_10_15_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep9_i_ess_LC_10_15_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep9_i_ess_LC_10_15_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep9_i_ess_LC_10_15_7  (
            .in0(N__9841),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9578),
            .lcout(WRITE_CYCLE_ACTIVE_rep9_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9392),
            .ce(N__9306),
            .sr(N__9239));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep13_i_ess_LC_10_16_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep13_i_ess_LC_10_16_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep13_i_ess_LC_10_16_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep13_i_ess_LC_10_16_4  (
            .in0(_gnd_net_),
            .in1(N__10040),
            .in2(_gnd_net_),
            .in3(N__9674),
            .lcout(WRITE_CYCLE_ACTIVE_rep13_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9388),
            .ce(N__9308),
            .sr(N__9241));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep6_i_ess_LC_10_16_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep6_i_ess_LC_10_16_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep6_i_ess_LC_10_16_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep6_i_ess_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(N__10041),
            .in2(_gnd_net_),
            .in3(N__9675),
            .lcout(WRITE_CYCLE_ACTIVE_rep6_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9388),
            .ce(N__9308),
            .sr(N__9241));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep7_i_ess_LC_10_17_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep7_i_ess_LC_10_17_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep7_i_ess_LC_10_17_0 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep7_i_ess_LC_10_17_0  (
            .in0(N__9683),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10043),
            .lcout(READ_CYCLE_ACTIVE_rep7_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9385),
            .ce(N__9310),
            .sr(N__9243));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep2_i_ess_LC_10_17_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep2_i_ess_LC_10_17_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep2_i_ess_LC_10_17_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep2_i_ess_LC_10_17_3  (
            .in0(N__10042),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9682),
            .lcout(READ_CYCLE_ACTIVE_rep2_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9385),
            .ce(N__9310),
            .sr(N__9243));
    defparam LBENn_c_sbtinv_LC_11_1_6.C_ON=1'b0;
    defparam LBENn_c_sbtinv_LC_11_1_6.SEQ_MODE=4'b0000;
    defparam LBENn_c_sbtinv_LC_11_1_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 LBENn_c_sbtinv_LC_11_1_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8015),
            .lcout(LBENn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep24_i_ess_LC_11_11_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep24_i_ess_LC_11_11_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep24_i_ess_LC_11_11_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep24_i_ess_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__10014),
            .in2(_gnd_net_),
            .in3(N__9707),
            .lcout(READ_CYCLE_ACTIVE_rep24_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9406),
            .ce(N__9298),
            .sr(N__9230));
    defparam \U111_CYCLE_SM.TA_DIS_RNO_0_LC_11_12_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_RNO_0_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_DIS_RNO_0_LC_11_12_0 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_RNO_0_LC_11_12_0  (
            .in0(N__6481),
            .in1(N__6498),
            .in2(_gnd_net_),
            .in3(N__6432),
            .lcout(\U111_CYCLE_SM.N_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_12_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_12_2 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_12_2  (
            .in0(N__6773),
            .in1(N__6836),
            .in2(N__7155),
            .in3(N__6939),
            .lcout(\U111_CYCLE_SM.N_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_11_12_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_11_12_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_11_12_3  (
            .in0(N__6835),
            .in1(N__7146),
            .in2(_gnd_net_),
            .in3(N__6772),
            .lcout(\U111_CYCLE_SM.N_75 ),
            .ltout(\U111_CYCLE_SM.N_75_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_11_12_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_11_12_4 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_1_LC_11_12_4  (
            .in0(N__6743),
            .in1(N__6358),
            .in2(N__6371),
            .in3(N__7037),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9402),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_3_LC_11_12_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_3_LC_11_12_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_3_LC_11_12_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_3_LC_11_12_5  (
            .in0(N__6893),
            .in1(N__6744),
            .in2(_gnd_net_),
            .in3(N__7234),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9402),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LATCH_EN_RNO_0_LC_11_12_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LATCH_EN_RNO_0_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LATCH_EN_RNO_0_LC_11_12_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U111_CYCLE_SM.LATCH_EN_RNO_0_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(N__6875),
            .in2(_gnd_net_),
            .in3(N__7081),
            .lcout(\U111_CYCLE_SM.LATCH_EN_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.BURST_LC_11_13_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_LC_11_13_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.BURST_LC_11_13_0 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U111_CYCLE_SM.BURST_LC_11_13_0  (
            .in0(N__6334),
            .in1(N__6356),
            .in2(N__6310),
            .in3(N__7036),
            .lcout(\U111_CYCLE_SM.BURSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9397),
            .ce(),
            .sr(N__9237));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI541Q_0_LC_11_13_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI541Q_0_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI541Q_0_LC_11_13_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNI541Q_0_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(N__7082),
            .in2(_gnd_net_),
            .in3(N__9567),
            .lcout(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ),
            .ltout(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.BURST_COUNT_0_LC_11_13_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_COUNT_0_LC_11_13_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.BURST_COUNT_0_LC_11_13_2 .LUT_INIT=16'b0000110000000011;
    LogicCell40 \U111_CYCLE_SM.BURST_COUNT_0_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__6891),
            .in2(N__6362),
            .in3(N__6976),
            .lcout(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9397),
            .ce(),
            .sr(N__9237));
    defparam \U111_CYCLE_SM.BURST_COUNT_1_LC_11_13_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_COUNT_1_LC_11_13_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.BURST_COUNT_1_LC_11_13_6 .LUT_INIT=16'b0010001000010010;
    LogicCell40 \U111_CYCLE_SM.BURST_COUNT_1_LC_11_13_6  (
            .in0(N__7052),
            .in1(N__6355),
            .in2(N__6980),
            .in3(N__6892),
            .lcout(\U111_CYCLE_SM.BURST_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9397),
            .ce(),
            .sr(N__9237));
    defparam \U111_CYCLE_SM.LW_TRANS_LC_11_13_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_TRANS_LC_11_13_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LW_TRANS_LC_11_13_7 .LUT_INIT=16'b1101011110000010;
    LogicCell40 \U111_CYCLE_SM.LW_TRANS_LC_11_13_7  (
            .in0(N__6357),
            .in1(N__6335),
            .in2(N__6311),
            .in3(N__6499),
            .lcout(\U111_CYCLE_SM.LW_TRANSZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9397),
            .ce(),
            .sr(N__9237));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_11_14_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_11_14_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_11_14_0 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_11_14_0  (
            .in0(N__6874),
            .in1(N__7084),
            .in2(N__10073),
            .in3(N__9568),
            .lcout(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9393),
            .ce(),
            .sr(N__9240));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep0_i_ess_LC_11_15_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep0_i_ess_LC_11_15_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep0_i_ess_LC_11_15_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep0_i_ess_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__9819),
            .in2(_gnd_net_),
            .in3(N__9642),
            .lcout(READ_CYCLE_ACTIVE_rep0_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9389),
            .ce(N__9309),
            .sr(N__9242));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep9_i_ess_LC_11_15_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep9_i_ess_LC_11_15_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep9_i_ess_LC_11_15_1 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep9_i_ess_LC_11_15_1  (
            .in0(N__9648),
            .in1(_gnd_net_),
            .in2(N__9898),
            .in3(_gnd_net_),
            .lcout(READ_CYCLE_ACTIVE_rep9_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9389),
            .ce(N__9309),
            .sr(N__9242));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep15_i_ess_LC_11_15_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep15_i_ess_LC_11_15_2 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep15_i_ess_LC_11_15_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep15_i_ess_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__9823),
            .in2(_gnd_net_),
            .in3(N__9644),
            .lcout(READ_CYCLE_ACTIVE_rep15_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9389),
            .ce(N__9309),
            .sr(N__9242));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep1_i_ess_LC_11_15_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep1_i_ess_LC_11_15_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep1_i_ess_LC_11_15_3 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep1_i_ess_LC_11_15_3  (
            .in0(N__9645),
            .in1(_gnd_net_),
            .in2(N__9896),
            .in3(_gnd_net_),
            .lcout(READ_CYCLE_ACTIVE_rep1_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9389),
            .ce(N__9309),
            .sr(N__9242));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep3_i_ess_LC_11_15_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep3_i_ess_LC_11_15_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep3_i_ess_LC_11_15_5 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep3_i_ess_LC_11_15_5  (
            .in0(N__9646),
            .in1(_gnd_net_),
            .in2(N__9897),
            .in3(_gnd_net_),
            .lcout(READ_CYCLE_ACTIVE_rep3_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9389),
            .ce(N__9309),
            .sr(N__9242));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep8_i_ess_LC_11_15_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep8_i_ess_LC_11_15_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep8_i_ess_LC_11_15_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep8_i_ess_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__9830),
            .in2(_gnd_net_),
            .in3(N__9647),
            .lcout(READ_CYCLE_ACTIVE_rep8_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9389),
            .ce(N__9309),
            .sr(N__9242));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep11_i_ess_LC_11_15_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep11_i_ess_LC_11_15_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep11_i_ess_LC_11_15_7 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep11_i_ess_LC_11_15_7  (
            .in0(N__9643),
            .in1(_gnd_net_),
            .in2(N__9895),
            .in3(_gnd_net_),
            .lcout(READ_CYCLE_ACTIVE_rep11_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9389),
            .ce(N__9309),
            .sr(N__9242));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep4_i_ess_LC_11_16_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep4_i_ess_LC_11_16_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep4_i_ess_LC_11_16_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep4_i_ess_LC_11_16_7  (
            .in0(N__10038),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9698),
            .lcout(READ_CYCLE_ACTIVE_rep4_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9386),
            .ce(N__9311),
            .sr(N__9244));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep12_i_ess_LC_11_17_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep12_i_ess_LC_11_17_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep12_i_ess_LC_11_17_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep12_i_ess_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__10039),
            .in2(_gnd_net_),
            .in3(N__9699),
            .lcout(READ_CYCLE_ACTIVE_rep12_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9384),
            .ce(N__9312),
            .sr(N__9245));
    defparam D_UU_040_iobuf_RNO_6_LC_11_18_3.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_6_LC_11_18_3.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_6_LC_11_18_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_040_iobuf_RNO_6_LC_11_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6404),
            .lcout(N_211_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_040_iobuf_RNO_2_LC_11_20_2.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_2_LC_11_20_2.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_2_LC_11_20_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_040_iobuf_RNO_2_LC_11_20_2 (
            .in0(N__6674),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_207_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_12_2_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_12_2_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_12_2_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_12_2_1  (
            .in0(N__9158),
            .in1(N__6650),
            .in2(_gnd_net_),
            .in3(N__11162),
            .lcout(un2_D_LL_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_12_3_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_12_3_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_12_3_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_12_3_3  (
            .in0(N__6611),
            .in1(N__8279),
            .in2(_gnd_net_),
            .in3(N__11161),
            .lcout(un2_D_LL_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_2_LC_12_3_6.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_2_LC_12_3_6.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_2_LC_12_3_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_040_iobuf_RNO_2_LC_12_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6569),
            .lcout(N_231_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_12_7_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_12_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_12_7_7  (
            .in0(N__6542),
            .in1(N__8687),
            .in2(_gnd_net_),
            .in3(N__11122),
            .lcout(un2_D_LL_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.PORT_MISMATCH_LC_12_9_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.PORT_MISMATCH_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.PORT_MISMATCH_LC_12_9_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \U111_CYCLE_SM.PORT_MISMATCH_LC_12_9_3  (
            .in0(N__7232),
            .in1(N__6506),
            .in2(N__6482),
            .in3(N__6440),
            .lcout(\U111_CYCLE_SM.PORT_MISMATCHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9408),
            .ce(),
            .sr(N__9234));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_2_LC_12_12_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_2_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_2_LC_12_12_0 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_1_2_LC_12_12_0  (
            .in0(N__6433),
            .in1(N__7233),
            .in2(N__7197),
            .in3(N__6959),
            .lcout(),
            .ltout(\U111_CYCLE_SM.N_60_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_2_LC_12_12_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_2_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_2_LC_12_12_1 .LUT_INIT=16'b0000100000001010;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_2_LC_12_12_1  (
            .in0(N__6745),
            .in1(N__6434),
            .in2(N__6407),
            .in3(N__6899),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9395),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_12_12_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_12_12_3 .LUT_INIT=16'b0101111101011111;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_12_12_3  (
            .in0(N__6770),
            .in1(_gnd_net_),
            .in2(N__6847),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\U111_CYCLE_SM.N_46_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_5_LC_12_12_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_5_LC_12_12_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_5_LC_12_12_4 .LUT_INIT=16'b1100110000001000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_5_LC_12_12_4  (
            .in0(N__7184),
            .in1(N__6747),
            .in2(N__6947),
            .in3(N__6913),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9395),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_12_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_12_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_12_5  (
            .in0(N__6746),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6944),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9395),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.BURST_RNILNBJ_LC_12_12_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_RNILNBJ_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.BURST_RNILNBJ_LC_12_12_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U111_CYCLE_SM.BURST_RNILNBJ_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(N__6769),
            .in2(_gnd_net_),
            .in3(N__7035),
            .lcout(\U111_CYCLE_SM.N_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_12_12_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_12_12_7 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_12_12_7  (
            .in0(N__6837),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7126),
            .lcout(\U111_CYCLE_SM.N_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_13_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_13_0 .LUT_INIT=16'b1111111100111111;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__6842),
            .in2(N__7127),
            .in3(N__7189),
            .lcout(\U111_CYCLE_SM.N_40 ),
            .ltout(\U111_CYCLE_SM.N_40_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTO81_LC_12_13_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTO81_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTO81_LC_12_13_1 .LUT_INIT=16'b0101010101011111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTO81_LC_12_13_1  (
            .in0(N__6749),
            .in1(_gnd_net_),
            .in2(N__6878),
            .in3(N__6870),
            .lcout(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81 ),
            .ltout(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI0BVS1_2_LC_12_13_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI0BVS1_2_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI0BVS1_2_LC_12_13_2 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNI0BVS1_2_LC_12_13_2  (
            .in0(N__7125),
            .in1(N__6841),
            .in2(N__6854),
            .in3(N__7188),
            .lcout(\U111_CYCLE_SM.N_40_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_12_13_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_12_13_3 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_12_13_3  (
            .in0(N__6843),
            .in1(N__6771),
            .in2(_gnd_net_),
            .in3(N__7123),
            .lcout(),
            .ltout(\U111_CYCLE_SM.N_55_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_13_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_13_4 .LUT_INIT=16'b1111011111110011;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_13_4  (
            .in0(N__7193),
            .in1(N__6748),
            .in2(N__7253),
            .in3(N__7246),
            .lcout(\U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_13_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_13_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_13_5  (
            .in0(N__7235),
            .in1(N__6958),
            .in2(N__7198),
            .in3(N__7124),
            .lcout(),
            .ltout(\U111_CYCLE_SM.N_57_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_13_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_13_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_13_6  (
            .in0(N__7083),
            .in1(N__9708),
            .in2(N__7103),
            .in3(N__7100),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9390),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_12_13_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_12_13_7 .LUT_INIT=16'b1011111100111111;
    LogicCell40 \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_12_13_7  (
            .in0(N__7051),
            .in1(N__7034),
            .in2(N__7013),
            .in3(N__6975),
            .lcout(\U111_CYCLE_SM.N_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_12_14_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_12_14_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_12_14_0  (
            .in0(N__7547),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9387),
            .ce(N__8234),
            .sr(N__8201));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_12_14_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_12_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_12_14_1  (
            .in0(N__8682),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9387),
            .ce(N__8234),
            .sr(N__8201));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_12_14_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_12_14_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_12_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7408),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9387),
            .ce(N__8234),
            .sr(N__8201));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_12_14_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_12_14_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_12_14_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_12_14_3  (
            .in0(N__7318),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9387),
            .ce(N__8234),
            .sr(N__8201));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_12_14_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_12_14_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_12_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7490),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9387),
            .ce(N__8234),
            .sr(N__8201));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_12_14_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_12_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8528),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9387),
            .ce(N__8234),
            .sr(N__8201));
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_15_4.C_ON=1'b0;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_15_4.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_15_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_15_4 (
            .in0(N__7715),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_CLK80_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_040_iobuf_RNO_5_LC_12_15_5.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_5_LC_12_15_5.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_5_LC_12_15_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_040_iobuf_RNO_5_LC_12_15_5 (
            .in0(N__7664),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_210_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_12_15_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_12_15_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_12_15_6  (
            .in0(N__7634),
            .in1(N__7606),
            .in2(_gnd_net_),
            .in3(N__11061),
            .lcout(un1_D_UM_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_12_16_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_12_16_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_12_16_2  (
            .in0(N__10367),
            .in1(N__7556),
            .in2(_gnd_net_),
            .in3(N__7546),
            .lcout(un1_D_UU_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_12_17_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_12_17_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_12_17_3  (
            .in0(N__7486),
            .in1(N__7442),
            .in2(_gnd_net_),
            .in3(N__10393),
            .lcout(un1_D_UM_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_12_18_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_12_18_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_12_18_2  (
            .in0(N__7401),
            .in1(N__7364),
            .in2(_gnd_net_),
            .in3(N__10394),
            .lcout(un1_D_UM_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_12_18_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_12_18_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_12_18_6  (
            .in0(N__7328),
            .in1(N__7317),
            .in2(_gnd_net_),
            .in3(N__10395),
            .lcout(un1_D_UU_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_040_iobuf_RNO_1_LC_12_18_7.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_1_LC_12_18_7.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_1_LC_12_18_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_040_iobuf_RNO_1_LC_12_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7262),
            .lcout(N_206_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_12_19_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_12_19_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_12_19_5  (
            .in0(N__8075),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8033),
            .lcout(TAn_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_12_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_12_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_12_20_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_12_20_7  (
            .in0(N__7957),
            .in1(N__7931),
            .in2(_gnd_net_),
            .in3(N__11121),
            .lcout(un1_D_UU_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_13_3_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_13_3_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_13_3_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_13_3_1  (
            .in0(N__11164),
            .in1(N__9029),
            .in2(_gnd_net_),
            .in3(N__7895),
            .lcout(un2_D_LL_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_13_3_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_13_3_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_13_3_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_13_3_6  (
            .in0(N__8527),
            .in1(N__7856),
            .in2(_gnd_net_),
            .in3(N__11165),
            .lcout(un2_D_LL_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_13_9_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_13_9_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_13_9_1  (
            .in0(N__7813),
            .in1(N__7772),
            .in2(_gnd_net_),
            .in3(N__11093),
            .lcout(un1_D_UM_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_11_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_11_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_11_1  (
            .in0(N__8243),
            .in1(N__8272),
            .in2(_gnd_net_),
            .in3(N__10350),
            .lcout(un1_D_UM_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_13_12_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_13_12_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_13_12_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_13_12_0  (
            .in0(N__8765),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9403),
            .ce(N__8236),
            .sr(N__8212));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_13_12_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_13_12_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_13_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9144),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9403),
            .ce(N__8236),
            .sr(N__8212));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_13_12_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_13_12_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_13_12_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_13_12_6  (
            .in0(N__8271),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9403),
            .ce(N__8236),
            .sr(N__8212));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_13_13_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_13_13_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_13_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9090),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9398),
            .ce(N__8235),
            .sr(N__8211));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_13_14_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_13_14_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_13_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_13_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8372),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9394),
            .ce(N__8237),
            .sr(N__8213));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_13_14_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_13_14_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_13_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8456),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9394),
            .ce(N__8237),
            .sr(N__8213));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_13_14_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_13_14_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_13_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_13_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8164),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9394),
            .ce(N__8237),
            .sr(N__8213));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_13_14_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_13_14_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_13_14_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_13_14_5  (
            .in0(N__8825),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9394),
            .ce(N__8237),
            .sr(N__8213));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_13_14_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_13_14_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_13_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_13_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9024),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9394),
            .ce(N__8237),
            .sr(N__8213));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_13_14_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_13_14_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_13_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_13_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10472),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9394),
            .ce(N__8237),
            .sr(N__8213));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_13_15_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_13_15_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_13_15_1  (
            .in0(N__8163),
            .in1(N__8123),
            .in2(_gnd_net_),
            .in3(N__10380),
            .lcout(un1_D_UU_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_13_18_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_13_18_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_13_18_4  (
            .in0(N__10403),
            .in1(N__8834),
            .in2(_gnd_net_),
            .in3(N__8824),
            .lcout(un1_D_UU_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_13_19_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_13_19_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_13_19_2  (
            .in0(N__10405),
            .in1(N__8774),
            .in2(_gnd_net_),
            .in3(N__8760),
            .lcout(un1_D_UU_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_13_19_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_13_19_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_13_19_5  (
            .in0(N__8686),
            .in1(N__8645),
            .in2(_gnd_net_),
            .in3(N__10404),
            .lcout(un1_D_UM_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_13_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_13_20_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_13_20_1  (
            .in0(N__11167),
            .in1(N__8618),
            .in2(_gnd_net_),
            .in3(N__8596),
            .lcout(un1_D_UU_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_13_20_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_13_20_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_13_20_2  (
            .in0(N__10407),
            .in1(N__8540),
            .in2(_gnd_net_),
            .in3(N__8517),
            .lcout(un1_D_UM_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_13_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_13_20_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_13_20_3  (
            .in0(N__8448),
            .in1(N__8408),
            .in2(_gnd_net_),
            .in3(N__10408),
            .lcout(un1_D_UU_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_13_20_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_13_20_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_13_20_4  (
            .in0(N__10409),
            .in1(N__8381),
            .in2(_gnd_net_),
            .in3(N__8371),
            .lcout(un1_D_UU_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_040_iobuf_RNO_3_LC_14_11_2.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_3_LC_14_11_2.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_3_LC_14_11_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_040_iobuf_RNO_3_LC_14_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9038),
            .lcout(N_224_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_14_12_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_14_12_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_14_12_2  (
            .in0(N__10327),
            .in1(N__9164),
            .in2(_gnd_net_),
            .in3(N__9145),
            .lcout(un1_D_UM_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_14_13_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_14_13_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_14_13_0  (
            .in0(N__9101),
            .in1(N__9094),
            .in2(_gnd_net_),
            .in3(N__10379),
            .lcout(un1_D_UM_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep19_i_ess_LC_14_14_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep19_i_ess_LC_14_14_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep19_i_ess_LC_14_14_1 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep19_i_ess_LC_14_14_1  (
            .in0(N__9701),
            .in1(_gnd_net_),
            .in2(N__10011),
            .in3(_gnd_net_),
            .lcout(READ_CYCLE_ACTIVE_rep19_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9399),
            .ce(N__9313),
            .sr(N__9246));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep16_i_ess_LC_14_14_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep16_i_ess_LC_14_14_2 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep16_i_ess_LC_14_14_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep16_i_ess_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(N__9939),
            .in2(_gnd_net_),
            .in3(N__9700),
            .lcout(READ_CYCLE_ACTIVE_rep16_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9399),
            .ce(N__9313),
            .sr(N__9246));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep29_i_ess_LC_14_14_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep29_i_ess_LC_14_14_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep29_i_ess_LC_14_14_5 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep29_i_ess_LC_14_14_5  (
            .in0(N__9702),
            .in1(_gnd_net_),
            .in2(N__10012),
            .in3(_gnd_net_),
            .lcout(READ_CYCLE_ACTIVE_rep29_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9399),
            .ce(N__9313),
            .sr(N__9246));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep31_i_ess_LC_14_14_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep31_i_ess_LC_14_14_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep31_i_ess_LC_14_14_7 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep31_i_ess_LC_14_14_7  (
            .in0(N__9703),
            .in1(_gnd_net_),
            .in2(N__10013),
            .in3(_gnd_net_),
            .lcout(READ_CYCLE_ACTIVE_rep31_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9399),
            .ce(N__9313),
            .sr(N__9246));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_14_15_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_14_15_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_14_15_1  (
            .in0(N__9025),
            .in1(N__8978),
            .in2(_gnd_net_),
            .in3(N__10381),
            .lcout(un1_D_UM_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_040_iobuf_RNO_3_LC_14_16_0.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_3_LC_14_16_0.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_3_LC_14_16_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_040_iobuf_RNO_3_LC_14_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8951),
            .lcout(N_216_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_14_18_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_14_18_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_14_18_4  (
            .in0(N__8920),
            .in1(N__8879),
            .in2(_gnd_net_),
            .in3(N__11168),
            .lcout(un1_D_UU_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_14_19_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_14_19_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_14_19_7  (
            .in0(N__10461),
            .in1(N__10421),
            .in2(_gnd_net_),
            .in3(N__10406),
            .lcout(un1_D_UU_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_040_iobuf_RNO_6_LC_15_12_4.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_6_LC_15_12_4.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_6_LC_15_12_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UM_040_iobuf_RNO_6_LC_15_12_4 (
            .in0(N__10271),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_219_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_040_iobuf_RNO_7_LC_15_18_1.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_7_LC_15_18_1.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_7_LC_15_18_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_040_iobuf_RNO_7_LC_15_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10241),
            .lcout(N_220_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_5_LC_16_7_3.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_5_LC_16_7_3.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_5_LC_16_7_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_040_iobuf_RNO_5_LC_16_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10208),
            .lcout(N_234_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_16_11_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_16_11_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_16_11_7  (
            .in0(N__10174),
            .in1(N__10133),
            .in2(_gnd_net_),
            .in3(N__11129),
            .lcout(un1_D_UM_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep10_i_ess_LC_16_14_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep10_i_ess_LC_16_14_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep10_i_ess_LC_16_14_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep10_i_ess_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(N__9860),
            .in2(_gnd_net_),
            .in3(N__9704),
            .lcout(READ_CYCLE_ACTIVE_rep10_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9407),
            .ce(N__9314),
            .sr(N__9247));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep20_i_ess_LC_16_14_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep20_i_ess_LC_16_14_2 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep20_i_ess_LC_16_14_2 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep20_i_ess_LC_16_14_2  (
            .in0(N__9705),
            .in1(_gnd_net_),
            .in2(N__9938),
            .in3(_gnd_net_),
            .lcout(READ_CYCLE_ACTIVE_rep20_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9407),
            .ce(N__9314),
            .sr(N__9247));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep22_i_ess_LC_16_14_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep22_i_ess_LC_16_14_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep22_i_ess_LC_16_14_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep22_i_ess_LC_16_14_5  (
            .in0(_gnd_net_),
            .in1(N__9864),
            .in2(_gnd_net_),
            .in3(N__9706),
            .lcout(READ_CYCLE_ACTIVE_rep22_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9407),
            .ce(N__9314),
            .sr(N__9247));
    defparam D_LL_040_iobuf_RNO_3_LC_17_1_4.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_3_LC_17_1_4.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_3_LC_17_1_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LL_040_iobuf_RNO_3_LC_17_1_4 (
            .in0(N__10793),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_232_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_040_iobuf_RNO_2_LC_17_6_3.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_2_LC_17_6_3.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_2_LC_17_6_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_040_iobuf_RNO_2_LC_17_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10760),
            .lcout(N_223_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_040_iobuf_RNO_0_LC_17_17_7.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_0_LC_17_17_7.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_0_LC_17_17_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_040_iobuf_RNO_0_LC_17_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10730),
            .lcout(N_205_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_040_iobuf_RNO_7_LC_17_18_5.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_7_LC_17_18_5.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_7_LC_17_18_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_040_iobuf_RNO_7_LC_17_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10694),
            .lcout(N_212_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_18_10_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_18_10_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_18_10_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_18_10_3  (
            .in0(N__10661),
            .in1(N__10639),
            .in2(_gnd_net_),
            .in3(N__11151),
            .lcout(un1_D_UM_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_7_LC_18_14_1.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_7_LC_18_14_1.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_7_LC_18_14_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LL_040_iobuf_RNO_7_LC_18_14_1 (
            .in0(N__10589),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_236_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_040_iobuf_RNO_6_LC_18_14_4.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_6_LC_18_14_4.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_6_LC_18_14_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LM_040_iobuf_RNO_6_LC_18_14_4 (
            .in0(N__10565),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_227_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_040_iobuf_RNO_5_LC_18_17_1.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_5_LC_18_17_1.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_5_LC_18_17_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_040_iobuf_RNO_5_LC_18_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10538),
            .lcout(N_218_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_040_iobuf_RNO_4_LC_18_17_2.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_4_LC_18_17_2.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_4_LC_18_17_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_040_iobuf_RNO_4_LC_18_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10505),
            .lcout(N_209_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_18_19_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_18_19_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_18_19_1  (
            .in0(N__11504),
            .in1(N__11482),
            .in2(_gnd_net_),
            .in3(N__11169),
            .lcout(un1_D_UM_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_4_LC_19_6_0.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_4_LC_19_6_0.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_4_LC_19_6_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LL_040_iobuf_RNO_4_LC_19_6_0 (
            .in0(N__11411),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_233_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_6_LC_19_6_2.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_6_LC_19_6_2.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_6_LC_19_6_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LL_040_iobuf_RNO_6_LC_19_6_2 (
            .in0(N__11384),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_235_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_040_iobuf_RNO_1_LC_19_6_6.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_1_LC_19_6_6.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_1_LC_19_6_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LM_040_iobuf_RNO_1_LC_19_6_6 (
            .in0(N__11351),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_222_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_19_19_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_19_19_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_19_19_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_19_19_5  (
            .in0(N__11321),
            .in1(N__11302),
            .in2(_gnd_net_),
            .in3(N__11170),
            .lcout(un1_D_UM_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_19_20_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_19_20_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_19_20_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_19_20_2  (
            .in0(N__11224),
            .in1(N__11189),
            .in2(_gnd_net_),
            .in3(N__11171),
            .lcout(un1_D_UM_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_1_LC_20_9_2.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_1_LC_20_9_2.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_1_LC_20_9_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LL_040_iobuf_RNO_1_LC_20_9_2 (
            .in0(N__10850),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_230_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_040_iobuf_RNO_2_LC_20_10_6.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_2_LC_20_10_6.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_2_LC_20_10_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_040_iobuf_RNO_2_LC_20_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10814),
            .lcout(N_215_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_040_iobuf_RNO_5_LC_20_11_2.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_5_LC_20_11_2.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_5_LC_20_11_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LM_040_iobuf_RNO_5_LC_20_11_2 (
            .in0(N__11750),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_226_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_0_LC_20_11_5.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_0_LC_20_11_5.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_0_LC_20_11_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_040_iobuf_RNO_0_LC_20_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11726),
            .lcout(N_229_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_040_iobuf_RNO_1_LC_20_15_6.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_1_LC_20_15_6.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_1_LC_20_15_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UM_040_iobuf_RNO_1_LC_20_15_6 (
            .in0(N__11690),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_214_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_040_iobuf_RNO_4_LC_20_18_2.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_4_LC_20_18_2.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_4_LC_20_18_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_040_iobuf_RNO_4_LC_20_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11657),
            .lcout(N_217_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_040_iobuf_RNO_0_LC_22_12_3.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_0_LC_22_12_3.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_0_LC_22_12_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_040_iobuf_RNO_0_LC_22_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11621),
            .lcout(N_213_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_040_iobuf_RNO_7_LC_22_15_6.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_7_LC_22_15_6.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_7_LC_22_15_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_040_iobuf_RNO_7_LC_22_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11591),
            .lcout(N_228_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_040_iobuf_RNO_4_LC_23_14_2.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_4_LC_23_14_2.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_4_LC_23_14_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_040_iobuf_RNO_4_LC_23_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11561),
            .lcout(N_225_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_040_iobuf_RNO_3_LC_23_19_4.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_3_LC_23_19_4.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_3_LC_23_19_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_040_iobuf_RNO_3_LC_23_19_4 (
            .in0(N__11531),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_208_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_040_iobuf_RNO_0_LC_24_7_2.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_0_LC_24_7_2.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_0_LC_24_7_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_040_iobuf_RNO_0_LC_24_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11783),
            .lcout(N_221_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U111_TOP

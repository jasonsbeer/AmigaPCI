// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Sep 11 2025 19:59:55

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U111_TOP" view "INTERFACE"

module U111_TOP (
    D_LM_AMIGA,
    D_UM_AMIGA,
    D_LL_AMIGA,
    D_UU_AMIGA,
    D_LL_040,
    D_UU_040,
    D_LM_040,
    D_UM_040,
    A_AMIGA,
    A_040,
    SIZ,
    TBIn,
    TEAn,
    TSn,
    RESETn,
    CLKRAMA,
    PORTSIZE,
    DMAAn,
    TEA_CPUn,
    LBENn,
    CLK40B,
    TBI_CPUn,
    TAn,
    CPUBGn,
    BUFENn,
    RnW,
    CLK80_CPU,
    BUFDIR,
    TCI_CPUn,
    TS_CPUn,
    CLKRAMB,
    CLK40A,
    TCIn,
    CLK40C,
    CLK40_IN,
    BBn,
    TACKn,
    BGn);

    inout [7:0] D_LM_AMIGA;
    inout [7:0] D_UM_AMIGA;
    inout [7:0] D_LL_AMIGA;
    inout [7:0] D_UU_AMIGA;
    inout [7:0] D_LL_040;
    inout [7:0] D_UU_040;
    inout [7:0] D_LM_040;
    inout [7:0] D_UM_040;
    output [1:0] A_AMIGA;
    input [1:0] A_040;
    input [1:0] SIZ;
    input TBIn;
    input TEAn;
    output TSn;
    input RESETn;
    output CLKRAMA;
    input PORTSIZE;
    output DMAAn;
    output TEA_CPUn;
    input LBENn;
    output CLK40B;
    output TBI_CPUn;
    inout TAn;
    output CPUBGn;
    output BUFENn;
    input RnW;
    output CLK80_CPU;
    output BUFDIR;
    output TCI_CPUn;
    inout TS_CPUn;
    output CLKRAMB;
    output CLK40A;
    input TCIn;
    output CLK40C;
    input CLK40_IN;
    input BBn;
    inout TACKn;
    input BGn;

    wire N__9524;
    wire N__9508;
    wire N__9507;
    wire N__9506;
    wire N__9499;
    wire N__9498;
    wire N__9497;
    wire N__9490;
    wire N__9489;
    wire N__9488;
    wire N__9481;
    wire N__9480;
    wire N__9479;
    wire N__9472;
    wire N__9471;
    wire N__9470;
    wire N__9463;
    wire N__9462;
    wire N__9461;
    wire N__9454;
    wire N__9453;
    wire N__9452;
    wire N__9445;
    wire N__9444;
    wire N__9443;
    wire N__9436;
    wire N__9435;
    wire N__9434;
    wire N__9427;
    wire N__9426;
    wire N__9425;
    wire N__9418;
    wire N__9417;
    wire N__9416;
    wire N__9409;
    wire N__9408;
    wire N__9407;
    wire N__9400;
    wire N__9399;
    wire N__9398;
    wire N__9391;
    wire N__9390;
    wire N__9389;
    wire N__9382;
    wire N__9381;
    wire N__9380;
    wire N__9373;
    wire N__9372;
    wire N__9371;
    wire N__9364;
    wire N__9363;
    wire N__9362;
    wire N__9355;
    wire N__9354;
    wire N__9353;
    wire N__9346;
    wire N__9345;
    wire N__9344;
    wire N__9337;
    wire N__9336;
    wire N__9335;
    wire N__9328;
    wire N__9327;
    wire N__9326;
    wire N__9319;
    wire N__9318;
    wire N__9317;
    wire N__9310;
    wire N__9309;
    wire N__9308;
    wire N__9301;
    wire N__9300;
    wire N__9299;
    wire N__9292;
    wire N__9291;
    wire N__9290;
    wire N__9283;
    wire N__9282;
    wire N__9281;
    wire N__9274;
    wire N__9273;
    wire N__9272;
    wire N__9265;
    wire N__9264;
    wire N__9263;
    wire N__9256;
    wire N__9255;
    wire N__9254;
    wire N__9247;
    wire N__9246;
    wire N__9245;
    wire N__9238;
    wire N__9237;
    wire N__9236;
    wire N__9229;
    wire N__9228;
    wire N__9227;
    wire N__9220;
    wire N__9219;
    wire N__9218;
    wire N__9211;
    wire N__9210;
    wire N__9209;
    wire N__9202;
    wire N__9201;
    wire N__9200;
    wire N__9193;
    wire N__9192;
    wire N__9191;
    wire N__9184;
    wire N__9183;
    wire N__9182;
    wire N__9175;
    wire N__9174;
    wire N__9173;
    wire N__9166;
    wire N__9165;
    wire N__9164;
    wire N__9157;
    wire N__9156;
    wire N__9155;
    wire N__9148;
    wire N__9147;
    wire N__9146;
    wire N__9139;
    wire N__9138;
    wire N__9137;
    wire N__9130;
    wire N__9129;
    wire N__9128;
    wire N__9121;
    wire N__9120;
    wire N__9119;
    wire N__9112;
    wire N__9111;
    wire N__9110;
    wire N__9103;
    wire N__9102;
    wire N__9101;
    wire N__9094;
    wire N__9093;
    wire N__9092;
    wire N__9085;
    wire N__9084;
    wire N__9083;
    wire N__9076;
    wire N__9075;
    wire N__9074;
    wire N__9067;
    wire N__9066;
    wire N__9065;
    wire N__9058;
    wire N__9057;
    wire N__9056;
    wire N__9049;
    wire N__9048;
    wire N__9047;
    wire N__9040;
    wire N__9039;
    wire N__9038;
    wire N__9031;
    wire N__9030;
    wire N__9029;
    wire N__9022;
    wire N__9021;
    wire N__9020;
    wire N__9013;
    wire N__9012;
    wire N__9011;
    wire N__9004;
    wire N__9003;
    wire N__9002;
    wire N__8995;
    wire N__8994;
    wire N__8993;
    wire N__8986;
    wire N__8985;
    wire N__8984;
    wire N__8977;
    wire N__8976;
    wire N__8975;
    wire N__8968;
    wire N__8967;
    wire N__8966;
    wire N__8959;
    wire N__8958;
    wire N__8957;
    wire N__8950;
    wire N__8949;
    wire N__8948;
    wire N__8941;
    wire N__8940;
    wire N__8939;
    wire N__8932;
    wire N__8931;
    wire N__8930;
    wire N__8923;
    wire N__8922;
    wire N__8921;
    wire N__8914;
    wire N__8913;
    wire N__8912;
    wire N__8905;
    wire N__8904;
    wire N__8903;
    wire N__8896;
    wire N__8895;
    wire N__8894;
    wire N__8887;
    wire N__8886;
    wire N__8885;
    wire N__8878;
    wire N__8877;
    wire N__8876;
    wire N__8869;
    wire N__8868;
    wire N__8867;
    wire N__8860;
    wire N__8859;
    wire N__8858;
    wire N__8851;
    wire N__8850;
    wire N__8849;
    wire N__8842;
    wire N__8841;
    wire N__8840;
    wire N__8833;
    wire N__8832;
    wire N__8831;
    wire N__8824;
    wire N__8823;
    wire N__8822;
    wire N__8815;
    wire N__8814;
    wire N__8813;
    wire N__8806;
    wire N__8805;
    wire N__8804;
    wire N__8797;
    wire N__8796;
    wire N__8795;
    wire N__8788;
    wire N__8787;
    wire N__8786;
    wire N__8779;
    wire N__8778;
    wire N__8777;
    wire N__8770;
    wire N__8769;
    wire N__8768;
    wire N__8761;
    wire N__8760;
    wire N__8759;
    wire N__8752;
    wire N__8751;
    wire N__8750;
    wire N__8743;
    wire N__8742;
    wire N__8741;
    wire N__8734;
    wire N__8733;
    wire N__8732;
    wire N__8725;
    wire N__8724;
    wire N__8723;
    wire N__8716;
    wire N__8715;
    wire N__8714;
    wire N__8707;
    wire N__8706;
    wire N__8705;
    wire N__8698;
    wire N__8697;
    wire N__8696;
    wire N__8689;
    wire N__8688;
    wire N__8687;
    wire N__8680;
    wire N__8679;
    wire N__8678;
    wire N__8671;
    wire N__8670;
    wire N__8669;
    wire N__8662;
    wire N__8661;
    wire N__8660;
    wire N__8653;
    wire N__8652;
    wire N__8651;
    wire N__8634;
    wire N__8631;
    wire N__8628;
    wire N__8625;
    wire N__8622;
    wire N__8619;
    wire N__8616;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8608;
    wire N__8605;
    wire N__8602;
    wire N__8599;
    wire N__8596;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8559;
    wire N__8556;
    wire N__8553;
    wire N__8550;
    wire N__8547;
    wire N__8544;
    wire N__8541;
    wire N__8538;
    wire N__8535;
    wire N__8532;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8519;
    wire N__8516;
    wire N__8513;
    wire N__8510;
    wire N__8507;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8484;
    wire N__8481;
    wire N__8478;
    wire N__8475;
    wire N__8472;
    wire N__8469;
    wire N__8466;
    wire N__8463;
    wire N__8460;
    wire N__8457;
    wire N__8454;
    wire N__8451;
    wire N__8448;
    wire N__8445;
    wire N__8442;
    wire N__8439;
    wire N__8436;
    wire N__8433;
    wire N__8430;
    wire N__8427;
    wire N__8426;
    wire N__8423;
    wire N__8422;
    wire N__8419;
    wire N__8416;
    wire N__8413;
    wire N__8410;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8382;
    wire N__8379;
    wire N__8376;
    wire N__8373;
    wire N__8370;
    wire N__8367;
    wire N__8364;
    wire N__8361;
    wire N__8358;
    wire N__8355;
    wire N__8352;
    wire N__8349;
    wire N__8348;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8330;
    wire N__8327;
    wire N__8324;
    wire N__8319;
    wire N__8316;
    wire N__8313;
    wire N__8310;
    wire N__8307;
    wire N__8304;
    wire N__8301;
    wire N__8298;
    wire N__8295;
    wire N__8292;
    wire N__8289;
    wire N__8286;
    wire N__8283;
    wire N__8280;
    wire N__8277;
    wire N__8274;
    wire N__8271;
    wire N__8268;
    wire N__8265;
    wire N__8264;
    wire N__8261;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8249;
    wire N__8246;
    wire N__8243;
    wire N__8240;
    wire N__8237;
    wire N__8234;
    wire N__8231;
    wire N__8228;
    wire N__8225;
    wire N__8222;
    wire N__8217;
    wire N__8216;
    wire N__8215;
    wire N__8214;
    wire N__8213;
    wire N__8212;
    wire N__8211;
    wire N__8210;
    wire N__8209;
    wire N__8208;
    wire N__8207;
    wire N__8206;
    wire N__8201;
    wire N__8198;
    wire N__8197;
    wire N__8192;
    wire N__8187;
    wire N__8186;
    wire N__8183;
    wire N__8178;
    wire N__8175;
    wire N__8174;
    wire N__8173;
    wire N__8172;
    wire N__8169;
    wire N__8168;
    wire N__8167;
    wire N__8162;
    wire N__8159;
    wire N__8156;
    wire N__8153;
    wire N__8150;
    wire N__8149;
    wire N__8148;
    wire N__8143;
    wire N__8140;
    wire N__8139;
    wire N__8138;
    wire N__8137;
    wire N__8136;
    wire N__8135;
    wire N__8134;
    wire N__8131;
    wire N__8130;
    wire N__8129;
    wire N__8126;
    wire N__8123;
    wire N__8120;
    wire N__8115;
    wire N__8110;
    wire N__8103;
    wire N__8098;
    wire N__8093;
    wire N__8090;
    wire N__8085;
    wire N__8080;
    wire N__8077;
    wire N__8074;
    wire N__8071;
    wire N__8068;
    wire N__8067;
    wire N__8062;
    wire N__8057;
    wire N__8054;
    wire N__8049;
    wire N__8044;
    wire N__8037;
    wire N__8030;
    wire N__8027;
    wire N__8026;
    wire N__8025;
    wire N__8024;
    wire N__8021;
    wire N__8018;
    wire N__8013;
    wire N__8006;
    wire N__8003;
    wire N__7998;
    wire N__7995;
    wire N__7980;
    wire N__7977;
    wire N__7974;
    wire N__7971;
    wire N__7968;
    wire N__7965;
    wire N__7962;
    wire N__7959;
    wire N__7956;
    wire N__7953;
    wire N__7952;
    wire N__7949;
    wire N__7946;
    wire N__7943;
    wire N__7942;
    wire N__7939;
    wire N__7936;
    wire N__7933;
    wire N__7930;
    wire N__7925;
    wire N__7922;
    wire N__7919;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7902;
    wire N__7899;
    wire N__7896;
    wire N__7893;
    wire N__7890;
    wire N__7887;
    wire N__7884;
    wire N__7883;
    wire N__7882;
    wire N__7881;
    wire N__7880;
    wire N__7877;
    wire N__7876;
    wire N__7867;
    wire N__7866;
    wire N__7865;
    wire N__7864;
    wire N__7863;
    wire N__7862;
    wire N__7861;
    wire N__7858;
    wire N__7855;
    wire N__7852;
    wire N__7845;
    wire N__7842;
    wire N__7837;
    wire N__7824;
    wire N__7821;
    wire N__7820;
    wire N__7817;
    wire N__7814;
    wire N__7811;
    wire N__7808;
    wire N__7807;
    wire N__7806;
    wire N__7805;
    wire N__7802;
    wire N__7799;
    wire N__7792;
    wire N__7791;
    wire N__7788;
    wire N__7785;
    wire N__7782;
    wire N__7779;
    wire N__7776;
    wire N__7775;
    wire N__7770;
    wire N__7769;
    wire N__7766;
    wire N__7763;
    wire N__7760;
    wire N__7757;
    wire N__7754;
    wire N__7751;
    wire N__7746;
    wire N__7741;
    wire N__7738;
    wire N__7735;
    wire N__7732;
    wire N__7725;
    wire N__7724;
    wire N__7721;
    wire N__7720;
    wire N__7719;
    wire N__7716;
    wire N__7713;
    wire N__7710;
    wire N__7705;
    wire N__7704;
    wire N__7701;
    wire N__7698;
    wire N__7695;
    wire N__7692;
    wire N__7689;
    wire N__7686;
    wire N__7681;
    wire N__7676;
    wire N__7673;
    wire N__7670;
    wire N__7667;
    wire N__7664;
    wire N__7661;
    wire N__7656;
    wire N__7655;
    wire N__7654;
    wire N__7653;
    wire N__7650;
    wire N__7647;
    wire N__7646;
    wire N__7645;
    wire N__7644;
    wire N__7641;
    wire N__7638;
    wire N__7637;
    wire N__7636;
    wire N__7635;
    wire N__7634;
    wire N__7633;
    wire N__7632;
    wire N__7631;
    wire N__7630;
    wire N__7629;
    wire N__7624;
    wire N__7621;
    wire N__7618;
    wire N__7615;
    wire N__7614;
    wire N__7611;
    wire N__7610;
    wire N__7607;
    wire N__7604;
    wire N__7601;
    wire N__7600;
    wire N__7597;
    wire N__7594;
    wire N__7591;
    wire N__7588;
    wire N__7585;
    wire N__7582;
    wire N__7579;
    wire N__7570;
    wire N__7567;
    wire N__7564;
    wire N__7561;
    wire N__7560;
    wire N__7559;
    wire N__7558;
    wire N__7551;
    wire N__7548;
    wire N__7547;
    wire N__7546;
    wire N__7541;
    wire N__7530;
    wire N__7529;
    wire N__7528;
    wire N__7527;
    wire N__7524;
    wire N__7521;
    wire N__7516;
    wire N__7513;
    wire N__7510;
    wire N__7507;
    wire N__7502;
    wire N__7499;
    wire N__7496;
    wire N__7495;
    wire N__7494;
    wire N__7491;
    wire N__7488;
    wire N__7485;
    wire N__7482;
    wire N__7481;
    wire N__7480;
    wire N__7479;
    wire N__7476;
    wire N__7473;
    wire N__7470;
    wire N__7461;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7443;
    wire N__7440;
    wire N__7437;
    wire N__7434;
    wire N__7431;
    wire N__7428;
    wire N__7425;
    wire N__7420;
    wire N__7415;
    wire N__7410;
    wire N__7403;
    wire N__7398;
    wire N__7395;
    wire N__7392;
    wire N__7389;
    wire N__7386;
    wire N__7383;
    wire N__7380;
    wire N__7373;
    wire N__7368;
    wire N__7365;
    wire N__7360;
    wire N__7357;
    wire N__7350;
    wire N__7349;
    wire N__7348;
    wire N__7345;
    wire N__7344;
    wire N__7343;
    wire N__7342;
    wire N__7341;
    wire N__7340;
    wire N__7339;
    wire N__7334;
    wire N__7333;
    wire N__7330;
    wire N__7327;
    wire N__7324;
    wire N__7323;
    wire N__7322;
    wire N__7321;
    wire N__7320;
    wire N__7319;
    wire N__7310;
    wire N__7309;
    wire N__7306;
    wire N__7303;
    wire N__7298;
    wire N__7295;
    wire N__7292;
    wire N__7289;
    wire N__7286;
    wire N__7281;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7269;
    wire N__7258;
    wire N__7255;
    wire N__7252;
    wire N__7247;
    wire N__7244;
    wire N__7239;
    wire N__7236;
    wire N__7227;
    wire N__7224;
    wire N__7221;
    wire N__7218;
    wire N__7215;
    wire N__7212;
    wire N__7211;
    wire N__7210;
    wire N__7207;
    wire N__7204;
    wire N__7201;
    wire N__7194;
    wire N__7191;
    wire N__7188;
    wire N__7185;
    wire N__7182;
    wire N__7179;
    wire N__7178;
    wire N__7177;
    wire N__7174;
    wire N__7171;
    wire N__7168;
    wire N__7161;
    wire N__7158;
    wire N__7155;
    wire N__7152;
    wire N__7149;
    wire N__7146;
    wire N__7143;
    wire N__7140;
    wire N__7137;
    wire N__7136;
    wire N__7135;
    wire N__7134;
    wire N__7133;
    wire N__7132;
    wire N__7131;
    wire N__7130;
    wire N__7129;
    wire N__7128;
    wire N__7127;
    wire N__7126;
    wire N__7125;
    wire N__7124;
    wire N__7123;
    wire N__7122;
    wire N__7089;
    wire N__7086;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7076;
    wire N__7075;
    wire N__7072;
    wire N__7069;
    wire N__7066;
    wire N__7063;
    wire N__7060;
    wire N__7057;
    wire N__7054;
    wire N__7047;
    wire N__7046;
    wire N__7043;
    wire N__7040;
    wire N__7039;
    wire N__7036;
    wire N__7033;
    wire N__7030;
    wire N__7027;
    wire N__7024;
    wire N__7021;
    wire N__7014;
    wire N__7011;
    wire N__7008;
    wire N__7007;
    wire N__7006;
    wire N__7003;
    wire N__7000;
    wire N__6997;
    wire N__6994;
    wire N__6989;
    wire N__6986;
    wire N__6983;
    wire N__6980;
    wire N__6977;
    wire N__6972;
    wire N__6969;
    wire N__6966;
    wire N__6963;
    wire N__6960;
    wire N__6957;
    wire N__6954;
    wire N__6951;
    wire N__6948;
    wire N__6945;
    wire N__6942;
    wire N__6941;
    wire N__6940;
    wire N__6937;
    wire N__6934;
    wire N__6931;
    wire N__6926;
    wire N__6923;
    wire N__6918;
    wire N__6915;
    wire N__6912;
    wire N__6909;
    wire N__6906;
    wire N__6903;
    wire N__6900;
    wire N__6897;
    wire N__6894;
    wire N__6891;
    wire N__6888;
    wire N__6885;
    wire N__6882;
    wire N__6879;
    wire N__6876;
    wire N__6875;
    wire N__6872;
    wire N__6869;
    wire N__6866;
    wire N__6863;
    wire N__6862;
    wire N__6861;
    wire N__6858;
    wire N__6855;
    wire N__6850;
    wire N__6849;
    wire N__6846;
    wire N__6843;
    wire N__6840;
    wire N__6839;
    wire N__6836;
    wire N__6835;
    wire N__6832;
    wire N__6829;
    wire N__6826;
    wire N__6823;
    wire N__6820;
    wire N__6817;
    wire N__6814;
    wire N__6807;
    wire N__6802;
    wire N__6797;
    wire N__6794;
    wire N__6789;
    wire N__6786;
    wire N__6783;
    wire N__6780;
    wire N__6777;
    wire N__6774;
    wire N__6771;
    wire N__6768;
    wire N__6765;
    wire N__6762;
    wire N__6759;
    wire N__6756;
    wire N__6753;
    wire N__6750;
    wire N__6747;
    wire N__6744;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6732;
    wire N__6729;
    wire N__6728;
    wire N__6725;
    wire N__6722;
    wire N__6719;
    wire N__6718;
    wire N__6715;
    wire N__6712;
    wire N__6709;
    wire N__6706;
    wire N__6701;
    wire N__6698;
    wire N__6695;
    wire N__6692;
    wire N__6689;
    wire N__6684;
    wire N__6681;
    wire N__6678;
    wire N__6675;
    wire N__6672;
    wire N__6669;
    wire N__6666;
    wire N__6663;
    wire N__6660;
    wire N__6657;
    wire N__6654;
    wire N__6651;
    wire N__6648;
    wire N__6645;
    wire N__6642;
    wire N__6639;
    wire N__6636;
    wire N__6633;
    wire N__6630;
    wire N__6627;
    wire N__6624;
    wire N__6621;
    wire N__6618;
    wire N__6615;
    wire N__6612;
    wire N__6609;
    wire N__6608;
    wire N__6605;
    wire N__6602;
    wire N__6599;
    wire N__6596;
    wire N__6591;
    wire N__6588;
    wire N__6585;
    wire N__6582;
    wire N__6579;
    wire N__6576;
    wire N__6573;
    wire N__6570;
    wire N__6567;
    wire N__6564;
    wire N__6561;
    wire N__6558;
    wire N__6555;
    wire N__6552;
    wire N__6549;
    wire N__6546;
    wire N__6543;
    wire N__6540;
    wire N__6537;
    wire N__6534;
    wire N__6531;
    wire N__6528;
    wire N__6525;
    wire N__6522;
    wire N__6519;
    wire N__6516;
    wire N__6513;
    wire N__6510;
    wire N__6507;
    wire N__6504;
    wire N__6503;
    wire N__6502;
    wire N__6499;
    wire N__6498;
    wire N__6495;
    wire N__6492;
    wire N__6491;
    wire N__6488;
    wire N__6485;
    wire N__6484;
    wire N__6481;
    wire N__6478;
    wire N__6475;
    wire N__6472;
    wire N__6469;
    wire N__6466;
    wire N__6459;
    wire N__6452;
    wire N__6449;
    wire N__6446;
    wire N__6443;
    wire N__6440;
    wire N__6435;
    wire N__6432;
    wire N__6429;
    wire N__6426;
    wire N__6423;
    wire N__6420;
    wire N__6417;
    wire N__6414;
    wire N__6411;
    wire N__6408;
    wire N__6405;
    wire N__6402;
    wire N__6401;
    wire N__6400;
    wire N__6397;
    wire N__6394;
    wire N__6391;
    wire N__6388;
    wire N__6383;
    wire N__6378;
    wire N__6375;
    wire N__6372;
    wire N__6369;
    wire N__6366;
    wire N__6365;
    wire N__6362;
    wire N__6361;
    wire N__6358;
    wire N__6355;
    wire N__6352;
    wire N__6345;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6337;
    wire N__6336;
    wire N__6335;
    wire N__6334;
    wire N__6333;
    wire N__6330;
    wire N__6327;
    wire N__6324;
    wire N__6321;
    wire N__6318;
    wire N__6313;
    wire N__6300;
    wire N__6299;
    wire N__6298;
    wire N__6297;
    wire N__6296;
    wire N__6295;
    wire N__6294;
    wire N__6293;
    wire N__6276;
    wire N__6273;
    wire N__6270;
    wire N__6269;
    wire N__6264;
    wire N__6263;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6255;
    wire N__6254;
    wire N__6253;
    wire N__6252;
    wire N__6249;
    wire N__6244;
    wire N__6239;
    wire N__6234;
    wire N__6231;
    wire N__6224;
    wire N__6221;
    wire N__6218;
    wire N__6215;
    wire N__6214;
    wire N__6211;
    wire N__6208;
    wire N__6205;
    wire N__6202;
    wire N__6197;
    wire N__6192;
    wire N__6189;
    wire N__6186;
    wire N__6185;
    wire N__6184;
    wire N__6183;
    wire N__6180;
    wire N__6177;
    wire N__6174;
    wire N__6171;
    wire N__6162;
    wire N__6159;
    wire N__6158;
    wire N__6157;
    wire N__6156;
    wire N__6155;
    wire N__6152;
    wire N__6151;
    wire N__6150;
    wire N__6149;
    wire N__6148;
    wire N__6139;
    wire N__6136;
    wire N__6129;
    wire N__6126;
    wire N__6117;
    wire N__6114;
    wire N__6111;
    wire N__6108;
    wire N__6105;
    wire N__6102;
    wire N__6099;
    wire N__6098;
    wire N__6095;
    wire N__6092;
    wire N__6089;
    wire N__6086;
    wire N__6083;
    wire N__6080;
    wire N__6077;
    wire N__6074;
    wire N__6071;
    wire N__6068;
    wire N__6065;
    wire N__6062;
    wire N__6057;
    wire N__6054;
    wire N__6051;
    wire N__6048;
    wire N__6045;
    wire N__6042;
    wire N__6039;
    wire N__6038;
    wire N__6035;
    wire N__6032;
    wire N__6029;
    wire N__6028;
    wire N__6025;
    wire N__6022;
    wire N__6019;
    wire N__6016;
    wire N__6011;
    wire N__6008;
    wire N__6005;
    wire N__6000;
    wire N__5997;
    wire N__5994;
    wire N__5991;
    wire N__5988;
    wire N__5987;
    wire N__5984;
    wire N__5981;
    wire N__5976;
    wire N__5973;
    wire N__5970;
    wire N__5967;
    wire N__5964;
    wire N__5961;
    wire N__5958;
    wire N__5955;
    wire N__5952;
    wire N__5949;
    wire N__5946;
    wire N__5943;
    wire N__5942;
    wire N__5939;
    wire N__5936;
    wire N__5933;
    wire N__5932;
    wire N__5929;
    wire N__5926;
    wire N__5923;
    wire N__5920;
    wire N__5915;
    wire N__5912;
    wire N__5909;
    wire N__5906;
    wire N__5903;
    wire N__5900;
    wire N__5897;
    wire N__5892;
    wire N__5889;
    wire N__5886;
    wire N__5883;
    wire N__5880;
    wire N__5877;
    wire N__5874;
    wire N__5871;
    wire N__5868;
    wire N__5865;
    wire N__5862;
    wire N__5859;
    wire N__5856;
    wire N__5855;
    wire N__5852;
    wire N__5849;
    wire N__5846;
    wire N__5843;
    wire N__5840;
    wire N__5837;
    wire N__5832;
    wire N__5829;
    wire N__5826;
    wire N__5823;
    wire N__5822;
    wire N__5819;
    wire N__5816;
    wire N__5811;
    wire N__5810;
    wire N__5807;
    wire N__5804;
    wire N__5801;
    wire N__5798;
    wire N__5797;
    wire N__5794;
    wire N__5791;
    wire N__5788;
    wire N__5785;
    wire N__5782;
    wire N__5779;
    wire N__5776;
    wire N__5771;
    wire N__5766;
    wire N__5763;
    wire N__5760;
    wire N__5757;
    wire N__5754;
    wire N__5753;
    wire N__5750;
    wire N__5747;
    wire N__5744;
    wire N__5741;
    wire N__5738;
    wire N__5735;
    wire N__5732;
    wire N__5729;
    wire N__5724;
    wire N__5721;
    wire N__5718;
    wire N__5715;
    wire N__5712;
    wire N__5709;
    wire N__5706;
    wire N__5703;
    wire N__5700;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5681;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5669;
    wire N__5664;
    wire N__5661;
    wire N__5658;
    wire N__5655;
    wire N__5652;
    wire N__5649;
    wire N__5646;
    wire N__5643;
    wire N__5640;
    wire N__5637;
    wire N__5634;
    wire N__5631;
    wire N__5628;
    wire N__5625;
    wire N__5624;
    wire N__5621;
    wire N__5618;
    wire N__5613;
    wire N__5610;
    wire N__5609;
    wire N__5606;
    wire N__5603;
    wire N__5602;
    wire N__5599;
    wire N__5596;
    wire N__5593;
    wire N__5590;
    wire N__5585;
    wire N__5580;
    wire N__5577;
    wire N__5574;
    wire N__5571;
    wire N__5568;
    wire N__5565;
    wire N__5562;
    wire N__5559;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5547;
    wire N__5544;
    wire N__5541;
    wire N__5538;
    wire N__5537;
    wire N__5534;
    wire N__5531;
    wire N__5526;
    wire N__5523;
    wire N__5520;
    wire N__5517;
    wire N__5514;
    wire N__5511;
    wire N__5508;
    wire N__5505;
    wire N__5504;
    wire N__5503;
    wire N__5500;
    wire N__5497;
    wire N__5494;
    wire N__5487;
    wire N__5486;
    wire N__5483;
    wire N__5480;
    wire N__5475;
    wire N__5472;
    wire N__5469;
    wire N__5468;
    wire N__5467;
    wire N__5466;
    wire N__5465;
    wire N__5464;
    wire N__5463;
    wire N__5462;
    wire N__5461;
    wire N__5458;
    wire N__5457;
    wire N__5454;
    wire N__5451;
    wire N__5448;
    wire N__5445;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5435;
    wire N__5434;
    wire N__5433;
    wire N__5432;
    wire N__5431;
    wire N__5430;
    wire N__5427;
    wire N__5424;
    wire N__5421;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5398;
    wire N__5397;
    wire N__5396;
    wire N__5395;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5374;
    wire N__5373;
    wire N__5372;
    wire N__5371;
    wire N__5370;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5351;
    wire N__5340;
    wire N__5337;
    wire N__5334;
    wire N__5331;
    wire N__5328;
    wire N__5327;
    wire N__5326;
    wire N__5325;
    wire N__5324;
    wire N__5323;
    wire N__5312;
    wire N__5301;
    wire N__5298;
    wire N__5295;
    wire N__5292;
    wire N__5289;
    wire N__5286;
    wire N__5285;
    wire N__5284;
    wire N__5281;
    wire N__5270;
    wire N__5267;
    wire N__5266;
    wire N__5263;
    wire N__5260;
    wire N__5257;
    wire N__5252;
    wire N__5249;
    wire N__5244;
    wire N__5239;
    wire N__5236;
    wire N__5233;
    wire N__5228;
    wire N__5223;
    wire N__5220;
    wire N__5219;
    wire N__5216;
    wire N__5213;
    wire N__5208;
    wire N__5205;
    wire N__5202;
    wire N__5199;
    wire N__5196;
    wire N__5193;
    wire N__5190;
    wire N__5189;
    wire N__5186;
    wire N__5183;
    wire N__5182;
    wire N__5181;
    wire N__5176;
    wire N__5173;
    wire N__5170;
    wire N__5163;
    wire N__5162;
    wire N__5159;
    wire N__5158;
    wire N__5155;
    wire N__5154;
    wire N__5151;
    wire N__5146;
    wire N__5143;
    wire N__5136;
    wire N__5133;
    wire N__5130;
    wire N__5129;
    wire N__5128;
    wire N__5127;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5115;
    wire N__5112;
    wire N__5103;
    wire N__5100;
    wire N__5097;
    wire N__5096;
    wire N__5095;
    wire N__5094;
    wire N__5093;
    wire N__5088;
    wire N__5085;
    wire N__5084;
    wire N__5081;
    wire N__5078;
    wire N__5075;
    wire N__5072;
    wire N__5069;
    wire N__5058;
    wire N__5055;
    wire N__5052;
    wire N__5051;
    wire N__5050;
    wire N__5049;
    wire N__5048;
    wire N__5045;
    wire N__5044;
    wire N__5043;
    wire N__5040;
    wire N__5037;
    wire N__5026;
    wire N__5019;
    wire N__5016;
    wire N__5013;
    wire N__5012;
    wire N__5009;
    wire N__5006;
    wire N__5003;
    wire N__5000;
    wire N__4997;
    wire N__4994;
    wire N__4989;
    wire N__4986;
    wire N__4983;
    wire N__4980;
    wire N__4977;
    wire N__4974;
    wire N__4971;
    wire N__4968;
    wire N__4965;
    wire N__4962;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4950;
    wire N__4947;
    wire N__4944;
    wire N__4941;
    wire N__4938;
    wire N__4937;
    wire N__4934;
    wire N__4931;
    wire N__4926;
    wire N__4923;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4905;
    wire N__4902;
    wire N__4899;
    wire N__4896;
    wire N__4893;
    wire N__4892;
    wire N__4891;
    wire N__4890;
    wire N__4887;
    wire N__4884;
    wire N__4879;
    wire N__4872;
    wire N__4871;
    wire N__4870;
    wire N__4869;
    wire N__4866;
    wire N__4863;
    wire N__4858;
    wire N__4851;
    wire N__4850;
    wire N__4849;
    wire N__4848;
    wire N__4847;
    wire N__4846;
    wire N__4843;
    wire N__4840;
    wire N__4837;
    wire N__4834;
    wire N__4829;
    wire N__4818;
    wire N__4815;
    wire N__4812;
    wire N__4809;
    wire N__4806;
    wire N__4803;
    wire N__4800;
    wire N__4797;
    wire N__4794;
    wire N__4791;
    wire N__4788;
    wire N__4785;
    wire N__4782;
    wire N__4779;
    wire N__4776;
    wire N__4773;
    wire N__4770;
    wire N__4767;
    wire N__4764;
    wire N__4761;
    wire N__4758;
    wire N__4755;
    wire N__4752;
    wire N__4749;
    wire N__4746;
    wire N__4743;
    wire N__4740;
    wire N__4737;
    wire N__4734;
    wire N__4731;
    wire N__4728;
    wire N__4725;
    wire N__4724;
    wire N__4721;
    wire N__4718;
    wire N__4715;
    wire N__4712;
    wire N__4709;
    wire N__4706;
    wire N__4703;
    wire N__4700;
    wire N__4697;
    wire N__4694;
    wire N__4691;
    wire N__4688;
    wire N__4685;
    wire N__4682;
    wire N__4677;
    wire N__4674;
    wire N__4671;
    wire N__4668;
    wire N__4665;
    wire N__4662;
    wire N__4659;
    wire N__4656;
    wire N__4653;
    wire N__4652;
    wire N__4649;
    wire N__4648;
    wire N__4645;
    wire N__4642;
    wire N__4639;
    wire N__4636;
    wire N__4633;
    wire N__4630;
    wire N__4627;
    wire N__4624;
    wire N__4621;
    wire N__4618;
    wire N__4613;
    wire N__4608;
    wire N__4605;
    wire N__4602;
    wire N__4601;
    wire N__4598;
    wire N__4595;
    wire N__4590;
    wire N__4587;
    wire N__4584;
    wire N__4581;
    wire N__4578;
    wire N__4575;
    wire N__4572;
    wire N__4569;
    wire N__4568;
    wire N__4565;
    wire N__4562;
    wire N__4557;
    wire N__4554;
    wire N__4551;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4539;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4527;
    wire N__4524;
    wire N__4521;
    wire N__4518;
    wire N__4515;
    wire N__4512;
    wire N__4509;
    wire N__4506;
    wire N__4503;
    wire N__4500;
    wire N__4497;
    wire N__4494;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4486;
    wire N__4483;
    wire N__4480;
    wire N__4477;
    wire N__4474;
    wire N__4469;
    wire N__4466;
    wire N__4463;
    wire N__4458;
    wire N__4455;
    wire N__4452;
    wire N__4449;
    wire N__4446;
    wire N__4445;
    wire N__4442;
    wire N__4439;
    wire N__4434;
    wire N__4431;
    wire N__4428;
    wire N__4425;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4407;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4397;
    wire N__4394;
    wire N__4391;
    wire N__4388;
    wire N__4385;
    wire N__4382;
    wire N__4379;
    wire N__4376;
    wire N__4373;
    wire N__4370;
    wire N__4365;
    wire N__4362;
    wire N__4359;
    wire N__4356;
    wire N__4353;
    wire N__4350;
    wire N__4347;
    wire N__4344;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4323;
    wire N__4322;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4310;
    wire N__4309;
    wire N__4304;
    wire N__4301;
    wire N__4298;
    wire N__4295;
    wire N__4290;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4278;
    wire N__4277;
    wire N__4274;
    wire N__4271;
    wire N__4266;
    wire N__4265;
    wire N__4260;
    wire N__4257;
    wire N__4254;
    wire N__4251;
    wire N__4248;
    wire N__4245;
    wire N__4242;
    wire N__4241;
    wire N__4238;
    wire N__4233;
    wire N__4230;
    wire N__4227;
    wire N__4224;
    wire N__4221;
    wire N__4218;
    wire N__4215;
    wire N__4214;
    wire N__4213;
    wire N__4210;
    wire N__4205;
    wire N__4202;
    wire N__4197;
    wire N__4194;
    wire N__4193;
    wire N__4192;
    wire N__4187;
    wire N__4184;
    wire N__4179;
    wire N__4178;
    wire N__4177;
    wire N__4176;
    wire N__4175;
    wire N__4170;
    wire N__4167;
    wire N__4162;
    wire N__4155;
    wire N__4154;
    wire N__4151;
    wire N__4148;
    wire N__4143;
    wire N__4142;
    wire N__4139;
    wire N__4136;
    wire N__4131;
    wire N__4128;
    wire N__4125;
    wire N__4122;
    wire N__4119;
    wire N__4116;
    wire N__4113;
    wire N__4110;
    wire N__4107;
    wire N__4106;
    wire N__4105;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4086;
    wire N__4083;
    wire N__4080;
    wire N__4077;
    wire N__4074;
    wire N__4071;
    wire N__4068;
    wire N__4065;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4053;
    wire N__4050;
    wire N__4047;
    wire N__4044;
    wire N__4041;
    wire N__4038;
    wire N__4035;
    wire N__4032;
    wire N__4029;
    wire N__4026;
    wire N__4023;
    wire N__4020;
    wire N__4017;
    wire N__4014;
    wire N__4011;
    wire N__4008;
    wire N__4005;
    wire N__4002;
    wire N__3999;
    wire N__3996;
    wire N__3993;
    wire N__3990;
    wire N__3987;
    wire N__3984;
    wire N__3981;
    wire N__3978;
    wire N__3975;
    wire N__3972;
    wire N__3969;
    wire N__3966;
    wire N__3965;
    wire N__3962;
    wire N__3959;
    wire N__3956;
    wire N__3953;
    wire N__3950;
    wire N__3947;
    wire N__3944;
    wire N__3941;
    wire N__3938;
    wire N__3935;
    wire N__3932;
    wire N__3929;
    wire N__3924;
    wire N__3921;
    wire N__3918;
    wire N__3915;
    wire N__3912;
    wire N__3909;
    wire N__3906;
    wire N__3903;
    wire N__3900;
    wire N__3897;
    wire N__3894;
    wire N__3891;
    wire N__3888;
    wire N__3885;
    wire N__3882;
    wire N__3879;
    wire N__3876;
    wire N__3873;
    wire N__3870;
    wire N__3867;
    wire N__3864;
    wire N__3861;
    wire N__3858;
    wire N__3855;
    wire N__3852;
    wire N__3849;
    wire N__3846;
    wire N__3843;
    wire N__3840;
    wire N__3837;
    wire N__3834;
    wire N__3831;
    wire N__3828;
    wire N__3825;
    wire N__3822;
    wire N__3819;
    wire N__3816;
    wire N__3813;
    wire N__3812;
    wire N__3807;
    wire N__3804;
    wire N__3801;
    wire N__3798;
    wire N__3797;
    wire N__3794;
    wire N__3791;
    wire N__3786;
    wire N__3783;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire N__3771;
    wire N__3768;
    wire N__3765;
    wire N__3762;
    wire N__3759;
    wire N__3756;
    wire N__3753;
    wire N__3750;
    wire N__3749;
    wire N__3746;
    wire N__3743;
    wire N__3740;
    wire N__3737;
    wire N__3734;
    wire N__3731;
    wire N__3728;
    wire N__3725;
    wire N__3720;
    wire N__3717;
    wire N__3714;
    wire N__3711;
    wire N__3708;
    wire N__3705;
    wire N__3702;
    wire N__3699;
    wire N__3696;
    wire N__3693;
    wire N__3690;
    wire N__3687;
    wire N__3684;
    wire N__3681;
    wire N__3678;
    wire N__3675;
    wire N__3672;
    wire N__3669;
    wire N__3666;
    wire N__3663;
    wire N__3660;
    wire N__3657;
    wire N__3654;
    wire N__3651;
    wire N__3648;
    wire N__3645;
    wire N__3642;
    wire N__3639;
    wire N__3636;
    wire N__3633;
    wire N__3630;
    wire N__3627;
    wire N__3624;
    wire N__3621;
    wire N__3618;
    wire N__3615;
    wire N__3612;
    wire N__3609;
    wire N__3606;
    wire N__3605;
    wire N__3604;
    wire N__3601;
    wire N__3596;
    wire N__3591;
    wire N__3588;
    wire N__3585;
    wire N__3582;
    wire N__3579;
    wire N__3576;
    wire N__3573;
    wire N__3570;
    wire N__3567;
    wire N__3564;
    wire N__3563;
    wire N__3560;
    wire N__3557;
    wire N__3556;
    wire N__3553;
    wire N__3552;
    wire N__3549;
    wire N__3546;
    wire N__3543;
    wire N__3540;
    wire N__3537;
    wire N__3534;
    wire N__3529;
    wire N__3526;
    wire N__3523;
    wire N__3520;
    wire N__3517;
    wire N__3514;
    wire N__3511;
    wire N__3508;
    wire N__3505;
    wire N__3502;
    wire N__3497;
    wire N__3492;
    wire N__3489;
    wire N__3486;
    wire N__3483;
    wire N__3480;
    wire N__3477;
    wire N__3474;
    wire N__3471;
    wire N__3468;
    wire N__3467;
    wire N__3464;
    wire N__3461;
    wire N__3456;
    wire N__3453;
    wire N__3450;
    wire N__3447;
    wire N__3444;
    wire N__3441;
    wire N__3438;
    wire N__3435;
    wire N__3432;
    wire N__3429;
    wire N__3426;
    wire N__3423;
    wire N__3420;
    wire N__3417;
    wire N__3414;
    wire N__3411;
    wire N__3408;
    wire N__3405;
    wire N__3402;
    wire N__3399;
    wire N__3396;
    wire N__3393;
    wire N__3390;
    wire N__3387;
    wire N__3384;
    wire N__3381;
    wire N__3378;
    wire N__3375;
    wire N__3372;
    wire N__3369;
    wire N__3366;
    wire N__3363;
    wire N__3360;
    wire N__3357;
    wire N__3354;
    wire N__3351;
    wire N__3348;
    wire N__3345;
    wire N__3342;
    wire N__3339;
    wire N__3336;
    wire N__3333;
    wire N__3332;
    wire N__3329;
    wire N__3326;
    wire N__3323;
    wire N__3320;
    wire N__3317;
    wire N__3314;
    wire N__3311;
    wire N__3308;
    wire N__3305;
    wire N__3302;
    wire N__3297;
    wire N__3294;
    wire N__3291;
    wire N__3288;
    wire N__3285;
    wire N__3282;
    wire N__3279;
    wire N__3276;
    wire N__3273;
    wire N__3270;
    wire N__3267;
    wire N__3264;
    wire N__3261;
    wire N__3258;
    wire N__3257;
    wire N__3254;
    wire N__3251;
    wire N__3248;
    wire N__3245;
    wire N__3242;
    wire N__3239;
    wire N__3236;
    wire N__3233;
    wire N__3230;
    wire N__3227;
    wire N__3224;
    wire N__3221;
    wire N__3218;
    wire N__3213;
    wire N__3210;
    wire N__3207;
    wire N__3204;
    wire N__3201;
    wire N__3198;
    wire N__3195;
    wire N__3192;
    wire N__3189;
    wire N__3186;
    wire N__3183;
    wire N__3180;
    wire N__3177;
    wire N__3174;
    wire N__3171;
    wire N__3168;
    wire N__3167;
    wire N__3164;
    wire N__3161;
    wire N__3158;
    wire N__3155;
    wire N__3152;
    wire N__3149;
    wire N__3146;
    wire N__3143;
    wire N__3138;
    wire N__3135;
    wire N__3132;
    wire N__3129;
    wire N__3126;
    wire N__3123;
    wire N__3120;
    wire N__3117;
    wire N__3114;
    wire N__3111;
    wire N__3108;
    wire N__3105;
    wire N__3102;
    wire N__3099;
    wire N__3096;
    wire N__3093;
    wire N__3090;
    wire N__3087;
    wire N__3084;
    wire N__3081;
    wire N__3078;
    wire N__3075;
    wire N__3072;
    wire N__3069;
    wire N__3066;
    wire N__3063;
    wire N__3060;
    wire N__3057;
    wire N__3054;
    wire N__3051;
    wire N__3048;
    wire N__3045;
    wire N__3042;
    wire N__3039;
    wire N__3036;
    wire N__3033;
    wire N__3030;
    wire N__3027;
    wire N__3026;
    wire N__3023;
    wire N__3020;
    wire N__3017;
    wire N__3014;
    wire N__3011;
    wire N__3008;
    wire N__3005;
    wire N__3002;
    wire N__2999;
    wire N__2996;
    wire N__2993;
    wire N__2990;
    wire N__2987;
    wire N__2982;
    wire N__2979;
    wire N__2976;
    wire N__2973;
    wire N__2970;
    wire N__2967;
    wire N__2964;
    wire N__2961;
    wire N__2958;
    wire N__2955;
    wire N__2952;
    wire N__2949;
    wire N__2946;
    wire N__2943;
    wire N__2940;
    wire N__2937;
    wire N__2934;
    wire N__2931;
    wire N__2930;
    wire N__2927;
    wire N__2924;
    wire N__2921;
    wire N__2918;
    wire N__2915;
    wire N__2912;
    wire N__2907;
    wire N__2904;
    wire N__2901;
    wire N__2898;
    wire N__2895;
    wire N__2892;
    wire N__2889;
    wire N__2886;
    wire N__2883;
    wire N__2880;
    wire N__2877;
    wire N__2874;
    wire N__2871;
    wire N__2868;
    wire N__2865;
    wire N__2862;
    wire N__2861;
    wire N__2858;
    wire N__2855;
    wire N__2852;
    wire N__2849;
    wire N__2846;
    wire N__2843;
    wire N__2840;
    wire N__2837;
    wire N__2834;
    wire N__2831;
    wire N__2828;
    wire N__2823;
    wire N__2820;
    wire N__2817;
    wire N__2814;
    wire N__2811;
    wire N__2808;
    wire N__2805;
    wire N__2802;
    wire N__2799;
    wire N__2796;
    wire N__2793;
    wire N__2790;
    wire N__2787;
    wire N__2784;
    wire N__2781;
    wire N__2778;
    wire N__2775;
    wire N__2772;
    wire N__2769;
    wire N__2766;
    wire N__2763;
    wire N__2760;
    wire N__2757;
    wire N__2754;
    wire N__2751;
    wire N__2748;
    wire N__2745;
    wire N__2742;
    wire N__2739;
    wire N__2736;
    wire N__2733;
    wire N__2730;
    wire N__2727;
    wire N__2724;
    wire N__2721;
    wire N__2718;
    wire N__2715;
    wire N__2712;
    wire N__2709;
    wire N__2706;
    wire N__2703;
    wire N__2700;
    wire N__2697;
    wire N__2694;
    wire N__2691;
    wire N__2688;
    wire N__2685;
    wire N__2682;
    wire N__2679;
    wire N__2676;
    wire N__2673;
    wire N__2670;
    wire N__2667;
    wire N__2664;
    wire N__2661;
    wire N__2658;
    wire N__2655;
    wire GNDG0;
    wire VCCG0;
    wire TAn_in;
    wire RESETn_c_i;
    wire U111_CYCLE_SM_A_AMIGA_0_i_1;
    wire A_040_c_0;
    wire A_AMIGA_c_0;
    wire D_UM_040_in_2;
    wire D_LL_040_in_2;
    wire un1_D_UM_040_2;
    wire D_UU_040_in_4;
    wire D_LM_040_in_4;
    wire un1_D_UU_040_4;
    wire D_UM_040_in_4;
    wire D_LL_040_in_4;
    wire un1_D_UM_040_4;
    wire D_LL_AMIGA_in_1;
    wire un2_D_LL_AMIGA_1;
    wire CPUBGn_c_i_0;
    wire D_LL_AMIGA_in_5;
    wire un2_D_LL_AMIGA_5;
    wire D_LL_AMIGA_in_7;
    wire un2_D_LL_AMIGA_7;
    wire A_040_c_1;
    wire D_LM_AMIGA_in_5;
    wire N_108;
    wire D_LM_AMIGA_in_3;
    wire N_110;
    wire D_LM_AMIGA_in_2;
    wire N_111;
    wire D_UM_040_in_6;
    wire D_LL_040_in_6;
    wire un1_D_UM_040_6;
    wire D_UU_040_in_0;
    wire D_LM_040_in_0;
    wire un1_D_UU_040_0;
    wire D_UU_040_in_6;
    wire D_LM_040_in_6;
    wire un1_D_UU_040_6;
    wire D_LL_AMIGA_in_4;
    wire un2_D_LL_AMIGA_4;
    wire D_LL_AMIGA_in_2;
    wire un2_D_LL_AMIGA_2;
    wire D_LL_040_in_0;
    wire D_UM_040_in_0;
    wire un1_D_UM_040_0;
    wire D_LM_AMIGA_in_1;
    wire N_112;
    wire N_96;
    wire N_94_i;
    wire BBn_c;
    wire BUFDIR_c;
    wire GB_BUFFER_CLK40_THRU_CO;
    wire \U111_CYCLE_SM.N_141 ;
    wire \U111_CYCLE_SM.TS_ENZ0 ;
    wire \INVU111_CYCLE_SM.TS_OUTC_net ;
    wire D_LM_AMIGA_in_7;
    wire N_106;
    wire D_LM_AMIGA_in_6;
    wire N_107;
    wire D_UM_040_in_3;
    wire D_LL_040_in_3;
    wire un1_D_UM_040_3;
    wire D_LL_AMIGA_in_3;
    wire un2_D_LL_AMIGA_3;
    wire LBENn_c_i;
    wire D_LM_AMIGA_in_0;
    wire un2_D_LM_AMIGA_0;
    wire \U111_CYCLE_SM.A2_ENZ0 ;
    wire \U111_CYCLE_SM.N_179 ;
    wire \U111_CYCLE_SM.N_179_cascade_ ;
    wire \U111_CYCLE_SM.N_101_cascade_ ;
    wire \U111_CYCLE_SM.N_98 ;
    wire \U111_CYCLE_SM.N_10 ;
    wire \U111_CYCLE_SM.N_101 ;
    wire \U111_CYCLE_SM.N_12_i_1_cascade_ ;
    wire \U111_CYCLE_SM.N_55 ;
    wire \U111_CYCLE_SM.BURST_COUNTZ0Z_1 ;
    wire SIZ_c_0;
    wire SIZ_c_1;
    wire \U111_CYCLE_SM.BURST_COUNTZ0Z_0 ;
    wire \U111_CYCLE_SM.LW_TRANSZ0 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ;
    wire PORTSIZE_c;
    wire TS_CPUn_in;
    wire D_LM_AMIGA_in_4;
    wire N_109;
    wire D_UU_040_in_2;
    wire D_LM_040_in_2;
    wire un1_D_UU_040_2;
    wire D_UU_AMIGA_in_2;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ;
    wire N_118;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ;
    wire D_UU_AMIGA_in_4;
    wire N_116;
    wire D_UU_AMIGA_in_7;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ;
    wire N_113;
    wire D_LM_040_in_3;
    wire D_UU_040_in_3;
    wire un1_D_UU_040_3;
    wire D_UU_AMIGA_in_5;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ;
    wire N_115;
    wire \U111_CYCLE_SM.CYCLE_STATE_srsts_i_i_o2_0_5_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ;
    wire \U111_CYCLE_SM.PORT_MISMATCHZ0 ;
    wire \U111_CYCLE_SM.BURSTZ0 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ;
    wire \U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_a3_2_0_0_cascade_ ;
    wire \U111_CYCLE_SM.N_133 ;
    wire \U111_CYCLE_SM.N_131 ;
    wire \U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_2_0_cascade_ ;
    wire \U111_CYCLE_SM.TS_DELAYZ0 ;
    wire \U111_CYCLE_SM.un4_TS_OUT_i_0_cascade_ ;
    wire TACKn_in;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ;
    wire \U111_CYCLE_SM.N_99_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ;
    wire \U111_CYCLE_SM.N_51 ;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ;
    wire D_LM_040_in_1;
    wire D_UU_040_in_1;
    wire un1_D_UU_040_1;
    wire TS_OUT;
    wire TSnz;
    wire D_LM_040_in_7;
    wire D_UU_040_in_7;
    wire un1_D_UU_040_7;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ;
    wire D_UU_AMIGA_in_6;
    wire N_114;
    wire CONSTANT_ONE_NET;
    wire BGn_c;
    wire \U111_CYCLE_SM.CYCLE_ENZ0 ;
    wire \U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0 ;
    wire U111_CYCLE_SM_OFFBOARD_EN_0;
    wire \U111_CYCLE_SM.un4_TS_OUT_i_0 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ;
    wire RESETn_c_i_g;
    wire RESETn_c;
    wire \U111_CYCLE_SM.N_99 ;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81_cascade_ ;
    wire \U111_CYCLE_SM.N_99_i ;
    wire D_UM_040_in_1;
    wire D_LL_040_in_1;
    wire un1_D_UM_040_1;
    wire D_UU_AMIGA_in_1;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ;
    wire N_119;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ;
    wire D_UM_AMIGA_in_4;
    wire un1_D_UM_AMIGA_4;
    wire CLK80;
    wire GB_BUFFER_CLK80_THRU_CO;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ;
    wire D_UU_AMIGA_in_0;
    wire un1_D_UU_AMIGA_0;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ;
    wire D_UU_AMIGA_in_3;
    wire N_117;
    wire D_LL_AMIGA_in_0;
    wire un2_D_LL_AMIGA_0;
    wire TBIn_c;
    wire U111_CYCLE_SM_TBI_CPUn_0_i;
    wire D_LL_AMIGA_in_6;
    wire un2_D_LL_AMIGA_6;
    wire un1_D_UM_AMIGA_2;
    wire un1_D_UM_AMIGA_0;
    wire TEAn_c;
    wire U111_CYCLE_SM_TEA_CPUn_0_i;
    wire D_UM_AMIGA_in_2;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ;
    wire D_UM_AMIGA_in_0;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ;
    wire CLK40;
    wire \U111_CYCLE_SM.N_99_i_0 ;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81 ;
    wire D_UM_AMIGA_in_1;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ;
    wire un1_D_UM_AMIGA_1;
    wire \U111_CYCLE_SM.TA_DISZ0 ;
    wire N_64;
    wire TCIn_c;
    wire LBENn_c;
    wire U111_CYCLE_SM_TCI_CPUn_0_i;
    wire D_UM_AMIGA_in_3;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ;
    wire un1_D_UM_AMIGA_3;
    wire D_LL_040_in_7;
    wire D_UM_040_in_7;
    wire un1_D_UM_040_7;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ;
    wire D_UM_AMIGA_in_7;
    wire un1_D_UM_AMIGA_7;
    wire D_LM_040_in_5;
    wire D_UU_040_in_5;
    wire un1_D_UU_040_5;
    wire D_UM_040_in_5;
    wire D_LL_040_in_5;
    wire \U111_CYCLE_SM.FLIP_WORDZ0 ;
    wire un1_D_UM_040_5;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ;
    wire D_UM_AMIGA_in_5;
    wire un1_D_UM_AMIGA_5;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ;
    wire CPUBGn_c;
    wire RnW_c;
    wire N_60_i;
    wire \U111_CYCLE_SM.LATCH_ENZ0 ;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ;
    wire D_UM_AMIGA_in_6;
    wire un1_D_UM_AMIGA_6;
    wire _gnd_net_;

    defparam pll_pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll_pll.TEST_MODE=1'b0;
    defparam pll_pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll_pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll_pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll_pll.FILTER_RANGE=3'b011;
    defparam pll_pll.FEEDBACK_PATH="SIMPLE";
    defparam pll_pll.FDA_RELATIVE=4'b0000;
    defparam pll_pll.FDA_FEEDBACK=4'b0000;
    defparam pll_pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll_pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll_pll.DIVR=4'b0000;
    defparam pll_pll.DIVQ=3'b011;
    defparam pll_pll.DIVF=7'b0001111;
    defparam pll_pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40_2F pll_pll (
            .SCLK(),
            .PLLOUTGLOBALA(CLK80),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALB(CLK40),
            .SDI(),
            .PLLOUTCOREA(),
            .BYPASS(),
            .RESETB(N__5553),
            .PLLOUTCOREB(),
            .LOCK(),
            .SDO(),
            .EXTFEEDBACK(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__9524));
    IO_PAD pll_iopad (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__9524),
            .PACKAGEPIN(CLK40_IN));
    IO_PAD LBENn_ibuf_iopad (
            .OE(N__9508),
            .DIN(N__9507),
            .DOUT(N__9506),
            .PACKAGEPIN(LBENn));
    defparam LBENn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam LBENn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO LBENn_ibuf_preio (
            .PADOEN(N__9508),
            .PADOUT(N__9507),
            .PADIN(N__9506),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(LBENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_obuft_iopad (
            .OE(N__9499),
            .DIN(N__9498),
            .DOUT(N__9497),
            .PACKAGEPIN(TSn));
    defparam TSn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TSn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TSn_obuft_preio (
            .PADOEN(N__9499),
            .PADOUT(N__9498),
            .PADIN(N__9497),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2763),
            .DIN0(),
            .DOUT0(N__5760),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_3_iopad (
            .OE(N__9490),
            .DIN(N__9489),
            .DOUT(N__9488),
            .PACKAGEPIN(D_UM_040[3]));
    defparam D_UM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_3_preio (
            .PADOEN(N__9490),
            .PADOUT(N__9489),
            .PADIN(N__9488),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7637),
            .DIN0(D_UM_040_in_3),
            .DOUT0(N__8556),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TAn_iobuf_iopad (
            .OE(N__9481),
            .DIN(N__9480),
            .DOUT(N__9479),
            .PACKAGEPIN(TAn));
    defparam TAn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TAn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TAn_iobuf_preio (
            .PADOEN(N__9481),
            .PADOUT(N__9480),
            .PADIN(N__9479),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6918),
            .DIN0(TAn_in),
            .DOUT0(N__5205),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_1_iopad (
            .OE(N__9472),
            .DIN(N__9471),
            .DOUT(N__9470),
            .PACKAGEPIN(D_LL_AMIGA[1]));
    defparam D_LL_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_1_preio (
            .PADOEN(N__9472),
            .PADOUT(N__9471),
            .PADIN(N__9470),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5435),
            .DIN0(D_LL_AMIGA_in_1),
            .DOUT0(N__6099),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_5_iopad (
            .OE(N__9463),
            .DIN(N__9462),
            .DOUT(N__9461),
            .PACKAGEPIN(D_UU_AMIGA[5]));
    defparam D_UU_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_5_preio (
            .PADOEN(N__9463),
            .PADOUT(N__9462),
            .PADIN(N__9461),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5475),
            .DIN0(D_UU_AMIGA_in_5),
            .DOUT0(N__8304),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_6_iopad (
            .OE(N__9454),
            .DIN(N__9453),
            .DOUT(N__9452),
            .PACKAGEPIN(D_UU_040[6]));
    defparam D_UU_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_6_preio (
            .PADOEN(N__9454),
            .PADOUT(N__9453),
            .PADIN(N__9452),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7646),
            .DIN0(D_UU_040_in_6),
            .DOUT0(N__5574),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CPUBGn_obuf_iopad (
            .OE(N__9445),
            .DIN(N__9444),
            .DOUT(N__9443),
            .PACKAGEPIN(CPUBGn));
    defparam CPUBGn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CPUBGn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CPUBGn_obuf_preio (
            .PADOEN(N__9445),
            .PADOUT(N__9444),
            .PADIN(N__9443),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7824),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_7_iopad (
            .OE(N__9436),
            .DIN(N__9435),
            .DOUT(N__9434),
            .PACKAGEPIN(D_LL_040[7]));
    defparam D_LL_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_7_preio (
            .PADOEN(N__9436),
            .PADOUT(N__9435),
            .PADIN(N__9434),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7528),
            .DIN0(D_LL_040_in_7),
            .DOUT0(N__2706),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_4_iopad (
            .OE(N__9427),
            .DIN(N__9426),
            .DOUT(N__9425),
            .PACKAGEPIN(D_LL_AMIGA[4]));
    defparam D_LL_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_4_preio (
            .PADOEN(N__9427),
            .PADOUT(N__9426),
            .PADIN(N__9425),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5434),
            .DIN0(D_LL_AMIGA_in_4),
            .DOUT0(N__2865),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_3_iopad (
            .OE(N__9418),
            .DIN(N__9417),
            .DOUT(N__9416),
            .PACKAGEPIN(D_UM_AMIGA[3]));
    defparam D_UM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_3_preio (
            .PADOEN(N__9418),
            .PADOUT(N__9417),
            .PADIN(N__9416),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5431),
            .DIN0(D_UM_AMIGA_in_3),
            .DOUT0(N__3921),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_3_iopad (
            .OE(N__9409),
            .DIN(N__9408),
            .DOUT(N__9407),
            .PACKAGEPIN(D_UU_040[3]));
    defparam D_UU_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_3_preio (
            .PADOEN(N__9409),
            .PADOUT(N__9408),
            .PADIN(N__9407),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7480),
            .DIN0(D_UU_040_in_3),
            .DOUT0(N__6678),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TEA_CPUn_obuf_iopad (
            .OE(N__9400),
            .DIN(N__9399),
            .DOUT(N__9398),
            .PACKAGEPIN(TEA_CPUn));
    defparam TEA_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TEA_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TEA_CPUn_obuf_preio (
            .PADOEN(N__9400),
            .PADOUT(N__9399),
            .PADIN(N__9398),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6432),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_1_iopad (
            .OE(N__9391),
            .DIN(N__9390),
            .DOUT(N__9389),
            .PACKAGEPIN(A_040[1]));
    defparam A_040_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_1_preio (
            .PADOEN(N__9391),
            .PADOUT(N__9390),
            .PADIN(N__9389),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_3_iopad (
            .OE(N__9382),
            .DIN(N__9381),
            .DOUT(N__9380),
            .PACKAGEPIN(D_LM_AMIGA[3]));
    defparam D_LM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_3_preio (
            .PADOEN(N__9382),
            .PADOUT(N__9381),
            .PADIN(N__9380),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5266),
            .DIN0(D_LM_AMIGA_in_3),
            .DOUT0(N__4413),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_0_iopad (
            .OE(N__9373),
            .DIN(N__9372),
            .DOUT(N__9371),
            .PACKAGEPIN(D_LM_040[0]));
    defparam D_LM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_0_preio (
            .PADOEN(N__9373),
            .PADOUT(N__9372),
            .PADIN(N__9371),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7529),
            .DIN0(D_LM_040_in_0),
            .DOUT0(N__3834),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_6_iopad (
            .OE(N__9364),
            .DIN(N__9363),
            .DOUT(N__9362),
            .PACKAGEPIN(D_UM_AMIGA[6]));
    defparam D_UM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_6_preio (
            .PADOEN(N__9364),
            .PADOUT(N__9363),
            .PADIN(N__9362),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5457),
            .DIN0(D_UM_AMIGA_in_6),
            .DOUT0(N__3294),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_4_iopad (
            .OE(N__9355),
            .DIN(N__9354),
            .DOUT(N__9353),
            .PACKAGEPIN(D_LM_AMIGA[4]));
    defparam D_LM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_4_preio (
            .PADOEN(N__9355),
            .PADOUT(N__9354),
            .PADIN(N__9353),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5326),
            .DIN0(D_LM_AMIGA_in_4),
            .DOUT0(N__2940),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_1_iopad (
            .OE(N__9346),
            .DIN(N__9345),
            .DOUT(N__9344),
            .PACKAGEPIN(A_AMIGA[1]));
    defparam A_AMIGA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_1_preio (
            .PADOEN(N__9346),
            .PADOUT(N__9345),
            .PADIN(N__9344),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3078),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_7_iopad (
            .OE(N__9337),
            .DIN(N__9336),
            .DOUT(N__9335),
            .PACKAGEPIN(D_LM_040[7]));
    defparam D_LM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_7_preio (
            .PADOEN(N__9337),
            .PADOUT(N__9336),
            .PADIN(N__9335),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7600),
            .DIN0(D_LM_040_in_7),
            .DOUT0(N__4035),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_4_iopad (
            .OE(N__9328),
            .DIN(N__9327),
            .DOUT(N__9326),
            .PACKAGEPIN(D_UM_040[4]));
    defparam D_UM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_4_preio (
            .PADOEN(N__9328),
            .PADOUT(N__9327),
            .PADIN(N__9326),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7481),
            .DIN0(D_UM_040_in_4),
            .DOUT0(N__5892),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_obuf_iopad (
            .OE(N__9319),
            .DIN(N__9318),
            .DOUT(N__9317),
            .PACKAGEPIN(CLK40B));
    defparam CLK40B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_obuf_preio (
            .PADOEN(N__9319),
            .PADOUT(N__9318),
            .PADIN(N__9317),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3552),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_0_iopad (
            .OE(N__9310),
            .DIN(N__9309),
            .DOUT(N__9308),
            .PACKAGEPIN(D_UU_AMIGA[0]));
    defparam D_UU_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_0_preio (
            .PADOEN(N__9310),
            .PADOUT(N__9309),
            .PADIN(N__9308),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5465),
            .DIN0(D_UU_AMIGA_in_0),
            .DOUT0(N__3210),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_1_iopad (
            .OE(N__9301),
            .DIN(N__9300),
            .DOUT(N__9299),
            .PACKAGEPIN(D_UM_040[1]));
    defparam D_UM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_1_preio (
            .PADOEN(N__9301),
            .PADOUT(N__9300),
            .PADIN(N__9299),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7479),
            .DIN0(D_UM_040_in_1),
            .DOUT0(N__6966),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_ibuf_iopad (
            .OE(N__9292),
            .DIN(N__9291),
            .DOUT(N__9290),
            .PACKAGEPIN(TBIn));
    defparam TBIn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TBIn_ibuf_preio (
            .PADOEN(N__9292),
            .PADOUT(N__9291),
            .PADIN(N__9290),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TBIn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_4_iopad (
            .OE(N__9283),
            .DIN(N__9282),
            .DOUT(N__9281),
            .PACKAGEPIN(D_LL_040[4]));
    defparam D_LL_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_4_preio (
            .PADOEN(N__9283),
            .PADOUT(N__9282),
            .PADIN(N__9281),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7633),
            .DIN0(D_LL_040_in_4),
            .DOUT0(N__3099),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_7_iopad (
            .OE(N__9274),
            .DIN(N__9273),
            .DOUT(N__9272),
            .PACKAGEPIN(D_LL_AMIGA[7]));
    defparam D_LL_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_7_preio (
            .PADOEN(N__9274),
            .PADOUT(N__9273),
            .PADIN(N__9272),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5395),
            .DIN0(D_LL_AMIGA_in_7),
            .DOUT0(N__8535),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_7_iopad (
            .OE(N__9265),
            .DIN(N__9264),
            .DOUT(N__9263),
            .PACKAGEPIN(D_UU_AMIGA[7]));
    defparam D_UU_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_7_preio (
            .PADOEN(N__9265),
            .PADOUT(N__9264),
            .PADIN(N__9263),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5467),
            .DIN0(D_UU_AMIGA_in_7),
            .DOUT0(N__5646),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFDIR_obuf_iopad (
            .OE(N__9256),
            .DIN(N__9255),
            .DOUT(N__9254),
            .PACKAGEPIN(BUFDIR));
    defparam BUFDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFDIR_obuf_preio (
            .PADOEN(N__9256),
            .PADOUT(N__9255),
            .PADIN(N__9254),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3582),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_4_iopad (
            .OE(N__9247),
            .DIN(N__9246),
            .DOUT(N__9245),
            .PACKAGEPIN(D_UU_040[4]));
    defparam D_UU_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_4_preio (
            .PADOEN(N__9247),
            .PADOUT(N__9246),
            .PADIN(N__9245),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7614),
            .DIN0(D_UU_040_in_4),
            .DOUT0(N__4515),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__9238),
            .DIN(N__9237),
            .DOUT(N__9236),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__9238),
            .PADOUT(N__9237),
            .PADIN(N__9236),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_1_iopad (
            .OE(N__9229),
            .DIN(N__9228),
            .DOUT(N__9227),
            .PACKAGEPIN(D_LL_040[1]));
    defparam D_LL_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_1_preio (
            .PADOEN(N__9229),
            .PADOUT(N__9228),
            .PADIN(N__9227),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7632),
            .DIN0(D_LL_040_in_1),
            .DOUT0(N__2787),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_5_iopad (
            .OE(N__9220),
            .DIN(N__9219),
            .DOUT(N__9218),
            .PACKAGEPIN(D_UM_AMIGA[5]));
    defparam D_UM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_5_preio (
            .PADOEN(N__9220),
            .PADOUT(N__9219),
            .PADIN(N__9218),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5466),
            .DIN0(D_UM_AMIGA_in_5),
            .DOUT0(N__7980),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_1_iopad (
            .OE(N__9211),
            .DIN(N__9210),
            .DOUT(N__9209),
            .PACKAGEPIN(D_UU_040[1]));
    defparam D_UU_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_1_preio (
            .PADOEN(N__9211),
            .PADOUT(N__9210),
            .PADIN(N__9209),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7653),
            .DIN0(D_UU_040_in_1),
            .DOUT0(N__5976),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_1_iopad (
            .OE(N__9202),
            .DIN(N__9201),
            .DOUT(N__9200),
            .PACKAGEPIN(D_LM_AMIGA[1]));
    defparam D_LM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_1_preio (
            .PADOEN(N__9202),
            .PADOUT(N__9201),
            .PADIN(N__9200),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5323),
            .DIN0(D_LM_AMIGA_in_1),
            .DOUT0(N__5019),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_2_iopad (
            .OE(N__9193),
            .DIN(N__9192),
            .DOUT(N__9191),
            .PACKAGEPIN(D_LM_040[2]));
    defparam D_LM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_2_preio (
            .PADOEN(N__9193),
            .PADOUT(N__9192),
            .PADIN(N__9191),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7495),
            .DIN0(D_LM_040_in_2),
            .DOUT0(N__3375),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__9184),
            .DIN(N__9183),
            .DOUT(N__9182),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__9184),
            .PADOUT(N__9183),
            .PADIN(N__9182),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3861),
            .DIN0(TACKn_in),
            .DOUT0(N__2685),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_2_iopad (
            .OE(N__9175),
            .DIN(N__9174),
            .DOUT(N__9173),
            .PACKAGEPIN(D_UM_040[2]));
    defparam D_UM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_2_preio (
            .PADOEN(N__9175),
            .PADOUT(N__9174),
            .PADIN(N__9173),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7558),
            .DIN0(D_UM_040_in_2),
            .DOUT0(N__6537),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMB_obuf_iopad (
            .OE(N__9166),
            .DIN(N__9165),
            .DOUT(N__9164),
            .PACKAGEPIN(CLKRAMB));
    defparam CLKRAMB_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMB_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMB_obuf_preio (
            .PADOEN(N__9166),
            .PADOUT(N__9165),
            .PADIN(N__9164),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5856),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_2_iopad (
            .OE(N__9157),
            .DIN(N__9156),
            .DOUT(N__9155),
            .PACKAGEPIN(D_LL_AMIGA[2]));
    defparam D_LL_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_2_preio (
            .PADOEN(N__9157),
            .PADOUT(N__9156),
            .PADIN(N__9155),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5285),
            .DIN0(D_LL_AMIGA_in_2),
            .DOUT0(N__3027),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_2_iopad (
            .OE(N__9148),
            .DIN(N__9147),
            .DOUT(N__9146),
            .PACKAGEPIN(D_UU_AMIGA[2]));
    defparam D_UU_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_2_preio (
            .PADOEN(N__9148),
            .PADOUT(N__9147),
            .PADIN(N__9146),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5464),
            .DIN0(D_UU_AMIGA_in_2),
            .DOUT0(N__4677),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TEAn_ibuf_iopad (
            .OE(N__9139),
            .DIN(N__9138),
            .DOUT(N__9137),
            .PACKAGEPIN(TEAn));
    defparam TEAn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TEAn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TEAn_ibuf_preio (
            .PADOEN(N__9139),
            .PADOUT(N__9138),
            .PADIN(N__9137),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TEAn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__9130),
            .DIN(N__9129),
            .DOUT(N__9128),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__9130),
            .PADOUT(N__9129),
            .PADIN(N__9128),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3624),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_6_iopad (
            .OE(N__9121),
            .DIN(N__9120),
            .DOUT(N__9119),
            .PACKAGEPIN(D_LL_040[6]));
    defparam D_LL_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_6_preio (
            .PADOEN(N__9121),
            .PADOUT(N__9120),
            .PADIN(N__9119),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7630),
            .DIN0(D_LL_040_in_6),
            .DOUT0(N__6558),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_5_iopad (
            .OE(N__9112),
            .DIN(N__9111),
            .DOUT(N__9110),
            .PACKAGEPIN(D_LL_AMIGA[5]));
    defparam D_LL_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_5_preio (
            .PADOEN(N__9112),
            .PADOUT(N__9111),
            .PADIN(N__9110),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5398),
            .DIN0(D_LL_AMIGA_in_5),
            .DOUT0(N__8268),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_0_iopad (
            .OE(N__9103),
            .DIN(N__9102),
            .DOUT(N__9101),
            .PACKAGEPIN(D_UM_AMIGA[0]));
    defparam D_UM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_0_preio (
            .PADOEN(N__9103),
            .PADOUT(N__9102),
            .PADIN(N__9101),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5325),
            .DIN0(D_UM_AMIGA_in_0),
            .DOUT0(N__3693),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_2_iopad (
            .OE(N__9094),
            .DIN(N__9093),
            .DOUT(N__9092),
            .PACKAGEPIN(D_UU_040[2]));
    defparam D_UU_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_2_preio (
            .PADOEN(N__9094),
            .PADOUT(N__9093),
            .PADIN(N__9092),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7527),
            .DIN0(D_UU_040_in_2),
            .DOUT0(N__4590),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_2_iopad (
            .OE(N__9085),
            .DIN(N__9084),
            .DOUT(N__9083),
            .PACKAGEPIN(D_LM_AMIGA[2]));
    defparam D_LM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_2_preio (
            .PADOEN(N__9085),
            .PADOUT(N__9084),
            .PADIN(N__9083),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5324),
            .DIN0(D_LM_AMIGA_in_2),
            .DOUT0(N__4725),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TS_CPUn_iobuf_iopad (
            .OE(N__9076),
            .DIN(N__9075),
            .DOUT(N__9074),
            .PACKAGEPIN(TS_CPUn));
    defparam TS_CPUn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TS_CPUn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TS_CPUn_iobuf_preio (
            .PADOEN(N__9076),
            .PADOUT(N__9075),
            .PADIN(N__9074),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7820),
            .DIN0(TS_CPUn_in),
            .DOUT0(N__5724),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK80_CPU_obuf_iopad (
            .OE(N__9067),
            .DIN(N__9066),
            .DOUT(N__9065),
            .PACKAGEPIN(CLK80_CPU));
    defparam CLK80_CPU_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK80_CPU_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK80_CPU_obuf_preio (
            .PADOEN(N__9067),
            .PADOUT(N__9066),
            .PADIN(N__9065),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5855),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_3_iopad (
            .OE(N__9058),
            .DIN(N__9057),
            .DOUT(N__9056),
            .PACKAGEPIN(D_LL_040[3]));
    defparam D_LL_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_3_preio (
            .PADOEN(N__9058),
            .PADOUT(N__9057),
            .PADIN(N__9056),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7634),
            .DIN0(D_LL_040_in_3),
            .DOUT0(N__3885),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_1_iopad (
            .OE(N__9049),
            .DIN(N__9048),
            .DOUT(N__9047),
            .PACKAGEPIN(D_LM_040[1]));
    defparam D_LM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_1_preio (
            .PADOEN(N__9049),
            .PADOUT(N__9048),
            .PADIN(N__9047),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7494),
            .DIN0(D_LM_040_in_1),
            .DOUT0(N__3663),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_7_iopad (
            .OE(N__9040),
            .DIN(N__9039),
            .DOUT(N__9038),
            .PACKAGEPIN(D_UM_AMIGA[7]));
    defparam D_UM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_7_preio (
            .PADOEN(N__9040),
            .PADOUT(N__9039),
            .PADIN(N__9038),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5432),
            .DIN0(D_UM_AMIGA_in_7),
            .DOUT0(N__8463),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_7_iopad (
            .OE(N__9031),
            .DIN(N__9030),
            .DOUT(N__9029),
            .PACKAGEPIN(D_LM_AMIGA[7]));
    defparam D_LM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_7_preio (
            .PADOEN(N__9031),
            .PADOUT(N__9030),
            .PADIN(N__9029),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5372),
            .DIN0(D_LM_AMIGA_in_7),
            .DOUT0(N__5706),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORTSIZE_ibuf_iopad (
            .OE(N__9022),
            .DIN(N__9021),
            .DOUT(N__9020),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO PORTSIZE_ibuf_preio (
            .PADOEN(N__9022),
            .PADOUT(N__9021),
            .PADIN(N__9020),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(PORTSIZE_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_0_iopad (
            .OE(N__9013),
            .DIN(N__9012),
            .DOUT(N__9011),
            .PACKAGEPIN(A_AMIGA[0]));
    defparam A_AMIGA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_0_preio (
            .PADOEN(N__9013),
            .PADOUT(N__9012),
            .PADIN(N__9011),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3054),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_4_iopad (
            .OE(N__9004),
            .DIN(N__9003),
            .DOUT(N__9002),
            .PACKAGEPIN(D_LM_040[4]));
    defparam D_LM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_4_preio (
            .PADOEN(N__9004),
            .PADOUT(N__9003),
            .PADIN(N__9002),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7610),
            .DIN0(D_LM_040_in_4),
            .DOUT0(N__4764),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_7_iopad (
            .OE(N__8995),
            .DIN(N__8994),
            .DOUT(N__8993),
            .PACKAGEPIN(D_UM_040[7]));
    defparam D_UM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_7_preio (
            .PADOEN(N__8995),
            .PADOUT(N__8994),
            .PADIN(N__8993),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7636),
            .DIN0(D_UM_040_in_7),
            .DOUT0(N__8382),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__8986),
            .DIN(N__8985),
            .DOUT(N__8984),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__8986),
            .PADOUT(N__8985),
            .PADIN(N__8984),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_1_iopad (
            .OE(N__8977),
            .DIN(N__8976),
            .DOUT(N__8975),
            .PACKAGEPIN(D_UU_AMIGA[1]));
    defparam D_UU_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_1_preio (
            .PADOEN(N__8977),
            .PADOUT(N__8976),
            .PADIN(N__8975),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5430),
            .DIN0(D_UU_AMIGA_in_1),
            .DOUT0(N__4968),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_obuf_iopad (
            .OE(N__8968),
            .DIN(N__8967),
            .DOUT(N__8966),
            .PACKAGEPIN(CLK40C));
    defparam CLK40C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_obuf_preio (
            .PADOEN(N__8968),
            .PADOUT(N__8967),
            .PADIN(N__8966),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3556),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_0_iopad (
            .OE(N__8959),
            .DIN(N__8958),
            .DOUT(N__8957),
            .PACKAGEPIN(D_UM_040[0]));
    defparam D_UM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_0_preio (
            .PADOEN(N__8959),
            .PADOUT(N__8958),
            .PADIN(N__8957),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7559),
            .DIN0(D_UM_040_in_0),
            .DOUT0(N__6525),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_0_iopad (
            .OE(N__8950),
            .DIN(N__8949),
            .DOUT(N__8948),
            .PACKAGEPIN(D_LL_AMIGA[0]));
    defparam D_LL_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_0_preio (
            .PADOEN(N__8950),
            .PADOUT(N__8949),
            .PADIN(N__8948),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5462),
            .DIN0(D_LL_AMIGA_in_0),
            .DOUT0(N__3753),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_4_iopad (
            .OE(N__8941),
            .DIN(N__8940),
            .DOUT(N__8939),
            .PACKAGEPIN(D_UU_AMIGA[4]));
    defparam D_UU_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_4_preio (
            .PADOEN(N__8941),
            .PADOUT(N__8940),
            .PADIN(N__8939),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5463),
            .DIN0(D_UU_AMIGA_in_4),
            .DOUT0(N__2901),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_7_iopad (
            .OE(N__8932),
            .DIN(N__8931),
            .DOUT(N__8930),
            .PACKAGEPIN(D_UU_040[7]));
    defparam D_UU_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_7_preio (
            .PADOEN(N__8932),
            .PADOUT(N__8931),
            .PADIN(N__8930),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7645),
            .DIN0(D_UU_040_in_7),
            .DOUT0(N__4434),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__8923),
            .DIN(N__8922),
            .DOUT(N__8921),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__8923),
            .PADOUT(N__8922),
            .PADIN(N__8921),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BGn_ibuf_iopad (
            .OE(N__8914),
            .DIN(N__8913),
            .DOUT(N__8912),
            .PACKAGEPIN(BGn));
    defparam BGn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BGn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BGn_ibuf_preio (
            .PADOEN(N__8914),
            .PADOUT(N__8913),
            .PADIN(N__8912),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(BGn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_0_iopad (
            .OE(N__8905),
            .DIN(N__8904),
            .DOUT(N__8903),
            .PACKAGEPIN(D_LL_040[0]));
    defparam D_LL_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_0_preio (
            .PADOEN(N__8905),
            .PADOUT(N__8904),
            .PADIN(N__8903),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7635),
            .DIN0(D_LL_040_in_0),
            .DOUT0(N__6639),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_2_iopad (
            .OE(N__8896),
            .DIN(N__8895),
            .DOUT(N__8894),
            .PACKAGEPIN(D_UM_AMIGA[2]));
    defparam D_UM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_2_preio (
            .PADOEN(N__8896),
            .PADOUT(N__8895),
            .PADIN(N__8894),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5327),
            .DIN0(D_UM_AMIGA_in_2),
            .DOUT0(N__2982),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_0_iopad (
            .OE(N__8887),
            .DIN(N__8886),
            .DOUT(N__8885),
            .PACKAGEPIN(D_UU_040[0]));
    defparam D_UU_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_0_preio (
            .PADOEN(N__8887),
            .PADOUT(N__8886),
            .PADIN(N__8885),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7644),
            .DIN0(D_UU_040_in_0),
            .DOUT0(N__6768),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_ibuf_iopad (
            .OE(N__8878),
            .DIN(N__8877),
            .DOUT(N__8876),
            .PACKAGEPIN(TCIn));
    defparam TCIn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TCIn_ibuf_preio (
            .PADOEN(N__8878),
            .PADOUT(N__8877),
            .PADIN(N__8876),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TCIn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_0_iopad (
            .OE(N__8869),
            .DIN(N__8868),
            .DOUT(N__8867),
            .PACKAGEPIN(A_040[0]));
    defparam A_040_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_0_preio (
            .PADOEN(N__8869),
            .PADOUT(N__8868),
            .PADIN(N__8867),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_0_iopad (
            .OE(N__8860),
            .DIN(N__8859),
            .DOUT(N__8858),
            .PACKAGEPIN(D_LM_AMIGA[0]));
    defparam D_LM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_0_preio (
            .PADOEN(N__8860),
            .PADOUT(N__8859),
            .PADIN(N__8858),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5396),
            .DIN0(D_LM_AMIGA_in_0),
            .DOUT0(N__3258),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBI_CPUn_obuf_iopad (
            .OE(N__8851),
            .DIN(N__8850),
            .DOUT(N__8849),
            .PACKAGEPIN(TBI_CPUn));
    defparam TBI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TBI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TBI_CPUn_obuf_preio (
            .PADOEN(N__8851),
            .PADOUT(N__8850),
            .PADIN(N__8849),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6588),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40A_obuf_iopad (
            .OE(N__8842),
            .DIN(N__8841),
            .DOUT(N__8840),
            .PACKAGEPIN(CLK40A));
    defparam CLK40A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40A_obuf_preio (
            .PADOEN(N__8842),
            .PADOUT(N__8841),
            .PADIN(N__8840),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3563),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_3_iopad (
            .OE(N__8833),
            .DIN(N__8832),
            .DOUT(N__8831),
            .PACKAGEPIN(D_LM_040[3]));
    defparam D_LM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_3_preio (
            .PADOEN(N__8833),
            .PADOUT(N__8832),
            .PADIN(N__8831),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7654),
            .DIN0(D_LM_040_in_3),
            .DOUT0(N__3411),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_5_iopad (
            .OE(N__8824),
            .DIN(N__8823),
            .DOUT(N__8822),
            .PACKAGEPIN(D_LM_AMIGA[5]));
    defparam D_LM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_5_preio (
            .PADOEN(N__8824),
            .PADOUT(N__8823),
            .PADIN(N__8822),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5370),
            .DIN0(D_LM_AMIGA_in_5),
            .DOUT0(N__8361),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_6_iopad (
            .OE(N__8815),
            .DIN(N__8814),
            .DOUT(N__8813),
            .PACKAGEPIN(D_LM_040[6]));
    defparam D_LM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_6_preio (
            .PADOEN(N__8815),
            .PADOUT(N__8814),
            .PADIN(N__8813),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7547),
            .DIN0(D_LM_040_in_6),
            .DOUT0(N__3999),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_5_iopad (
            .OE(N__8806),
            .DIN(N__8805),
            .DOUT(N__8804),
            .PACKAGEPIN(D_UM_040[5]));
    defparam D_UM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_5_preio (
            .PADOEN(N__8806),
            .PADOUT(N__8805),
            .PADIN(N__8804),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7655),
            .DIN0(D_UM_040_in_5),
            .DOUT0(N__7902),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_3_iopad (
            .OE(N__8797),
            .DIN(N__8796),
            .DOUT(N__8795),
            .PACKAGEPIN(D_LL_AMIGA[3]));
    defparam D_LL_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_3_preio (
            .PADOEN(N__8797),
            .PADOUT(N__8796),
            .PADIN(N__8795),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5284),
            .DIN0(D_LL_AMIGA_in_3),
            .DOUT0(N__3965),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_3_iopad (
            .OE(N__8788),
            .DIN(N__8787),
            .DOUT(N__8786),
            .PACKAGEPIN(D_UU_AMIGA[3]));
    defparam D_UU_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_3_preio (
            .PADOEN(N__8788),
            .PADOUT(N__8787),
            .PADIN(N__8786),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5461),
            .DIN0(D_UU_AMIGA_in_3),
            .DOUT0(N__4344),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_5_iopad (
            .OE(N__8779),
            .DIN(N__8778),
            .DOUT(N__8777),
            .PACKAGEPIN(D_LL_040[5]));
    defparam D_LL_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_5_preio (
            .PADOEN(N__8779),
            .PADOUT(N__8778),
            .PADIN(N__8777),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7629),
            .DIN0(D_LL_040_in_5),
            .DOUT0(N__2733),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_6_iopad (
            .OE(N__8770),
            .DIN(N__8769),
            .DOUT(N__8768),
            .PACKAGEPIN(D_LL_AMIGA[6]));
    defparam D_LL_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_6_preio (
            .PADOEN(N__8770),
            .PADOUT(N__8769),
            .PADIN(N__8768),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5397),
            .DIN0(D_LL_AMIGA_in_6),
            .DOUT0(N__3339),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_6_iopad (
            .OE(N__8761),
            .DIN(N__8760),
            .DOUT(N__8759),
            .PACKAGEPIN(D_UU_AMIGA[6]));
    defparam D_UU_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_6_preio (
            .PADOEN(N__8761),
            .PADOUT(N__8760),
            .PADIN(N__8759),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5468),
            .DIN0(D_UU_AMIGA_in_6),
            .DOUT0(N__3132),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_1_iopad (
            .OE(N__8752),
            .DIN(N__8751),
            .DOUT(N__8750),
            .PACKAGEPIN(D_UM_AMIGA[1]));
    defparam D_UM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_1_preio (
            .PADOEN(N__8752),
            .PADOUT(N__8751),
            .PADIN(N__8750),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5371),
            .DIN0(D_UM_AMIGA_in_1),
            .DOUT0(N__6054),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_5_iopad (
            .OE(N__8743),
            .DIN(N__8742),
            .DOUT(N__8741),
            .PACKAGEPIN(D_UU_040[5]));
    defparam D_UU_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_5_preio (
            .PADOEN(N__8743),
            .PADOUT(N__8742),
            .PADIN(N__8741),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7656),
            .DIN0(D_UU_040_in_5),
            .DOUT0(N__4926),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMA_obuf_iopad (
            .OE(N__8734),
            .DIN(N__8733),
            .DOUT(N__8732),
            .PACKAGEPIN(CLKRAMA));
    defparam CLKRAMA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMA_obuf_preio (
            .PADOEN(N__8734),
            .PADOUT(N__8733),
            .PADIN(N__8732),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3564),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_2_iopad (
            .OE(N__8725),
            .DIN(N__8724),
            .DOUT(N__8723),
            .PACKAGEPIN(D_LL_040[2]));
    defparam D_LL_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_2_preio (
            .PADOEN(N__8725),
            .PADOUT(N__8724),
            .PADIN(N__8723),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7631),
            .DIN0(D_LL_040_in_2),
            .DOUT0(N__3768),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCI_CPUn_obuf_iopad (
            .OE(N__8716),
            .DIN(N__8715),
            .DOUT(N__8714),
            .PACKAGEPIN(TCI_CPUn));
    defparam TCI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TCI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TCI_CPUn_obuf_preio (
            .PADOEN(N__8716),
            .PADOUT(N__8715),
            .PADIN(N__8714),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6789),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BBn_ibuf_iopad (
            .OE(N__8707),
            .DIN(N__8706),
            .DOUT(N__8705),
            .PACKAGEPIN(BBn));
    defparam BBn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BBn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BBn_ibuf_preio (
            .PADOEN(N__8707),
            .PADOUT(N__8706),
            .PADIN(N__8705),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(BBn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMAAn_obuf_iopad (
            .OE(N__8698),
            .DIN(N__8697),
            .DOUT(N__8696),
            .PACKAGEPIN(DMAAn));
    defparam DMAAn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMAAn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMAAn_obuf_preio (
            .PADOEN(N__8698),
            .PADOUT(N__8697),
            .PADIN(N__8696),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3642),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_4_iopad (
            .OE(N__8689),
            .DIN(N__8688),
            .DOUT(N__8687),
            .PACKAGEPIN(D_UM_AMIGA[4]));
    defparam D_UM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_4_preio (
            .PADOEN(N__8689),
            .PADOUT(N__8688),
            .PADIN(N__8687),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5433),
            .DIN0(D_UM_AMIGA_in_4),
            .DOUT0(N__2823),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_6_iopad (
            .OE(N__8680),
            .DIN(N__8679),
            .DOUT(N__8678),
            .PACKAGEPIN(D_LM_AMIGA[6]));
    defparam D_LM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_6_preio (
            .PADOEN(N__8680),
            .PADOUT(N__8679),
            .PADIN(N__8678),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5373),
            .DIN0(D_LM_AMIGA_in_6),
            .DOUT0(N__3171),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__8671),
            .DIN(N__8670),
            .DOUT(N__8669),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__8671),
            .PADOUT(N__8670),
            .PADIN(N__8669),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_5_iopad (
            .OE(N__8662),
            .DIN(N__8661),
            .DOUT(N__8660),
            .PACKAGEPIN(D_LM_040[5]));
    defparam D_LM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_5_preio (
            .PADOEN(N__8662),
            .PADOUT(N__8661),
            .PADIN(N__8660),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7560),
            .DIN0(D_LM_040_in_5),
            .DOUT0(N__3438),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_6_iopad (
            .OE(N__8653),
            .DIN(N__8652),
            .DOUT(N__8651),
            .PACKAGEPIN(D_UM_040[6]));
    defparam D_UM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_6_preio (
            .PADOEN(N__8653),
            .PADOUT(N__8652),
            .PADIN(N__8651),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7546),
            .DIN0(D_UM_040_in_6),
            .DOUT0(N__8634),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IoInMux I__2218 (
            .O(N__8634),
            .I(N__8631));
    LocalMux I__2217 (
            .O(N__8631),
            .I(N__8628));
    Span4Mux_s2_h I__2216 (
            .O(N__8628),
            .I(N__8625));
    Sp12to4 I__2215 (
            .O(N__8625),
            .I(N__8622));
    Span12Mux_v I__2214 (
            .O(N__8622),
            .I(N__8619));
    Odrv12 I__2213 (
            .O(N__8619),
            .I(un1_D_UM_AMIGA_6));
    InMux I__2212 (
            .O(N__8616),
            .I(N__8612));
    InMux I__2211 (
            .O(N__8615),
            .I(N__8609));
    LocalMux I__2210 (
            .O(N__8612),
            .I(N__8605));
    LocalMux I__2209 (
            .O(N__8609),
            .I(N__8602));
    InMux I__2208 (
            .O(N__8608),
            .I(N__8599));
    Span4Mux_v I__2207 (
            .O(N__8605),
            .I(N__8596));
    Span4Mux_v I__2206 (
            .O(N__8602),
            .I(N__8591));
    LocalMux I__2205 (
            .O(N__8599),
            .I(N__8591));
    Sp12to4 I__2204 (
            .O(N__8596),
            .I(N__8588));
    Span4Mux_v I__2203 (
            .O(N__8591),
            .I(N__8585));
    Span12Mux_h I__2202 (
            .O(N__8588),
            .I(N__8582));
    Span4Mux_v I__2201 (
            .O(N__8585),
            .I(N__8579));
    Span12Mux_v I__2200 (
            .O(N__8582),
            .I(N__8576));
    Sp12to4 I__2199 (
            .O(N__8579),
            .I(N__8573));
    Span12Mux_v I__2198 (
            .O(N__8576),
            .I(N__8568));
    Span12Mux_h I__2197 (
            .O(N__8573),
            .I(N__8568));
    Odrv12 I__2196 (
            .O(N__8568),
            .I(D_UM_AMIGA_in_3));
    InMux I__2195 (
            .O(N__8565),
            .I(N__8562));
    LocalMux I__2194 (
            .O(N__8562),
            .I(N__8559));
    Odrv4 I__2193 (
            .O(N__8559),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ));
    IoInMux I__2192 (
            .O(N__8556),
            .I(N__8553));
    LocalMux I__2191 (
            .O(N__8553),
            .I(N__8550));
    IoSpan4Mux I__2190 (
            .O(N__8550),
            .I(N__8547));
    Span4Mux_s0_h I__2189 (
            .O(N__8547),
            .I(N__8544));
    Sp12to4 I__2188 (
            .O(N__8544),
            .I(N__8541));
    Span12Mux_h I__2187 (
            .O(N__8541),
            .I(N__8538));
    Odrv12 I__2186 (
            .O(N__8538),
            .I(un1_D_UM_AMIGA_3));
    IoInMux I__2185 (
            .O(N__8535),
            .I(N__8532));
    LocalMux I__2184 (
            .O(N__8532),
            .I(N__8528));
    InMux I__2183 (
            .O(N__8531),
            .I(N__8525));
    IoSpan4Mux I__2182 (
            .O(N__8528),
            .I(N__8522));
    LocalMux I__2181 (
            .O(N__8525),
            .I(N__8519));
    Span4Mux_s3_h I__2180 (
            .O(N__8522),
            .I(N__8516));
    Span4Mux_h I__2179 (
            .O(N__8519),
            .I(N__8513));
    Sp12to4 I__2178 (
            .O(N__8516),
            .I(N__8510));
    Sp12to4 I__2177 (
            .O(N__8513),
            .I(N__8507));
    Span12Mux_v I__2176 (
            .O(N__8510),
            .I(N__8504));
    Span12Mux_v I__2175 (
            .O(N__8507),
            .I(N__8501));
    Span12Mux_h I__2174 (
            .O(N__8504),
            .I(N__8498));
    Span12Mux_v I__2173 (
            .O(N__8501),
            .I(N__8495));
    Span12Mux_h I__2172 (
            .O(N__8498),
            .I(N__8492));
    Span12Mux_h I__2171 (
            .O(N__8495),
            .I(N__8489));
    Odrv12 I__2170 (
            .O(N__8492),
            .I(D_LL_040_in_7));
    Odrv12 I__2169 (
            .O(N__8489),
            .I(D_LL_040_in_7));
    InMux I__2168 (
            .O(N__8484),
            .I(N__8481));
    LocalMux I__2167 (
            .O(N__8481),
            .I(N__8478));
    Span4Mux_v I__2166 (
            .O(N__8478),
            .I(N__8475));
    Span4Mux_v I__2165 (
            .O(N__8475),
            .I(N__8472));
    Sp12to4 I__2164 (
            .O(N__8472),
            .I(N__8469));
    Span12Mux_h I__2163 (
            .O(N__8469),
            .I(N__8466));
    Odrv12 I__2162 (
            .O(N__8466),
            .I(D_UM_040_in_7));
    IoInMux I__2161 (
            .O(N__8463),
            .I(N__8460));
    LocalMux I__2160 (
            .O(N__8460),
            .I(N__8457));
    IoSpan4Mux I__2159 (
            .O(N__8457),
            .I(N__8454));
    Span4Mux_s0_h I__2158 (
            .O(N__8454),
            .I(N__8451));
    Sp12to4 I__2157 (
            .O(N__8451),
            .I(N__8448));
    Span12Mux_s11_h I__2156 (
            .O(N__8448),
            .I(N__8445));
    Odrv12 I__2155 (
            .O(N__8445),
            .I(un1_D_UM_040_7));
    InMux I__2154 (
            .O(N__8442),
            .I(N__8439));
    LocalMux I__2153 (
            .O(N__8439),
            .I(N__8436));
    Span12Mux_s9_v I__2152 (
            .O(N__8436),
            .I(N__8433));
    Odrv12 I__2151 (
            .O(N__8433),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ));
    InMux I__2150 (
            .O(N__8430),
            .I(N__8427));
    LocalMux I__2149 (
            .O(N__8427),
            .I(N__8423));
    InMux I__2148 (
            .O(N__8426),
            .I(N__8419));
    Span4Mux_v I__2147 (
            .O(N__8423),
            .I(N__8416));
    InMux I__2146 (
            .O(N__8422),
            .I(N__8413));
    LocalMux I__2145 (
            .O(N__8419),
            .I(N__8410));
    Span4Mux_v I__2144 (
            .O(N__8416),
            .I(N__8405));
    LocalMux I__2143 (
            .O(N__8413),
            .I(N__8405));
    Span4Mux_v I__2142 (
            .O(N__8410),
            .I(N__8402));
    Span4Mux_v I__2141 (
            .O(N__8405),
            .I(N__8399));
    Sp12to4 I__2140 (
            .O(N__8402),
            .I(N__8396));
    Sp12to4 I__2139 (
            .O(N__8399),
            .I(N__8393));
    Span12Mux_v I__2138 (
            .O(N__8396),
            .I(N__8390));
    Span12Mux_h I__2137 (
            .O(N__8393),
            .I(N__8387));
    Odrv12 I__2136 (
            .O(N__8390),
            .I(D_UM_AMIGA_in_7));
    Odrv12 I__2135 (
            .O(N__8387),
            .I(D_UM_AMIGA_in_7));
    IoInMux I__2134 (
            .O(N__8382),
            .I(N__8379));
    LocalMux I__2133 (
            .O(N__8379),
            .I(N__8376));
    IoSpan4Mux I__2132 (
            .O(N__8376),
            .I(N__8373));
    IoSpan4Mux I__2131 (
            .O(N__8373),
            .I(N__8370));
    Span4Mux_s3_h I__2130 (
            .O(N__8370),
            .I(N__8367));
    Sp12to4 I__2129 (
            .O(N__8367),
            .I(N__8364));
    Odrv12 I__2128 (
            .O(N__8364),
            .I(un1_D_UM_AMIGA_7));
    IoInMux I__2127 (
            .O(N__8361),
            .I(N__8358));
    LocalMux I__2126 (
            .O(N__8358),
            .I(N__8355));
    IoSpan4Mux I__2125 (
            .O(N__8355),
            .I(N__8352));
    IoSpan4Mux I__2124 (
            .O(N__8352),
            .I(N__8349));
    Span4Mux_s2_h I__2123 (
            .O(N__8349),
            .I(N__8345));
    InMux I__2122 (
            .O(N__8348),
            .I(N__8342));
    Sp12to4 I__2121 (
            .O(N__8345),
            .I(N__8339));
    LocalMux I__2120 (
            .O(N__8342),
            .I(N__8336));
    Span12Mux_h I__2119 (
            .O(N__8339),
            .I(N__8333));
    Span12Mux_v I__2118 (
            .O(N__8336),
            .I(N__8330));
    Span12Mux_h I__2117 (
            .O(N__8333),
            .I(N__8327));
    Span12Mux_h I__2116 (
            .O(N__8330),
            .I(N__8324));
    Odrv12 I__2115 (
            .O(N__8327),
            .I(D_LM_040_in_5));
    Odrv12 I__2114 (
            .O(N__8324),
            .I(D_LM_040_in_5));
    InMux I__2113 (
            .O(N__8319),
            .I(N__8316));
    LocalMux I__2112 (
            .O(N__8316),
            .I(N__8313));
    Span12Mux_v I__2111 (
            .O(N__8313),
            .I(N__8310));
    Span12Mux_h I__2110 (
            .O(N__8310),
            .I(N__8307));
    Odrv12 I__2109 (
            .O(N__8307),
            .I(D_UU_040_in_5));
    IoInMux I__2108 (
            .O(N__8304),
            .I(N__8301));
    LocalMux I__2107 (
            .O(N__8301),
            .I(N__8298));
    Span4Mux_s2_h I__2106 (
            .O(N__8298),
            .I(N__8295));
    Span4Mux_v I__2105 (
            .O(N__8295),
            .I(N__8292));
    Sp12to4 I__2104 (
            .O(N__8292),
            .I(N__8289));
    Span12Mux_s10_h I__2103 (
            .O(N__8289),
            .I(N__8286));
    Odrv12 I__2102 (
            .O(N__8286),
            .I(un1_D_UU_040_5));
    InMux I__2101 (
            .O(N__8283),
            .I(N__8280));
    LocalMux I__2100 (
            .O(N__8280),
            .I(N__8277));
    Span12Mux_s7_v I__2099 (
            .O(N__8277),
            .I(N__8274));
    Span12Mux_h I__2098 (
            .O(N__8274),
            .I(N__8271));
    Odrv12 I__2097 (
            .O(N__8271),
            .I(D_UM_040_in_5));
    IoInMux I__2096 (
            .O(N__8268),
            .I(N__8265));
    LocalMux I__2095 (
            .O(N__8265),
            .I(N__8261));
    InMux I__2094 (
            .O(N__8264),
            .I(N__8258));
    IoSpan4Mux I__2093 (
            .O(N__8261),
            .I(N__8255));
    LocalMux I__2092 (
            .O(N__8258),
            .I(N__8252));
    Span4Mux_s3_h I__2091 (
            .O(N__8255),
            .I(N__8249));
    Span4Mux_h I__2090 (
            .O(N__8252),
            .I(N__8246));
    Sp12to4 I__2089 (
            .O(N__8249),
            .I(N__8243));
    Sp12to4 I__2088 (
            .O(N__8246),
            .I(N__8240));
    Span12Mux_v I__2087 (
            .O(N__8243),
            .I(N__8237));
    Span12Mux_v I__2086 (
            .O(N__8240),
            .I(N__8234));
    Span12Mux_h I__2085 (
            .O(N__8237),
            .I(N__8231));
    Span12Mux_v I__2084 (
            .O(N__8234),
            .I(N__8228));
    Span12Mux_h I__2083 (
            .O(N__8231),
            .I(N__8225));
    Span12Mux_h I__2082 (
            .O(N__8228),
            .I(N__8222));
    Odrv12 I__2081 (
            .O(N__8225),
            .I(D_LL_040_in_5));
    Odrv12 I__2080 (
            .O(N__8222),
            .I(D_LL_040_in_5));
    InMux I__2079 (
            .O(N__8217),
            .I(N__8201));
    InMux I__2078 (
            .O(N__8216),
            .I(N__8201));
    InMux I__2077 (
            .O(N__8215),
            .I(N__8198));
    InMux I__2076 (
            .O(N__8214),
            .I(N__8192));
    InMux I__2075 (
            .O(N__8213),
            .I(N__8192));
    InMux I__2074 (
            .O(N__8212),
            .I(N__8187));
    InMux I__2073 (
            .O(N__8211),
            .I(N__8187));
    InMux I__2072 (
            .O(N__8210),
            .I(N__8183));
    InMux I__2071 (
            .O(N__8209),
            .I(N__8178));
    InMux I__2070 (
            .O(N__8208),
            .I(N__8178));
    InMux I__2069 (
            .O(N__8207),
            .I(N__8175));
    InMux I__2068 (
            .O(N__8206),
            .I(N__8169));
    LocalMux I__2067 (
            .O(N__8201),
            .I(N__8162));
    LocalMux I__2066 (
            .O(N__8198),
            .I(N__8162));
    InMux I__2065 (
            .O(N__8197),
            .I(N__8159));
    LocalMux I__2064 (
            .O(N__8192),
            .I(N__8156));
    LocalMux I__2063 (
            .O(N__8187),
            .I(N__8153));
    InMux I__2062 (
            .O(N__8186),
            .I(N__8150));
    LocalMux I__2061 (
            .O(N__8183),
            .I(N__8143));
    LocalMux I__2060 (
            .O(N__8178),
            .I(N__8143));
    LocalMux I__2059 (
            .O(N__8175),
            .I(N__8140));
    InMux I__2058 (
            .O(N__8174),
            .I(N__8131));
    InMux I__2057 (
            .O(N__8173),
            .I(N__8126));
    InMux I__2056 (
            .O(N__8172),
            .I(N__8123));
    LocalMux I__2055 (
            .O(N__8169),
            .I(N__8120));
    InMux I__2054 (
            .O(N__8168),
            .I(N__8115));
    InMux I__2053 (
            .O(N__8167),
            .I(N__8115));
    Span4Mux_v I__2052 (
            .O(N__8162),
            .I(N__8110));
    LocalMux I__2051 (
            .O(N__8159),
            .I(N__8110));
    Span4Mux_h I__2050 (
            .O(N__8156),
            .I(N__8103));
    Span4Mux_h I__2049 (
            .O(N__8153),
            .I(N__8103));
    LocalMux I__2048 (
            .O(N__8150),
            .I(N__8103));
    InMux I__2047 (
            .O(N__8149),
            .I(N__8098));
    InMux I__2046 (
            .O(N__8148),
            .I(N__8098));
    Span4Mux_v I__2045 (
            .O(N__8143),
            .I(N__8093));
    Span4Mux_v I__2044 (
            .O(N__8140),
            .I(N__8093));
    InMux I__2043 (
            .O(N__8139),
            .I(N__8090));
    InMux I__2042 (
            .O(N__8138),
            .I(N__8085));
    InMux I__2041 (
            .O(N__8137),
            .I(N__8085));
    InMux I__2040 (
            .O(N__8136),
            .I(N__8080));
    InMux I__2039 (
            .O(N__8135),
            .I(N__8080));
    InMux I__2038 (
            .O(N__8134),
            .I(N__8077));
    LocalMux I__2037 (
            .O(N__8131),
            .I(N__8074));
    InMux I__2036 (
            .O(N__8130),
            .I(N__8071));
    InMux I__2035 (
            .O(N__8129),
            .I(N__8068));
    LocalMux I__2034 (
            .O(N__8126),
            .I(N__8062));
    LocalMux I__2033 (
            .O(N__8123),
            .I(N__8062));
    Span4Mux_h I__2032 (
            .O(N__8120),
            .I(N__8057));
    LocalMux I__2031 (
            .O(N__8115),
            .I(N__8057));
    Span4Mux_v I__2030 (
            .O(N__8110),
            .I(N__8054));
    Span4Mux_v I__2029 (
            .O(N__8103),
            .I(N__8049));
    LocalMux I__2028 (
            .O(N__8098),
            .I(N__8049));
    Span4Mux_v I__2027 (
            .O(N__8093),
            .I(N__8044));
    LocalMux I__2026 (
            .O(N__8090),
            .I(N__8044));
    LocalMux I__2025 (
            .O(N__8085),
            .I(N__8037));
    LocalMux I__2024 (
            .O(N__8080),
            .I(N__8037));
    LocalMux I__2023 (
            .O(N__8077),
            .I(N__8037));
    Span4Mux_v I__2022 (
            .O(N__8074),
            .I(N__8030));
    LocalMux I__2021 (
            .O(N__8071),
            .I(N__8030));
    LocalMux I__2020 (
            .O(N__8068),
            .I(N__8030));
    InMux I__2019 (
            .O(N__8067),
            .I(N__8027));
    Span12Mux_v I__2018 (
            .O(N__8062),
            .I(N__8021));
    Span4Mux_v I__2017 (
            .O(N__8057),
            .I(N__8018));
    Span4Mux_h I__2016 (
            .O(N__8054),
            .I(N__8013));
    Span4Mux_v I__2015 (
            .O(N__8049),
            .I(N__8013));
    Span4Mux_v I__2014 (
            .O(N__8044),
            .I(N__8006));
    Span4Mux_v I__2013 (
            .O(N__8037),
            .I(N__8006));
    Span4Mux_v I__2012 (
            .O(N__8030),
            .I(N__8006));
    LocalMux I__2011 (
            .O(N__8027),
            .I(N__8003));
    InMux I__2010 (
            .O(N__8026),
            .I(N__7998));
    InMux I__2009 (
            .O(N__8025),
            .I(N__7998));
    InMux I__2008 (
            .O(N__8024),
            .I(N__7995));
    Odrv12 I__2007 (
            .O(N__8021),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv4 I__2006 (
            .O(N__8018),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv4 I__2005 (
            .O(N__8013),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv4 I__2004 (
            .O(N__8006),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv4 I__2003 (
            .O(N__8003),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    LocalMux I__2002 (
            .O(N__7998),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    LocalMux I__2001 (
            .O(N__7995),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    IoInMux I__2000 (
            .O(N__7980),
            .I(N__7977));
    LocalMux I__1999 (
            .O(N__7977),
            .I(N__7974));
    Span12Mux_s6_v I__1998 (
            .O(N__7974),
            .I(N__7971));
    Span12Mux_h I__1997 (
            .O(N__7971),
            .I(N__7968));
    Odrv12 I__1996 (
            .O(N__7968),
            .I(un1_D_UM_040_5));
    InMux I__1995 (
            .O(N__7965),
            .I(N__7962));
    LocalMux I__1994 (
            .O(N__7962),
            .I(N__7959));
    Sp12to4 I__1993 (
            .O(N__7959),
            .I(N__7956));
    Odrv12 I__1992 (
            .O(N__7956),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ));
    InMux I__1991 (
            .O(N__7953),
            .I(N__7949));
    InMux I__1990 (
            .O(N__7952),
            .I(N__7946));
    LocalMux I__1989 (
            .O(N__7949),
            .I(N__7943));
    LocalMux I__1988 (
            .O(N__7946),
            .I(N__7939));
    Span4Mux_v I__1987 (
            .O(N__7943),
            .I(N__7936));
    InMux I__1986 (
            .O(N__7942),
            .I(N__7933));
    Span4Mux_v I__1985 (
            .O(N__7939),
            .I(N__7930));
    Span4Mux_v I__1984 (
            .O(N__7936),
            .I(N__7925));
    LocalMux I__1983 (
            .O(N__7933),
            .I(N__7925));
    Sp12to4 I__1982 (
            .O(N__7930),
            .I(N__7922));
    Span4Mux_v I__1981 (
            .O(N__7925),
            .I(N__7919));
    Span12Mux_h I__1980 (
            .O(N__7922),
            .I(N__7916));
    Sp12to4 I__1979 (
            .O(N__7919),
            .I(N__7913));
    Span12Mux_v I__1978 (
            .O(N__7916),
            .I(N__7910));
    Span12Mux_h I__1977 (
            .O(N__7913),
            .I(N__7907));
    Odrv12 I__1976 (
            .O(N__7910),
            .I(D_UM_AMIGA_in_5));
    Odrv12 I__1975 (
            .O(N__7907),
            .I(D_UM_AMIGA_in_5));
    IoInMux I__1974 (
            .O(N__7902),
            .I(N__7899));
    LocalMux I__1973 (
            .O(N__7899),
            .I(N__7896));
    Span12Mux_s11_v I__1972 (
            .O(N__7896),
            .I(N__7893));
    Span12Mux_h I__1971 (
            .O(N__7893),
            .I(N__7890));
    Odrv12 I__1970 (
            .O(N__7890),
            .I(un1_D_UM_AMIGA_5));
    InMux I__1969 (
            .O(N__7887),
            .I(N__7884));
    LocalMux I__1968 (
            .O(N__7884),
            .I(N__7877));
    InMux I__1967 (
            .O(N__7883),
            .I(N__7867));
    InMux I__1966 (
            .O(N__7882),
            .I(N__7867));
    InMux I__1965 (
            .O(N__7881),
            .I(N__7867));
    InMux I__1964 (
            .O(N__7880),
            .I(N__7867));
    Span4Mux_v I__1963 (
            .O(N__7877),
            .I(N__7858));
    InMux I__1962 (
            .O(N__7876),
            .I(N__7855));
    LocalMux I__1961 (
            .O(N__7867),
            .I(N__7852));
    InMux I__1960 (
            .O(N__7866),
            .I(N__7845));
    InMux I__1959 (
            .O(N__7865),
            .I(N__7845));
    InMux I__1958 (
            .O(N__7864),
            .I(N__7845));
    InMux I__1957 (
            .O(N__7863),
            .I(N__7842));
    InMux I__1956 (
            .O(N__7862),
            .I(N__7837));
    InMux I__1955 (
            .O(N__7861),
            .I(N__7837));
    Odrv4 I__1954 (
            .O(N__7858),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    LocalMux I__1953 (
            .O(N__7855),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    Odrv4 I__1952 (
            .O(N__7852),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    LocalMux I__1951 (
            .O(N__7845),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    LocalMux I__1950 (
            .O(N__7842),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    LocalMux I__1949 (
            .O(N__7837),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    IoInMux I__1948 (
            .O(N__7824),
            .I(N__7821));
    LocalMux I__1947 (
            .O(N__7821),
            .I(N__7817));
    IoInMux I__1946 (
            .O(N__7820),
            .I(N__7814));
    Span4Mux_s0_h I__1945 (
            .O(N__7817),
            .I(N__7811));
    LocalMux I__1944 (
            .O(N__7814),
            .I(N__7808));
    Span4Mux_h I__1943 (
            .O(N__7811),
            .I(N__7802));
    IoSpan4Mux I__1942 (
            .O(N__7808),
            .I(N__7799));
    InMux I__1941 (
            .O(N__7807),
            .I(N__7792));
    InMux I__1940 (
            .O(N__7806),
            .I(N__7792));
    InMux I__1939 (
            .O(N__7805),
            .I(N__7792));
    Span4Mux_h I__1938 (
            .O(N__7802),
            .I(N__7788));
    Span4Mux_s2_v I__1937 (
            .O(N__7799),
            .I(N__7785));
    LocalMux I__1936 (
            .O(N__7792),
            .I(N__7782));
    InMux I__1935 (
            .O(N__7791),
            .I(N__7779));
    Span4Mux_h I__1934 (
            .O(N__7788),
            .I(N__7776));
    Span4Mux_v I__1933 (
            .O(N__7785),
            .I(N__7770));
    Span4Mux_h I__1932 (
            .O(N__7782),
            .I(N__7770));
    LocalMux I__1931 (
            .O(N__7779),
            .I(N__7766));
    Span4Mux_h I__1930 (
            .O(N__7776),
            .I(N__7763));
    InMux I__1929 (
            .O(N__7775),
            .I(N__7760));
    Span4Mux_v I__1928 (
            .O(N__7770),
            .I(N__7757));
    InMux I__1927 (
            .O(N__7769),
            .I(N__7754));
    Span4Mux_h I__1926 (
            .O(N__7766),
            .I(N__7751));
    Span4Mux_v I__1925 (
            .O(N__7763),
            .I(N__7746));
    LocalMux I__1924 (
            .O(N__7760),
            .I(N__7746));
    Span4Mux_v I__1923 (
            .O(N__7757),
            .I(N__7741));
    LocalMux I__1922 (
            .O(N__7754),
            .I(N__7741));
    Sp12to4 I__1921 (
            .O(N__7751),
            .I(N__7738));
    Span4Mux_v I__1920 (
            .O(N__7746),
            .I(N__7735));
    Span4Mux_h I__1919 (
            .O(N__7741),
            .I(N__7732));
    Odrv12 I__1918 (
            .O(N__7738),
            .I(CPUBGn_c));
    Odrv4 I__1917 (
            .O(N__7735),
            .I(CPUBGn_c));
    Odrv4 I__1916 (
            .O(N__7732),
            .I(CPUBGn_c));
    InMux I__1915 (
            .O(N__7725),
            .I(N__7721));
    CascadeMux I__1914 (
            .O(N__7724),
            .I(N__7716));
    LocalMux I__1913 (
            .O(N__7721),
            .I(N__7713));
    CascadeMux I__1912 (
            .O(N__7720),
            .I(N__7710));
    InMux I__1911 (
            .O(N__7719),
            .I(N__7705));
    InMux I__1910 (
            .O(N__7716),
            .I(N__7705));
    Span4Mux_v I__1909 (
            .O(N__7713),
            .I(N__7701));
    InMux I__1908 (
            .O(N__7710),
            .I(N__7698));
    LocalMux I__1907 (
            .O(N__7705),
            .I(N__7695));
    InMux I__1906 (
            .O(N__7704),
            .I(N__7692));
    Span4Mux_h I__1905 (
            .O(N__7701),
            .I(N__7689));
    LocalMux I__1904 (
            .O(N__7698),
            .I(N__7686));
    Span4Mux_h I__1903 (
            .O(N__7695),
            .I(N__7681));
    LocalMux I__1902 (
            .O(N__7692),
            .I(N__7681));
    Span4Mux_v I__1901 (
            .O(N__7689),
            .I(N__7676));
    Span4Mux_v I__1900 (
            .O(N__7686),
            .I(N__7676));
    Span4Mux_v I__1899 (
            .O(N__7681),
            .I(N__7673));
    Sp12to4 I__1898 (
            .O(N__7676),
            .I(N__7670));
    Sp12to4 I__1897 (
            .O(N__7673),
            .I(N__7667));
    Span12Mux_h I__1896 (
            .O(N__7670),
            .I(N__7664));
    Span12Mux_h I__1895 (
            .O(N__7667),
            .I(N__7661));
    Odrv12 I__1894 (
            .O(N__7664),
            .I(RnW_c));
    Odrv12 I__1893 (
            .O(N__7661),
            .I(RnW_c));
    IoInMux I__1892 (
            .O(N__7656),
            .I(N__7650));
    IoInMux I__1891 (
            .O(N__7655),
            .I(N__7647));
    IoInMux I__1890 (
            .O(N__7654),
            .I(N__7641));
    IoInMux I__1889 (
            .O(N__7653),
            .I(N__7638));
    LocalMux I__1888 (
            .O(N__7650),
            .I(N__7624));
    LocalMux I__1887 (
            .O(N__7647),
            .I(N__7624));
    IoInMux I__1886 (
            .O(N__7646),
            .I(N__7621));
    IoInMux I__1885 (
            .O(N__7645),
            .I(N__7618));
    IoInMux I__1884 (
            .O(N__7644),
            .I(N__7615));
    LocalMux I__1883 (
            .O(N__7641),
            .I(N__7611));
    LocalMux I__1882 (
            .O(N__7638),
            .I(N__7607));
    IoInMux I__1881 (
            .O(N__7637),
            .I(N__7604));
    IoInMux I__1880 (
            .O(N__7636),
            .I(N__7601));
    IoInMux I__1879 (
            .O(N__7635),
            .I(N__7597));
    IoInMux I__1878 (
            .O(N__7634),
            .I(N__7594));
    IoInMux I__1877 (
            .O(N__7633),
            .I(N__7591));
    IoInMux I__1876 (
            .O(N__7632),
            .I(N__7588));
    IoInMux I__1875 (
            .O(N__7631),
            .I(N__7585));
    IoInMux I__1874 (
            .O(N__7630),
            .I(N__7582));
    IoInMux I__1873 (
            .O(N__7629),
            .I(N__7579));
    IoSpan4Mux I__1872 (
            .O(N__7624),
            .I(N__7570));
    LocalMux I__1871 (
            .O(N__7621),
            .I(N__7570));
    LocalMux I__1870 (
            .O(N__7618),
            .I(N__7570));
    LocalMux I__1869 (
            .O(N__7615),
            .I(N__7570));
    IoInMux I__1868 (
            .O(N__7614),
            .I(N__7567));
    Span4Mux_s2_h I__1867 (
            .O(N__7611),
            .I(N__7564));
    IoInMux I__1866 (
            .O(N__7610),
            .I(N__7561));
    IoSpan4Mux I__1865 (
            .O(N__7607),
            .I(N__7551));
    LocalMux I__1864 (
            .O(N__7604),
            .I(N__7551));
    LocalMux I__1863 (
            .O(N__7601),
            .I(N__7551));
    IoInMux I__1862 (
            .O(N__7600),
            .I(N__7548));
    LocalMux I__1861 (
            .O(N__7597),
            .I(N__7541));
    LocalMux I__1860 (
            .O(N__7594),
            .I(N__7541));
    LocalMux I__1859 (
            .O(N__7591),
            .I(N__7530));
    LocalMux I__1858 (
            .O(N__7588),
            .I(N__7530));
    LocalMux I__1857 (
            .O(N__7585),
            .I(N__7530));
    LocalMux I__1856 (
            .O(N__7582),
            .I(N__7530));
    LocalMux I__1855 (
            .O(N__7579),
            .I(N__7530));
    IoSpan4Mux I__1854 (
            .O(N__7570),
            .I(N__7524));
    LocalMux I__1853 (
            .O(N__7567),
            .I(N__7521));
    Span4Mux_v I__1852 (
            .O(N__7564),
            .I(N__7516));
    LocalMux I__1851 (
            .O(N__7561),
            .I(N__7516));
    IoInMux I__1850 (
            .O(N__7560),
            .I(N__7513));
    IoInMux I__1849 (
            .O(N__7559),
            .I(N__7510));
    IoInMux I__1848 (
            .O(N__7558),
            .I(N__7507));
    IoSpan4Mux I__1847 (
            .O(N__7551),
            .I(N__7502));
    LocalMux I__1846 (
            .O(N__7548),
            .I(N__7502));
    IoInMux I__1845 (
            .O(N__7547),
            .I(N__7499));
    IoInMux I__1844 (
            .O(N__7546),
            .I(N__7496));
    Span4Mux_s3_h I__1843 (
            .O(N__7541),
            .I(N__7491));
    IoSpan4Mux I__1842 (
            .O(N__7530),
            .I(N__7488));
    IoInMux I__1841 (
            .O(N__7529),
            .I(N__7485));
    IoInMux I__1840 (
            .O(N__7528),
            .I(N__7482));
    IoInMux I__1839 (
            .O(N__7527),
            .I(N__7476));
    Span4Mux_s2_v I__1838 (
            .O(N__7524),
            .I(N__7473));
    Span4Mux_s2_v I__1837 (
            .O(N__7521),
            .I(N__7470));
    IoSpan4Mux I__1836 (
            .O(N__7516),
            .I(N__7461));
    LocalMux I__1835 (
            .O(N__7513),
            .I(N__7461));
    LocalMux I__1834 (
            .O(N__7510),
            .I(N__7461));
    LocalMux I__1833 (
            .O(N__7507),
            .I(N__7461));
    IoSpan4Mux I__1832 (
            .O(N__7502),
            .I(N__7454));
    LocalMux I__1831 (
            .O(N__7499),
            .I(N__7454));
    LocalMux I__1830 (
            .O(N__7496),
            .I(N__7454));
    IoInMux I__1829 (
            .O(N__7495),
            .I(N__7451));
    IoInMux I__1828 (
            .O(N__7494),
            .I(N__7448));
    Span4Mux_v I__1827 (
            .O(N__7491),
            .I(N__7443));
    Span4Mux_s3_h I__1826 (
            .O(N__7488),
            .I(N__7443));
    LocalMux I__1825 (
            .O(N__7485),
            .I(N__7440));
    LocalMux I__1824 (
            .O(N__7482),
            .I(N__7437));
    IoInMux I__1823 (
            .O(N__7481),
            .I(N__7434));
    IoInMux I__1822 (
            .O(N__7480),
            .I(N__7431));
    IoInMux I__1821 (
            .O(N__7479),
            .I(N__7428));
    LocalMux I__1820 (
            .O(N__7476),
            .I(N__7425));
    Span4Mux_v I__1819 (
            .O(N__7473),
            .I(N__7420));
    Span4Mux_v I__1818 (
            .O(N__7470),
            .I(N__7420));
    IoSpan4Mux I__1817 (
            .O(N__7461),
            .I(N__7415));
    IoSpan4Mux I__1816 (
            .O(N__7454),
            .I(N__7415));
    LocalMux I__1815 (
            .O(N__7451),
            .I(N__7410));
    LocalMux I__1814 (
            .O(N__7448),
            .I(N__7410));
    Sp12to4 I__1813 (
            .O(N__7443),
            .I(N__7403));
    Sp12to4 I__1812 (
            .O(N__7440),
            .I(N__7403));
    Span12Mux_s1_h I__1811 (
            .O(N__7437),
            .I(N__7403));
    LocalMux I__1810 (
            .O(N__7434),
            .I(N__7398));
    LocalMux I__1809 (
            .O(N__7431),
            .I(N__7398));
    LocalMux I__1808 (
            .O(N__7428),
            .I(N__7395));
    Span4Mux_s3_v I__1807 (
            .O(N__7425),
            .I(N__7392));
    Span4Mux_v I__1806 (
            .O(N__7420),
            .I(N__7389));
    Span4Mux_s2_h I__1805 (
            .O(N__7415),
            .I(N__7386));
    Span12Mux_s8_h I__1804 (
            .O(N__7410),
            .I(N__7383));
    Span12Mux_h I__1803 (
            .O(N__7403),
            .I(N__7380));
    Span12Mux_s3_v I__1802 (
            .O(N__7398),
            .I(N__7373));
    Sp12to4 I__1801 (
            .O(N__7395),
            .I(N__7373));
    Sp12to4 I__1800 (
            .O(N__7392),
            .I(N__7373));
    Span4Mux_v I__1799 (
            .O(N__7389),
            .I(N__7368));
    Span4Mux_h I__1798 (
            .O(N__7386),
            .I(N__7368));
    Span12Mux_v I__1797 (
            .O(N__7383),
            .I(N__7365));
    Span12Mux_v I__1796 (
            .O(N__7380),
            .I(N__7360));
    Span12Mux_h I__1795 (
            .O(N__7373),
            .I(N__7360));
    Span4Mux_h I__1794 (
            .O(N__7368),
            .I(N__7357));
    Odrv12 I__1793 (
            .O(N__7365),
            .I(N_60_i));
    Odrv12 I__1792 (
            .O(N__7360),
            .I(N_60_i));
    Odrv4 I__1791 (
            .O(N__7357),
            .I(N_60_i));
    InMux I__1790 (
            .O(N__7350),
            .I(N__7345));
    InMux I__1789 (
            .O(N__7349),
            .I(N__7334));
    InMux I__1788 (
            .O(N__7348),
            .I(N__7334));
    LocalMux I__1787 (
            .O(N__7345),
            .I(N__7330));
    InMux I__1786 (
            .O(N__7344),
            .I(N__7327));
    InMux I__1785 (
            .O(N__7343),
            .I(N__7324));
    InMux I__1784 (
            .O(N__7342),
            .I(N__7310));
    InMux I__1783 (
            .O(N__7341),
            .I(N__7310));
    InMux I__1782 (
            .O(N__7340),
            .I(N__7310));
    InMux I__1781 (
            .O(N__7339),
            .I(N__7310));
    LocalMux I__1780 (
            .O(N__7334),
            .I(N__7306));
    InMux I__1779 (
            .O(N__7333),
            .I(N__7303));
    Span4Mux_v I__1778 (
            .O(N__7330),
            .I(N__7298));
    LocalMux I__1777 (
            .O(N__7327),
            .I(N__7298));
    LocalMux I__1776 (
            .O(N__7324),
            .I(N__7295));
    InMux I__1775 (
            .O(N__7323),
            .I(N__7292));
    InMux I__1774 (
            .O(N__7322),
            .I(N__7289));
    InMux I__1773 (
            .O(N__7321),
            .I(N__7286));
    InMux I__1772 (
            .O(N__7320),
            .I(N__7281));
    InMux I__1771 (
            .O(N__7319),
            .I(N__7281));
    LocalMux I__1770 (
            .O(N__7310),
            .I(N__7277));
    InMux I__1769 (
            .O(N__7309),
            .I(N__7274));
    Span4Mux_v I__1768 (
            .O(N__7306),
            .I(N__7269));
    LocalMux I__1767 (
            .O(N__7303),
            .I(N__7269));
    Span4Mux_v I__1766 (
            .O(N__7298),
            .I(N__7258));
    Span4Mux_h I__1765 (
            .O(N__7295),
            .I(N__7258));
    LocalMux I__1764 (
            .O(N__7292),
            .I(N__7258));
    LocalMux I__1763 (
            .O(N__7289),
            .I(N__7258));
    LocalMux I__1762 (
            .O(N__7286),
            .I(N__7258));
    LocalMux I__1761 (
            .O(N__7281),
            .I(N__7255));
    CascadeMux I__1760 (
            .O(N__7280),
            .I(N__7252));
    Sp12to4 I__1759 (
            .O(N__7277),
            .I(N__7247));
    LocalMux I__1758 (
            .O(N__7274),
            .I(N__7247));
    Span4Mux_v I__1757 (
            .O(N__7269),
            .I(N__7244));
    Span4Mux_v I__1756 (
            .O(N__7258),
            .I(N__7239));
    Span4Mux_v I__1755 (
            .O(N__7255),
            .I(N__7239));
    InMux I__1754 (
            .O(N__7252),
            .I(N__7236));
    Odrv12 I__1753 (
            .O(N__7247),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    Odrv4 I__1752 (
            .O(N__7244),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    Odrv4 I__1751 (
            .O(N__7239),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    LocalMux I__1750 (
            .O(N__7236),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    InMux I__1749 (
            .O(N__7227),
            .I(N__7224));
    LocalMux I__1748 (
            .O(N__7224),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ));
    InMux I__1747 (
            .O(N__7221),
            .I(N__7218));
    LocalMux I__1746 (
            .O(N__7218),
            .I(N__7215));
    Span4Mux_v I__1745 (
            .O(N__7215),
            .I(N__7212));
    Span4Mux_v I__1744 (
            .O(N__7212),
            .I(N__7207));
    InMux I__1743 (
            .O(N__7211),
            .I(N__7204));
    InMux I__1742 (
            .O(N__7210),
            .I(N__7201));
    Sp12to4 I__1741 (
            .O(N__7207),
            .I(N__7194));
    LocalMux I__1740 (
            .O(N__7204),
            .I(N__7194));
    LocalMux I__1739 (
            .O(N__7201),
            .I(N__7194));
    Span12Mux_h I__1738 (
            .O(N__7194),
            .I(N__7191));
    Span12Mux_v I__1737 (
            .O(N__7191),
            .I(N__7188));
    Odrv12 I__1736 (
            .O(N__7188),
            .I(D_UM_AMIGA_in_6));
    InMux I__1735 (
            .O(N__7185),
            .I(N__7182));
    LocalMux I__1734 (
            .O(N__7182),
            .I(N__7179));
    Span4Mux_v I__1733 (
            .O(N__7179),
            .I(N__7174));
    InMux I__1732 (
            .O(N__7178),
            .I(N__7171));
    InMux I__1731 (
            .O(N__7177),
            .I(N__7168));
    Span4Mux_v I__1730 (
            .O(N__7174),
            .I(N__7161));
    LocalMux I__1729 (
            .O(N__7171),
            .I(N__7161));
    LocalMux I__1728 (
            .O(N__7168),
            .I(N__7161));
    Span4Mux_v I__1727 (
            .O(N__7161),
            .I(N__7158));
    Sp12to4 I__1726 (
            .O(N__7158),
            .I(N__7155));
    Span12Mux_h I__1725 (
            .O(N__7155),
            .I(N__7152));
    Odrv12 I__1724 (
            .O(N__7152),
            .I(D_UM_AMIGA_in_0));
    InMux I__1723 (
            .O(N__7149),
            .I(N__7146));
    LocalMux I__1722 (
            .O(N__7146),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ));
    InMux I__1721 (
            .O(N__7143),
            .I(N__7140));
    LocalMux I__1720 (
            .O(N__7140),
            .I(N__7137));
    Glb2LocalMux I__1719 (
            .O(N__7137),
            .I(N__7089));
    ClkMux I__1718 (
            .O(N__7136),
            .I(N__7089));
    ClkMux I__1717 (
            .O(N__7135),
            .I(N__7089));
    ClkMux I__1716 (
            .O(N__7134),
            .I(N__7089));
    ClkMux I__1715 (
            .O(N__7133),
            .I(N__7089));
    ClkMux I__1714 (
            .O(N__7132),
            .I(N__7089));
    ClkMux I__1713 (
            .O(N__7131),
            .I(N__7089));
    ClkMux I__1712 (
            .O(N__7130),
            .I(N__7089));
    ClkMux I__1711 (
            .O(N__7129),
            .I(N__7089));
    ClkMux I__1710 (
            .O(N__7128),
            .I(N__7089));
    ClkMux I__1709 (
            .O(N__7127),
            .I(N__7089));
    ClkMux I__1708 (
            .O(N__7126),
            .I(N__7089));
    ClkMux I__1707 (
            .O(N__7125),
            .I(N__7089));
    ClkMux I__1706 (
            .O(N__7124),
            .I(N__7089));
    ClkMux I__1705 (
            .O(N__7123),
            .I(N__7089));
    ClkMux I__1704 (
            .O(N__7122),
            .I(N__7089));
    GlobalMux I__1703 (
            .O(N__7089),
            .I(CLK40));
    CEMux I__1702 (
            .O(N__7086),
            .I(N__7082));
    CEMux I__1701 (
            .O(N__7085),
            .I(N__7079));
    LocalMux I__1700 (
            .O(N__7082),
            .I(N__7076));
    LocalMux I__1699 (
            .O(N__7079),
            .I(N__7072));
    Span4Mux_v I__1698 (
            .O(N__7076),
            .I(N__7069));
    CEMux I__1697 (
            .O(N__7075),
            .I(N__7066));
    Span4Mux_v I__1696 (
            .O(N__7072),
            .I(N__7063));
    Span4Mux_h I__1695 (
            .O(N__7069),
            .I(N__7060));
    LocalMux I__1694 (
            .O(N__7066),
            .I(N__7057));
    Span4Mux_h I__1693 (
            .O(N__7063),
            .I(N__7054));
    Odrv4 I__1692 (
            .O(N__7060),
            .I(\U111_CYCLE_SM.N_99_i_0 ));
    Odrv12 I__1691 (
            .O(N__7057),
            .I(\U111_CYCLE_SM.N_99_i_0 ));
    Odrv4 I__1690 (
            .O(N__7054),
            .I(\U111_CYCLE_SM.N_99_i_0 ));
    SRMux I__1689 (
            .O(N__7047),
            .I(N__7043));
    SRMux I__1688 (
            .O(N__7046),
            .I(N__7040));
    LocalMux I__1687 (
            .O(N__7043),
            .I(N__7036));
    LocalMux I__1686 (
            .O(N__7040),
            .I(N__7033));
    SRMux I__1685 (
            .O(N__7039),
            .I(N__7030));
    Span4Mux_h I__1684 (
            .O(N__7036),
            .I(N__7027));
    Span4Mux_h I__1683 (
            .O(N__7033),
            .I(N__7024));
    LocalMux I__1682 (
            .O(N__7030),
            .I(N__7021));
    Odrv4 I__1681 (
            .O(N__7027),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81 ));
    Odrv4 I__1680 (
            .O(N__7024),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81 ));
    Odrv12 I__1679 (
            .O(N__7021),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81 ));
    InMux I__1678 (
            .O(N__7014),
            .I(N__7011));
    LocalMux I__1677 (
            .O(N__7011),
            .I(N__7008));
    Span4Mux_v I__1676 (
            .O(N__7008),
            .I(N__7003));
    InMux I__1675 (
            .O(N__7007),
            .I(N__7000));
    InMux I__1674 (
            .O(N__7006),
            .I(N__6997));
    Sp12to4 I__1673 (
            .O(N__7003),
            .I(N__6994));
    LocalMux I__1672 (
            .O(N__7000),
            .I(N__6989));
    LocalMux I__1671 (
            .O(N__6997),
            .I(N__6989));
    Span12Mux_h I__1670 (
            .O(N__6994),
            .I(N__6986));
    Span12Mux_v I__1669 (
            .O(N__6989),
            .I(N__6983));
    Span12Mux_v I__1668 (
            .O(N__6986),
            .I(N__6980));
    Span12Mux_h I__1667 (
            .O(N__6983),
            .I(N__6977));
    Odrv12 I__1666 (
            .O(N__6980),
            .I(D_UM_AMIGA_in_1));
    Odrv12 I__1665 (
            .O(N__6977),
            .I(D_UM_AMIGA_in_1));
    InMux I__1664 (
            .O(N__6972),
            .I(N__6969));
    LocalMux I__1663 (
            .O(N__6969),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ));
    IoInMux I__1662 (
            .O(N__6966),
            .I(N__6963));
    LocalMux I__1661 (
            .O(N__6963),
            .I(N__6960));
    Span4Mux_s2_h I__1660 (
            .O(N__6960),
            .I(N__6957));
    Sp12to4 I__1659 (
            .O(N__6957),
            .I(N__6954));
    Span12Mux_s11_v I__1658 (
            .O(N__6954),
            .I(N__6951));
    Span12Mux_h I__1657 (
            .O(N__6951),
            .I(N__6948));
    Odrv12 I__1656 (
            .O(N__6948),
            .I(un1_D_UM_AMIGA_1));
    InMux I__1655 (
            .O(N__6945),
            .I(N__6942));
    LocalMux I__1654 (
            .O(N__6942),
            .I(N__6937));
    InMux I__1653 (
            .O(N__6941),
            .I(N__6934));
    CascadeMux I__1652 (
            .O(N__6940),
            .I(N__6931));
    Span4Mux_v I__1651 (
            .O(N__6937),
            .I(N__6926));
    LocalMux I__1650 (
            .O(N__6934),
            .I(N__6926));
    InMux I__1649 (
            .O(N__6931),
            .I(N__6923));
    Odrv4 I__1648 (
            .O(N__6926),
            .I(\U111_CYCLE_SM.TA_DISZ0 ));
    LocalMux I__1647 (
            .O(N__6923),
            .I(\U111_CYCLE_SM.TA_DISZ0 ));
    IoInMux I__1646 (
            .O(N__6918),
            .I(N__6915));
    LocalMux I__1645 (
            .O(N__6915),
            .I(N__6912));
    Span4Mux_s1_v I__1644 (
            .O(N__6912),
            .I(N__6909));
    Span4Mux_v I__1643 (
            .O(N__6909),
            .I(N__6906));
    Span4Mux_v I__1642 (
            .O(N__6906),
            .I(N__6903));
    Span4Mux_v I__1641 (
            .O(N__6903),
            .I(N__6900));
    Odrv4 I__1640 (
            .O(N__6900),
            .I(N_64));
    InMux I__1639 (
            .O(N__6897),
            .I(N__6894));
    LocalMux I__1638 (
            .O(N__6894),
            .I(N__6891));
    Span4Mux_v I__1637 (
            .O(N__6891),
            .I(N__6888));
    Sp12to4 I__1636 (
            .O(N__6888),
            .I(N__6885));
    Span12Mux_h I__1635 (
            .O(N__6885),
            .I(N__6882));
    Span12Mux_v I__1634 (
            .O(N__6882),
            .I(N__6879));
    Odrv12 I__1633 (
            .O(N__6879),
            .I(TCIn_c));
    CascadeMux I__1632 (
            .O(N__6876),
            .I(N__6872));
    InMux I__1631 (
            .O(N__6875),
            .I(N__6869));
    InMux I__1630 (
            .O(N__6872),
            .I(N__6866));
    LocalMux I__1629 (
            .O(N__6869),
            .I(N__6863));
    LocalMux I__1628 (
            .O(N__6866),
            .I(N__6858));
    Span4Mux_v I__1627 (
            .O(N__6863),
            .I(N__6855));
    InMux I__1626 (
            .O(N__6862),
            .I(N__6850));
    InMux I__1625 (
            .O(N__6861),
            .I(N__6850));
    Span4Mux_v I__1624 (
            .O(N__6858),
            .I(N__6846));
    Span4Mux_v I__1623 (
            .O(N__6855),
            .I(N__6843));
    LocalMux I__1622 (
            .O(N__6850),
            .I(N__6840));
    InMux I__1621 (
            .O(N__6849),
            .I(N__6836));
    Span4Mux_v I__1620 (
            .O(N__6846),
            .I(N__6832));
    Sp12to4 I__1619 (
            .O(N__6843),
            .I(N__6829));
    Span4Mux_h I__1618 (
            .O(N__6840),
            .I(N__6826));
    InMux I__1617 (
            .O(N__6839),
            .I(N__6823));
    LocalMux I__1616 (
            .O(N__6836),
            .I(N__6820));
    InMux I__1615 (
            .O(N__6835),
            .I(N__6817));
    Sp12to4 I__1614 (
            .O(N__6832),
            .I(N__6814));
    Span12Mux_h I__1613 (
            .O(N__6829),
            .I(N__6807));
    Sp12to4 I__1612 (
            .O(N__6826),
            .I(N__6807));
    LocalMux I__1611 (
            .O(N__6823),
            .I(N__6807));
    Span4Mux_h I__1610 (
            .O(N__6820),
            .I(N__6802));
    LocalMux I__1609 (
            .O(N__6817),
            .I(N__6802));
    Span12Mux_h I__1608 (
            .O(N__6814),
            .I(N__6797));
    Span12Mux_v I__1607 (
            .O(N__6807),
            .I(N__6797));
    Span4Mux_v I__1606 (
            .O(N__6802),
            .I(N__6794));
    Odrv12 I__1605 (
            .O(N__6797),
            .I(LBENn_c));
    Odrv4 I__1604 (
            .O(N__6794),
            .I(LBENn_c));
    IoInMux I__1603 (
            .O(N__6789),
            .I(N__6786));
    LocalMux I__1602 (
            .O(N__6786),
            .I(N__6783));
    Span4Mux_s3_h I__1601 (
            .O(N__6783),
            .I(N__6780));
    Span4Mux_v I__1600 (
            .O(N__6780),
            .I(N__6777));
    Span4Mux_v I__1599 (
            .O(N__6777),
            .I(N__6774));
    Sp12to4 I__1598 (
            .O(N__6774),
            .I(N__6771));
    Odrv12 I__1597 (
            .O(N__6771),
            .I(U111_CYCLE_SM_TCI_CPUn_0_i));
    IoInMux I__1596 (
            .O(N__6768),
            .I(N__6765));
    LocalMux I__1595 (
            .O(N__6765),
            .I(N__6762));
    Span4Mux_s2_v I__1594 (
            .O(N__6762),
            .I(N__6759));
    Span4Mux_h I__1593 (
            .O(N__6759),
            .I(N__6756));
    Span4Mux_h I__1592 (
            .O(N__6756),
            .I(N__6753));
    Span4Mux_v I__1591 (
            .O(N__6753),
            .I(N__6750));
    Odrv4 I__1590 (
            .O(N__6750),
            .I(un1_D_UU_AMIGA_0));
    InMux I__1589 (
            .O(N__6747),
            .I(N__6744));
    LocalMux I__1588 (
            .O(N__6744),
            .I(N__6740));
    InMux I__1587 (
            .O(N__6743),
            .I(N__6737));
    Odrv12 I__1586 (
            .O(N__6740),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ));
    LocalMux I__1585 (
            .O(N__6737),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ));
    CascadeMux I__1584 (
            .O(N__6732),
            .I(N__6729));
    InMux I__1583 (
            .O(N__6729),
            .I(N__6725));
    InMux I__1582 (
            .O(N__6728),
            .I(N__6722));
    LocalMux I__1581 (
            .O(N__6725),
            .I(N__6719));
    LocalMux I__1580 (
            .O(N__6722),
            .I(N__6715));
    Span4Mux_v I__1579 (
            .O(N__6719),
            .I(N__6712));
    InMux I__1578 (
            .O(N__6718),
            .I(N__6709));
    Span4Mux_v I__1577 (
            .O(N__6715),
            .I(N__6706));
    Span4Mux_v I__1576 (
            .O(N__6712),
            .I(N__6701));
    LocalMux I__1575 (
            .O(N__6709),
            .I(N__6701));
    Span4Mux_v I__1574 (
            .O(N__6706),
            .I(N__6698));
    Span4Mux_v I__1573 (
            .O(N__6701),
            .I(N__6695));
    Span4Mux_v I__1572 (
            .O(N__6698),
            .I(N__6692));
    Span4Mux_h I__1571 (
            .O(N__6695),
            .I(N__6689));
    Sp12to4 I__1570 (
            .O(N__6692),
            .I(N__6684));
    Sp12to4 I__1569 (
            .O(N__6689),
            .I(N__6684));
    Span12Mux_h I__1568 (
            .O(N__6684),
            .I(N__6681));
    Odrv12 I__1567 (
            .O(N__6681),
            .I(D_UU_AMIGA_in_3));
    IoInMux I__1566 (
            .O(N__6678),
            .I(N__6675));
    LocalMux I__1565 (
            .O(N__6675),
            .I(N__6672));
    IoSpan4Mux I__1564 (
            .O(N__6672),
            .I(N__6669));
    IoSpan4Mux I__1563 (
            .O(N__6669),
            .I(N__6666));
    IoSpan4Mux I__1562 (
            .O(N__6666),
            .I(N__6663));
    Span4Mux_s2_v I__1561 (
            .O(N__6663),
            .I(N__6660));
    Span4Mux_v I__1560 (
            .O(N__6660),
            .I(N__6657));
    Odrv4 I__1559 (
            .O(N__6657),
            .I(N_117));
    InMux I__1558 (
            .O(N__6654),
            .I(N__6651));
    LocalMux I__1557 (
            .O(N__6651),
            .I(N__6648));
    Span12Mux_v I__1556 (
            .O(N__6648),
            .I(N__6645));
    Span12Mux_h I__1555 (
            .O(N__6645),
            .I(N__6642));
    Odrv12 I__1554 (
            .O(N__6642),
            .I(D_LL_AMIGA_in_0));
    IoInMux I__1553 (
            .O(N__6639),
            .I(N__6636));
    LocalMux I__1552 (
            .O(N__6636),
            .I(N__6633));
    Span4Mux_s2_h I__1551 (
            .O(N__6633),
            .I(N__6630));
    Span4Mux_h I__1550 (
            .O(N__6630),
            .I(N__6627));
    Sp12to4 I__1549 (
            .O(N__6627),
            .I(N__6624));
    Span12Mux_s6_v I__1548 (
            .O(N__6624),
            .I(N__6621));
    Odrv12 I__1547 (
            .O(N__6621),
            .I(un2_D_LL_AMIGA_0));
    InMux I__1546 (
            .O(N__6618),
            .I(N__6615));
    LocalMux I__1545 (
            .O(N__6615),
            .I(N__6612));
    Span4Mux_h I__1544 (
            .O(N__6612),
            .I(N__6609));
    Span4Mux_h I__1543 (
            .O(N__6609),
            .I(N__6605));
    InMux I__1542 (
            .O(N__6608),
            .I(N__6602));
    Sp12to4 I__1541 (
            .O(N__6605),
            .I(N__6599));
    LocalMux I__1540 (
            .O(N__6602),
            .I(N__6596));
    Span12Mux_v I__1539 (
            .O(N__6599),
            .I(N__6591));
    Span12Mux_h I__1538 (
            .O(N__6596),
            .I(N__6591));
    Odrv12 I__1537 (
            .O(N__6591),
            .I(TBIn_c));
    IoInMux I__1536 (
            .O(N__6588),
            .I(N__6585));
    LocalMux I__1535 (
            .O(N__6585),
            .I(N__6582));
    Span12Mux_s6_v I__1534 (
            .O(N__6582),
            .I(N__6579));
    Odrv12 I__1533 (
            .O(N__6579),
            .I(U111_CYCLE_SM_TBI_CPUn_0_i));
    InMux I__1532 (
            .O(N__6576),
            .I(N__6573));
    LocalMux I__1531 (
            .O(N__6573),
            .I(N__6570));
    Span4Mux_v I__1530 (
            .O(N__6570),
            .I(N__6567));
    Sp12to4 I__1529 (
            .O(N__6567),
            .I(N__6564));
    Span12Mux_h I__1528 (
            .O(N__6564),
            .I(N__6561));
    Odrv12 I__1527 (
            .O(N__6561),
            .I(D_LL_AMIGA_in_6));
    IoInMux I__1526 (
            .O(N__6558),
            .I(N__6555));
    LocalMux I__1525 (
            .O(N__6555),
            .I(N__6552));
    Span4Mux_s3_h I__1524 (
            .O(N__6552),
            .I(N__6549));
    Span4Mux_v I__1523 (
            .O(N__6549),
            .I(N__6546));
    Span4Mux_v I__1522 (
            .O(N__6546),
            .I(N__6543));
    Sp12to4 I__1521 (
            .O(N__6543),
            .I(N__6540));
    Odrv12 I__1520 (
            .O(N__6540),
            .I(un2_D_LL_AMIGA_6));
    IoInMux I__1519 (
            .O(N__6537),
            .I(N__6534));
    LocalMux I__1518 (
            .O(N__6534),
            .I(N__6531));
    Span12Mux_s3_h I__1517 (
            .O(N__6531),
            .I(N__6528));
    Odrv12 I__1516 (
            .O(N__6528),
            .I(un1_D_UM_AMIGA_2));
    IoInMux I__1515 (
            .O(N__6525),
            .I(N__6522));
    LocalMux I__1514 (
            .O(N__6522),
            .I(N__6519));
    IoSpan4Mux I__1513 (
            .O(N__6519),
            .I(N__6516));
    Span4Mux_s3_h I__1512 (
            .O(N__6516),
            .I(N__6513));
    Span4Mux_h I__1511 (
            .O(N__6513),
            .I(N__6510));
    Span4Mux_h I__1510 (
            .O(N__6510),
            .I(N__6507));
    Odrv4 I__1509 (
            .O(N__6507),
            .I(un1_D_UM_AMIGA_0));
    InMux I__1508 (
            .O(N__6504),
            .I(N__6499));
    InMux I__1507 (
            .O(N__6503),
            .I(N__6495));
    InMux I__1506 (
            .O(N__6502),
            .I(N__6492));
    LocalMux I__1505 (
            .O(N__6499),
            .I(N__6488));
    InMux I__1504 (
            .O(N__6498),
            .I(N__6485));
    LocalMux I__1503 (
            .O(N__6495),
            .I(N__6481));
    LocalMux I__1502 (
            .O(N__6492),
            .I(N__6478));
    InMux I__1501 (
            .O(N__6491),
            .I(N__6475));
    Span4Mux_v I__1500 (
            .O(N__6488),
            .I(N__6472));
    LocalMux I__1499 (
            .O(N__6485),
            .I(N__6469));
    InMux I__1498 (
            .O(N__6484),
            .I(N__6466));
    Span4Mux_v I__1497 (
            .O(N__6481),
            .I(N__6459));
    Span4Mux_h I__1496 (
            .O(N__6478),
            .I(N__6459));
    LocalMux I__1495 (
            .O(N__6475),
            .I(N__6459));
    Span4Mux_h I__1494 (
            .O(N__6472),
            .I(N__6452));
    Span4Mux_v I__1493 (
            .O(N__6469),
            .I(N__6452));
    LocalMux I__1492 (
            .O(N__6466),
            .I(N__6452));
    Span4Mux_v I__1491 (
            .O(N__6459),
            .I(N__6449));
    Span4Mux_v I__1490 (
            .O(N__6452),
            .I(N__6446));
    Sp12to4 I__1489 (
            .O(N__6449),
            .I(N__6443));
    Span4Mux_h I__1488 (
            .O(N__6446),
            .I(N__6440));
    Span12Mux_h I__1487 (
            .O(N__6443),
            .I(N__6435));
    Sp12to4 I__1486 (
            .O(N__6440),
            .I(N__6435));
    Odrv12 I__1485 (
            .O(N__6435),
            .I(TEAn_c));
    IoInMux I__1484 (
            .O(N__6432),
            .I(N__6429));
    LocalMux I__1483 (
            .O(N__6429),
            .I(N__6426));
    IoSpan4Mux I__1482 (
            .O(N__6426),
            .I(N__6423));
    Span4Mux_s3_v I__1481 (
            .O(N__6423),
            .I(N__6420));
    Sp12to4 I__1480 (
            .O(N__6420),
            .I(N__6417));
    Span12Mux_v I__1479 (
            .O(N__6417),
            .I(N__6414));
    Odrv12 I__1478 (
            .O(N__6414),
            .I(U111_CYCLE_SM_TEA_CPUn_0_i));
    InMux I__1477 (
            .O(N__6411),
            .I(N__6408));
    LocalMux I__1476 (
            .O(N__6408),
            .I(N__6405));
    Span4Mux_v I__1475 (
            .O(N__6405),
            .I(N__6402));
    Span4Mux_v I__1474 (
            .O(N__6402),
            .I(N__6397));
    InMux I__1473 (
            .O(N__6401),
            .I(N__6394));
    InMux I__1472 (
            .O(N__6400),
            .I(N__6391));
    Span4Mux_v I__1471 (
            .O(N__6397),
            .I(N__6388));
    LocalMux I__1470 (
            .O(N__6394),
            .I(N__6383));
    LocalMux I__1469 (
            .O(N__6391),
            .I(N__6383));
    Sp12to4 I__1468 (
            .O(N__6388),
            .I(N__6378));
    Span12Mux_v I__1467 (
            .O(N__6383),
            .I(N__6378));
    Span12Mux_h I__1466 (
            .O(N__6378),
            .I(N__6375));
    Odrv12 I__1465 (
            .O(N__6375),
            .I(D_UM_AMIGA_in_2));
    InMux I__1464 (
            .O(N__6372),
            .I(N__6369));
    LocalMux I__1463 (
            .O(N__6369),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ));
    InMux I__1462 (
            .O(N__6366),
            .I(N__6362));
    InMux I__1461 (
            .O(N__6365),
            .I(N__6358));
    LocalMux I__1460 (
            .O(N__6362),
            .I(N__6355));
    InMux I__1459 (
            .O(N__6361),
            .I(N__6352));
    LocalMux I__1458 (
            .O(N__6358),
            .I(\U111_CYCLE_SM.un4_TS_OUT_i_0 ));
    Odrv4 I__1457 (
            .O(N__6355),
            .I(\U111_CYCLE_SM.un4_TS_OUT_i_0 ));
    LocalMux I__1456 (
            .O(N__6352),
            .I(\U111_CYCLE_SM.un4_TS_OUT_i_0 ));
    InMux I__1455 (
            .O(N__6345),
            .I(N__6341));
    InMux I__1454 (
            .O(N__6344),
            .I(N__6338));
    LocalMux I__1453 (
            .O(N__6341),
            .I(N__6330));
    LocalMux I__1452 (
            .O(N__6338),
            .I(N__6327));
    InMux I__1451 (
            .O(N__6337),
            .I(N__6324));
    InMux I__1450 (
            .O(N__6336),
            .I(N__6321));
    InMux I__1449 (
            .O(N__6335),
            .I(N__6318));
    InMux I__1448 (
            .O(N__6334),
            .I(N__6313));
    InMux I__1447 (
            .O(N__6333),
            .I(N__6313));
    Odrv4 I__1446 (
            .O(N__6330),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    Odrv4 I__1445 (
            .O(N__6327),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1444 (
            .O(N__6324),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1443 (
            .O(N__6321),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1442 (
            .O(N__6318),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1441 (
            .O(N__6313),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    SRMux I__1440 (
            .O(N__6300),
            .I(N__6276));
    SRMux I__1439 (
            .O(N__6299),
            .I(N__6276));
    SRMux I__1438 (
            .O(N__6298),
            .I(N__6276));
    SRMux I__1437 (
            .O(N__6297),
            .I(N__6276));
    SRMux I__1436 (
            .O(N__6296),
            .I(N__6276));
    SRMux I__1435 (
            .O(N__6295),
            .I(N__6276));
    SRMux I__1434 (
            .O(N__6294),
            .I(N__6276));
    SRMux I__1433 (
            .O(N__6293),
            .I(N__6276));
    GlobalMux I__1432 (
            .O(N__6276),
            .I(N__6273));
    gio2CtrlBuf I__1431 (
            .O(N__6273),
            .I(RESETn_c_i_g));
    InMux I__1430 (
            .O(N__6270),
            .I(N__6264));
    InMux I__1429 (
            .O(N__6269),
            .I(N__6264));
    LocalMux I__1428 (
            .O(N__6264),
            .I(N__6259));
    InMux I__1427 (
            .O(N__6263),
            .I(N__6256));
    InMux I__1426 (
            .O(N__6262),
            .I(N__6249));
    Span4Mux_v I__1425 (
            .O(N__6259),
            .I(N__6244));
    LocalMux I__1424 (
            .O(N__6256),
            .I(N__6244));
    InMux I__1423 (
            .O(N__6255),
            .I(N__6239));
    InMux I__1422 (
            .O(N__6254),
            .I(N__6239));
    InMux I__1421 (
            .O(N__6253),
            .I(N__6234));
    InMux I__1420 (
            .O(N__6252),
            .I(N__6234));
    LocalMux I__1419 (
            .O(N__6249),
            .I(N__6231));
    Span4Mux_h I__1418 (
            .O(N__6244),
            .I(N__6224));
    LocalMux I__1417 (
            .O(N__6239),
            .I(N__6224));
    LocalMux I__1416 (
            .O(N__6234),
            .I(N__6224));
    Span4Mux_v I__1415 (
            .O(N__6231),
            .I(N__6221));
    Span4Mux_v I__1414 (
            .O(N__6224),
            .I(N__6218));
    Span4Mux_h I__1413 (
            .O(N__6221),
            .I(N__6215));
    Span4Mux_h I__1412 (
            .O(N__6218),
            .I(N__6211));
    Span4Mux_h I__1411 (
            .O(N__6215),
            .I(N__6208));
    InMux I__1410 (
            .O(N__6214),
            .I(N__6205));
    Span4Mux_h I__1409 (
            .O(N__6211),
            .I(N__6202));
    Sp12to4 I__1408 (
            .O(N__6208),
            .I(N__6197));
    LocalMux I__1407 (
            .O(N__6205),
            .I(N__6197));
    Sp12to4 I__1406 (
            .O(N__6202),
            .I(N__6192));
    Span12Mux_s7_h I__1405 (
            .O(N__6197),
            .I(N__6192));
    Span12Mux_v I__1404 (
            .O(N__6192),
            .I(N__6189));
    Odrv12 I__1403 (
            .O(N__6189),
            .I(RESETn_c));
    InMux I__1402 (
            .O(N__6186),
            .I(N__6180));
    InMux I__1401 (
            .O(N__6185),
            .I(N__6177));
    InMux I__1400 (
            .O(N__6184),
            .I(N__6174));
    InMux I__1399 (
            .O(N__6183),
            .I(N__6171));
    LocalMux I__1398 (
            .O(N__6180),
            .I(\U111_CYCLE_SM.N_99 ));
    LocalMux I__1397 (
            .O(N__6177),
            .I(\U111_CYCLE_SM.N_99 ));
    LocalMux I__1396 (
            .O(N__6174),
            .I(\U111_CYCLE_SM.N_99 ));
    LocalMux I__1395 (
            .O(N__6171),
            .I(\U111_CYCLE_SM.N_99 ));
    CascadeMux I__1394 (
            .O(N__6162),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81_cascade_ ));
    InMux I__1393 (
            .O(N__6159),
            .I(N__6152));
    InMux I__1392 (
            .O(N__6158),
            .I(N__6139));
    InMux I__1391 (
            .O(N__6157),
            .I(N__6139));
    InMux I__1390 (
            .O(N__6156),
            .I(N__6139));
    InMux I__1389 (
            .O(N__6155),
            .I(N__6139));
    LocalMux I__1388 (
            .O(N__6152),
            .I(N__6136));
    InMux I__1387 (
            .O(N__6151),
            .I(N__6129));
    InMux I__1386 (
            .O(N__6150),
            .I(N__6129));
    InMux I__1385 (
            .O(N__6149),
            .I(N__6129));
    InMux I__1384 (
            .O(N__6148),
            .I(N__6126));
    LocalMux I__1383 (
            .O(N__6139),
            .I(\U111_CYCLE_SM.N_99_i ));
    Odrv4 I__1382 (
            .O(N__6136),
            .I(\U111_CYCLE_SM.N_99_i ));
    LocalMux I__1381 (
            .O(N__6129),
            .I(\U111_CYCLE_SM.N_99_i ));
    LocalMux I__1380 (
            .O(N__6126),
            .I(\U111_CYCLE_SM.N_99_i ));
    InMux I__1379 (
            .O(N__6117),
            .I(N__6114));
    LocalMux I__1378 (
            .O(N__6114),
            .I(N__6111));
    Sp12to4 I__1377 (
            .O(N__6111),
            .I(N__6108));
    Span12Mux_v I__1376 (
            .O(N__6108),
            .I(N__6105));
    Span12Mux_h I__1375 (
            .O(N__6105),
            .I(N__6102));
    Odrv12 I__1374 (
            .O(N__6102),
            .I(D_UM_040_in_1));
    IoInMux I__1373 (
            .O(N__6099),
            .I(N__6095));
    InMux I__1372 (
            .O(N__6098),
            .I(N__6092));
    LocalMux I__1371 (
            .O(N__6095),
            .I(N__6089));
    LocalMux I__1370 (
            .O(N__6092),
            .I(N__6086));
    Span4Mux_s3_h I__1369 (
            .O(N__6089),
            .I(N__6083));
    Span4Mux_v I__1368 (
            .O(N__6086),
            .I(N__6080));
    Sp12to4 I__1367 (
            .O(N__6083),
            .I(N__6077));
    Span4Mux_v I__1366 (
            .O(N__6080),
            .I(N__6074));
    Span12Mux_v I__1365 (
            .O(N__6077),
            .I(N__6071));
    Sp12to4 I__1364 (
            .O(N__6074),
            .I(N__6068));
    Span12Mux_h I__1363 (
            .O(N__6071),
            .I(N__6065));
    Span12Mux_h I__1362 (
            .O(N__6068),
            .I(N__6062));
    Span12Mux_h I__1361 (
            .O(N__6065),
            .I(N__6057));
    Span12Mux_v I__1360 (
            .O(N__6062),
            .I(N__6057));
    Odrv12 I__1359 (
            .O(N__6057),
            .I(D_LL_040_in_1));
    IoInMux I__1358 (
            .O(N__6054),
            .I(N__6051));
    LocalMux I__1357 (
            .O(N__6051),
            .I(N__6048));
    Span12Mux_s4_h I__1356 (
            .O(N__6048),
            .I(N__6045));
    Span12Mux_h I__1355 (
            .O(N__6045),
            .I(N__6042));
    Odrv12 I__1354 (
            .O(N__6042),
            .I(un1_D_UM_040_1));
    CascadeMux I__1353 (
            .O(N__6039),
            .I(N__6035));
    InMux I__1352 (
            .O(N__6038),
            .I(N__6032));
    InMux I__1351 (
            .O(N__6035),
            .I(N__6029));
    LocalMux I__1350 (
            .O(N__6032),
            .I(N__6025));
    LocalMux I__1349 (
            .O(N__6029),
            .I(N__6022));
    InMux I__1348 (
            .O(N__6028),
            .I(N__6019));
    Span4Mux_v I__1347 (
            .O(N__6025),
            .I(N__6016));
    Span4Mux_v I__1346 (
            .O(N__6022),
            .I(N__6011));
    LocalMux I__1345 (
            .O(N__6019),
            .I(N__6011));
    Span4Mux_v I__1344 (
            .O(N__6016),
            .I(N__6008));
    Span4Mux_v I__1343 (
            .O(N__6011),
            .I(N__6005));
    Span4Mux_v I__1342 (
            .O(N__6008),
            .I(N__6000));
    Span4Mux_v I__1341 (
            .O(N__6005),
            .I(N__6000));
    Sp12to4 I__1340 (
            .O(N__6000),
            .I(N__5997));
    Span12Mux_h I__1339 (
            .O(N__5997),
            .I(N__5994));
    Odrv12 I__1338 (
            .O(N__5994),
            .I(D_UU_AMIGA_in_1));
    InMux I__1337 (
            .O(N__5991),
            .I(N__5988));
    LocalMux I__1336 (
            .O(N__5988),
            .I(N__5984));
    InMux I__1335 (
            .O(N__5987),
            .I(N__5981));
    Odrv12 I__1334 (
            .O(N__5984),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ));
    LocalMux I__1333 (
            .O(N__5981),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ));
    IoInMux I__1332 (
            .O(N__5976),
            .I(N__5973));
    LocalMux I__1331 (
            .O(N__5973),
            .I(N__5970));
    Span4Mux_s3_h I__1330 (
            .O(N__5970),
            .I(N__5967));
    Sp12to4 I__1329 (
            .O(N__5967),
            .I(N__5964));
    Span12Mux_v I__1328 (
            .O(N__5964),
            .I(N__5961));
    Span12Mux_h I__1327 (
            .O(N__5961),
            .I(N__5958));
    Odrv12 I__1326 (
            .O(N__5958),
            .I(N_119));
    InMux I__1325 (
            .O(N__5955),
            .I(N__5952));
    LocalMux I__1324 (
            .O(N__5952),
            .I(N__5949));
    Span12Mux_v I__1323 (
            .O(N__5949),
            .I(N__5946));
    Odrv12 I__1322 (
            .O(N__5946),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ));
    InMux I__1321 (
            .O(N__5943),
            .I(N__5939));
    InMux I__1320 (
            .O(N__5942),
            .I(N__5936));
    LocalMux I__1319 (
            .O(N__5939),
            .I(N__5933));
    LocalMux I__1318 (
            .O(N__5936),
            .I(N__5929));
    Span4Mux_h I__1317 (
            .O(N__5933),
            .I(N__5926));
    InMux I__1316 (
            .O(N__5932),
            .I(N__5923));
    Sp12to4 I__1315 (
            .O(N__5929),
            .I(N__5920));
    Span4Mux_v I__1314 (
            .O(N__5926),
            .I(N__5915));
    LocalMux I__1313 (
            .O(N__5923),
            .I(N__5915));
    Span12Mux_v I__1312 (
            .O(N__5920),
            .I(N__5912));
    Sp12to4 I__1311 (
            .O(N__5915),
            .I(N__5909));
    Span12Mux_h I__1310 (
            .O(N__5912),
            .I(N__5906));
    Span12Mux_v I__1309 (
            .O(N__5909),
            .I(N__5903));
    Span12Mux_v I__1308 (
            .O(N__5906),
            .I(N__5900));
    Span12Mux_h I__1307 (
            .O(N__5903),
            .I(N__5897));
    Odrv12 I__1306 (
            .O(N__5900),
            .I(D_UM_AMIGA_in_4));
    Odrv12 I__1305 (
            .O(N__5897),
            .I(D_UM_AMIGA_in_4));
    IoInMux I__1304 (
            .O(N__5892),
            .I(N__5889));
    LocalMux I__1303 (
            .O(N__5889),
            .I(N__5886));
    IoSpan4Mux I__1302 (
            .O(N__5886),
            .I(N__5883));
    IoSpan4Mux I__1301 (
            .O(N__5883),
            .I(N__5880));
    Span4Mux_s2_v I__1300 (
            .O(N__5880),
            .I(N__5877));
    Sp12to4 I__1299 (
            .O(N__5877),
            .I(N__5874));
    Span12Mux_s8_v I__1298 (
            .O(N__5874),
            .I(N__5871));
    Odrv12 I__1297 (
            .O(N__5871),
            .I(un1_D_UM_AMIGA_4));
    InMux I__1296 (
            .O(N__5868),
            .I(N__5865));
    LocalMux I__1295 (
            .O(N__5865),
            .I(N__5862));
    Glb2LocalMux I__1294 (
            .O(N__5862),
            .I(N__5859));
    GlobalMux I__1293 (
            .O(N__5859),
            .I(CLK80));
    IoInMux I__1292 (
            .O(N__5856),
            .I(N__5852));
    IoInMux I__1291 (
            .O(N__5855),
            .I(N__5849));
    LocalMux I__1290 (
            .O(N__5852),
            .I(N__5846));
    LocalMux I__1289 (
            .O(N__5849),
            .I(N__5843));
    Span12Mux_s4_v I__1288 (
            .O(N__5846),
            .I(N__5840));
    Span12Mux_s3_h I__1287 (
            .O(N__5843),
            .I(N__5837));
    Span12Mux_v I__1286 (
            .O(N__5840),
            .I(N__5832));
    Span12Mux_h I__1285 (
            .O(N__5837),
            .I(N__5832));
    Odrv12 I__1284 (
            .O(N__5832),
            .I(GB_BUFFER_CLK80_THRU_CO));
    InMux I__1283 (
            .O(N__5829),
            .I(N__5826));
    LocalMux I__1282 (
            .O(N__5826),
            .I(N__5823));
    Span12Mux_s11_v I__1281 (
            .O(N__5823),
            .I(N__5819));
    InMux I__1280 (
            .O(N__5822),
            .I(N__5816));
    Odrv12 I__1279 (
            .O(N__5819),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ));
    LocalMux I__1278 (
            .O(N__5816),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ));
    InMux I__1277 (
            .O(N__5811),
            .I(N__5807));
    CascadeMux I__1276 (
            .O(N__5810),
            .I(N__5804));
    LocalMux I__1275 (
            .O(N__5807),
            .I(N__5801));
    InMux I__1274 (
            .O(N__5804),
            .I(N__5798));
    Span4Mux_v I__1273 (
            .O(N__5801),
            .I(N__5794));
    LocalMux I__1272 (
            .O(N__5798),
            .I(N__5791));
    InMux I__1271 (
            .O(N__5797),
            .I(N__5788));
    Span4Mux_v I__1270 (
            .O(N__5794),
            .I(N__5785));
    Span4Mux_v I__1269 (
            .O(N__5791),
            .I(N__5782));
    LocalMux I__1268 (
            .O(N__5788),
            .I(N__5779));
    Span4Mux_v I__1267 (
            .O(N__5785),
            .I(N__5776));
    Span4Mux_v I__1266 (
            .O(N__5782),
            .I(N__5771));
    Span4Mux_v I__1265 (
            .O(N__5779),
            .I(N__5771));
    Sp12to4 I__1264 (
            .O(N__5776),
            .I(N__5766));
    Sp12to4 I__1263 (
            .O(N__5771),
            .I(N__5766));
    Span12Mux_h I__1262 (
            .O(N__5766),
            .I(N__5763));
    Odrv12 I__1261 (
            .O(N__5763),
            .I(D_UU_AMIGA_in_0));
    IoInMux I__1260 (
            .O(N__5760),
            .I(N__5757));
    LocalMux I__1259 (
            .O(N__5757),
            .I(N__5754));
    IoSpan4Mux I__1258 (
            .O(N__5754),
            .I(N__5750));
    InMux I__1257 (
            .O(N__5753),
            .I(N__5747));
    Span4Mux_s3_v I__1256 (
            .O(N__5750),
            .I(N__5744));
    LocalMux I__1255 (
            .O(N__5747),
            .I(N__5741));
    Sp12to4 I__1254 (
            .O(N__5744),
            .I(N__5738));
    Span4Mux_v I__1253 (
            .O(N__5741),
            .I(N__5735));
    Span12Mux_v I__1252 (
            .O(N__5738),
            .I(N__5732));
    Span4Mux_v I__1251 (
            .O(N__5735),
            .I(N__5729));
    Odrv12 I__1250 (
            .O(N__5732),
            .I(TS_OUT));
    Odrv4 I__1249 (
            .O(N__5729),
            .I(TS_OUT));
    IoInMux I__1248 (
            .O(N__5724),
            .I(N__5721));
    LocalMux I__1247 (
            .O(N__5721),
            .I(N__5718));
    Span4Mux_s0_v I__1246 (
            .O(N__5718),
            .I(N__5715));
    Span4Mux_v I__1245 (
            .O(N__5715),
            .I(N__5712));
    Span4Mux_v I__1244 (
            .O(N__5712),
            .I(N__5709));
    Odrv4 I__1243 (
            .O(N__5709),
            .I(TSnz));
    IoInMux I__1242 (
            .O(N__5706),
            .I(N__5703));
    LocalMux I__1241 (
            .O(N__5703),
            .I(N__5700));
    IoSpan4Mux I__1240 (
            .O(N__5700),
            .I(N__5696));
    InMux I__1239 (
            .O(N__5699),
            .I(N__5693));
    Span4Mux_s2_h I__1238 (
            .O(N__5696),
            .I(N__5690));
    LocalMux I__1237 (
            .O(N__5693),
            .I(N__5687));
    Sp12to4 I__1236 (
            .O(N__5690),
            .I(N__5684));
    Span4Mux_v I__1235 (
            .O(N__5687),
            .I(N__5681));
    Span12Mux_h I__1234 (
            .O(N__5684),
            .I(N__5678));
    Sp12to4 I__1233 (
            .O(N__5681),
            .I(N__5675));
    Span12Mux_h I__1232 (
            .O(N__5678),
            .I(N__5672));
    Span12Mux_h I__1231 (
            .O(N__5675),
            .I(N__5669));
    Odrv12 I__1230 (
            .O(N__5672),
            .I(D_LM_040_in_7));
    Odrv12 I__1229 (
            .O(N__5669),
            .I(D_LM_040_in_7));
    InMux I__1228 (
            .O(N__5664),
            .I(N__5661));
    LocalMux I__1227 (
            .O(N__5661),
            .I(N__5658));
    Span4Mux_v I__1226 (
            .O(N__5658),
            .I(N__5655));
    Sp12to4 I__1225 (
            .O(N__5655),
            .I(N__5652));
    Span12Mux_h I__1224 (
            .O(N__5652),
            .I(N__5649));
    Odrv12 I__1223 (
            .O(N__5649),
            .I(D_UU_040_in_7));
    IoInMux I__1222 (
            .O(N__5646),
            .I(N__5643));
    LocalMux I__1221 (
            .O(N__5643),
            .I(N__5640));
    Span12Mux_s9_v I__1220 (
            .O(N__5640),
            .I(N__5637));
    Span12Mux_h I__1219 (
            .O(N__5637),
            .I(N__5634));
    Odrv12 I__1218 (
            .O(N__5634),
            .I(un1_D_UU_040_7));
    InMux I__1217 (
            .O(N__5631),
            .I(N__5628));
    LocalMux I__1216 (
            .O(N__5628),
            .I(N__5625));
    Sp12to4 I__1215 (
            .O(N__5625),
            .I(N__5621));
    InMux I__1214 (
            .O(N__5624),
            .I(N__5618));
    Odrv12 I__1213 (
            .O(N__5621),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ));
    LocalMux I__1212 (
            .O(N__5618),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ));
    InMux I__1211 (
            .O(N__5613),
            .I(N__5610));
    LocalMux I__1210 (
            .O(N__5610),
            .I(N__5606));
    CascadeMux I__1209 (
            .O(N__5609),
            .I(N__5603));
    Span4Mux_v I__1208 (
            .O(N__5606),
            .I(N__5599));
    InMux I__1207 (
            .O(N__5603),
            .I(N__5596));
    InMux I__1206 (
            .O(N__5602),
            .I(N__5593));
    Span4Mux_v I__1205 (
            .O(N__5599),
            .I(N__5590));
    LocalMux I__1204 (
            .O(N__5596),
            .I(N__5585));
    LocalMux I__1203 (
            .O(N__5593),
            .I(N__5585));
    Sp12to4 I__1202 (
            .O(N__5590),
            .I(N__5580));
    Span12Mux_v I__1201 (
            .O(N__5585),
            .I(N__5580));
    Span12Mux_h I__1200 (
            .O(N__5580),
            .I(N__5577));
    Odrv12 I__1199 (
            .O(N__5577),
            .I(D_UU_AMIGA_in_6));
    IoInMux I__1198 (
            .O(N__5574),
            .I(N__5571));
    LocalMux I__1197 (
            .O(N__5571),
            .I(N__5568));
    Span4Mux_s3_v I__1196 (
            .O(N__5568),
            .I(N__5565));
    Span4Mux_h I__1195 (
            .O(N__5565),
            .I(N__5562));
    Span4Mux_h I__1194 (
            .O(N__5562),
            .I(N__5559));
    Span4Mux_h I__1193 (
            .O(N__5559),
            .I(N__5556));
    Odrv4 I__1192 (
            .O(N__5556),
            .I(N_114));
    IoInMux I__1191 (
            .O(N__5553),
            .I(N__5550));
    LocalMux I__1190 (
            .O(N__5550),
            .I(N__5547));
    Span4Mux_s2_v I__1189 (
            .O(N__5547),
            .I(N__5544));
    Span4Mux_v I__1188 (
            .O(N__5544),
            .I(N__5541));
    Odrv4 I__1187 (
            .O(N__5541),
            .I(CONSTANT_ONE_NET));
    InMux I__1186 (
            .O(N__5538),
            .I(N__5534));
    InMux I__1185 (
            .O(N__5537),
            .I(N__5531));
    LocalMux I__1184 (
            .O(N__5534),
            .I(N__5526));
    LocalMux I__1183 (
            .O(N__5531),
            .I(N__5526));
    Span4Mux_v I__1182 (
            .O(N__5526),
            .I(N__5523));
    Sp12to4 I__1181 (
            .O(N__5523),
            .I(N__5520));
    Span12Mux_h I__1180 (
            .O(N__5520),
            .I(N__5517));
    Odrv12 I__1179 (
            .O(N__5517),
            .I(BGn_c));
    CascadeMux I__1178 (
            .O(N__5514),
            .I(N__5511));
    InMux I__1177 (
            .O(N__5511),
            .I(N__5508));
    LocalMux I__1176 (
            .O(N__5508),
            .I(N__5505));
    Span4Mux_v I__1175 (
            .O(N__5505),
            .I(N__5500));
    InMux I__1174 (
            .O(N__5504),
            .I(N__5497));
    InMux I__1173 (
            .O(N__5503),
            .I(N__5494));
    Odrv4 I__1172 (
            .O(N__5500),
            .I(\U111_CYCLE_SM.CYCLE_ENZ0 ));
    LocalMux I__1171 (
            .O(N__5497),
            .I(\U111_CYCLE_SM.CYCLE_ENZ0 ));
    LocalMux I__1170 (
            .O(N__5494),
            .I(\U111_CYCLE_SM.CYCLE_ENZ0 ));
    InMux I__1169 (
            .O(N__5487),
            .I(N__5483));
    InMux I__1168 (
            .O(N__5486),
            .I(N__5480));
    LocalMux I__1167 (
            .O(N__5483),
            .I(\U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0 ));
    LocalMux I__1166 (
            .O(N__5480),
            .I(\U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0 ));
    IoInMux I__1165 (
            .O(N__5475),
            .I(N__5472));
    LocalMux I__1164 (
            .O(N__5472),
            .I(N__5469));
    IoSpan4Mux I__1163 (
            .O(N__5469),
            .I(N__5458));
    IoInMux I__1162 (
            .O(N__5468),
            .I(N__5454));
    IoInMux I__1161 (
            .O(N__5467),
            .I(N__5451));
    IoInMux I__1160 (
            .O(N__5466),
            .I(N__5448));
    IoInMux I__1159 (
            .O(N__5465),
            .I(N__5445));
    IoInMux I__1158 (
            .O(N__5464),
            .I(N__5442));
    IoInMux I__1157 (
            .O(N__5463),
            .I(N__5439));
    IoInMux I__1156 (
            .O(N__5462),
            .I(N__5436));
    IoInMux I__1155 (
            .O(N__5461),
            .I(N__5427));
    Span4Mux_s3_h I__1154 (
            .O(N__5458),
            .I(N__5424));
    IoInMux I__1153 (
            .O(N__5457),
            .I(N__5421));
    LocalMux I__1152 (
            .O(N__5454),
            .I(N__5408));
    LocalMux I__1151 (
            .O(N__5451),
            .I(N__5408));
    LocalMux I__1150 (
            .O(N__5448),
            .I(N__5408));
    LocalMux I__1149 (
            .O(N__5445),
            .I(N__5408));
    LocalMux I__1148 (
            .O(N__5442),
            .I(N__5408));
    LocalMux I__1147 (
            .O(N__5439),
            .I(N__5408));
    LocalMux I__1146 (
            .O(N__5436),
            .I(N__5405));
    IoInMux I__1145 (
            .O(N__5435),
            .I(N__5402));
    IoInMux I__1144 (
            .O(N__5434),
            .I(N__5399));
    IoInMux I__1143 (
            .O(N__5433),
            .I(N__5392));
    IoInMux I__1142 (
            .O(N__5432),
            .I(N__5389));
    IoInMux I__1141 (
            .O(N__5431),
            .I(N__5386));
    IoInMux I__1140 (
            .O(N__5430),
            .I(N__5383));
    LocalMux I__1139 (
            .O(N__5427),
            .I(N__5374));
    IoSpan4Mux I__1138 (
            .O(N__5424),
            .I(N__5374));
    LocalMux I__1137 (
            .O(N__5421),
            .I(N__5374));
    IoSpan4Mux I__1136 (
            .O(N__5408),
            .I(N__5374));
    IoSpan4Mux I__1135 (
            .O(N__5405),
            .I(N__5363));
    LocalMux I__1134 (
            .O(N__5402),
            .I(N__5363));
    LocalMux I__1133 (
            .O(N__5399),
            .I(N__5363));
    IoInMux I__1132 (
            .O(N__5398),
            .I(N__5360));
    IoInMux I__1131 (
            .O(N__5397),
            .I(N__5357));
    IoInMux I__1130 (
            .O(N__5396),
            .I(N__5354));
    IoInMux I__1129 (
            .O(N__5395),
            .I(N__5351));
    LocalMux I__1128 (
            .O(N__5392),
            .I(N__5340));
    LocalMux I__1127 (
            .O(N__5389),
            .I(N__5340));
    LocalMux I__1126 (
            .O(N__5386),
            .I(N__5340));
    LocalMux I__1125 (
            .O(N__5383),
            .I(N__5340));
    IoSpan4Mux I__1124 (
            .O(N__5374),
            .I(N__5340));
    IoInMux I__1123 (
            .O(N__5373),
            .I(N__5337));
    IoInMux I__1122 (
            .O(N__5372),
            .I(N__5334));
    IoInMux I__1121 (
            .O(N__5371),
            .I(N__5331));
    IoInMux I__1120 (
            .O(N__5370),
            .I(N__5328));
    IoSpan4Mux I__1119 (
            .O(N__5363),
            .I(N__5312));
    LocalMux I__1118 (
            .O(N__5360),
            .I(N__5312));
    LocalMux I__1117 (
            .O(N__5357),
            .I(N__5312));
    LocalMux I__1116 (
            .O(N__5354),
            .I(N__5312));
    LocalMux I__1115 (
            .O(N__5351),
            .I(N__5312));
    IoSpan4Mux I__1114 (
            .O(N__5340),
            .I(N__5301));
    LocalMux I__1113 (
            .O(N__5337),
            .I(N__5301));
    LocalMux I__1112 (
            .O(N__5334),
            .I(N__5301));
    LocalMux I__1111 (
            .O(N__5331),
            .I(N__5301));
    LocalMux I__1110 (
            .O(N__5328),
            .I(N__5301));
    IoInMux I__1109 (
            .O(N__5327),
            .I(N__5298));
    IoInMux I__1108 (
            .O(N__5326),
            .I(N__5295));
    IoInMux I__1107 (
            .O(N__5325),
            .I(N__5292));
    IoInMux I__1106 (
            .O(N__5324),
            .I(N__5289));
    IoInMux I__1105 (
            .O(N__5323),
            .I(N__5286));
    IoSpan4Mux I__1104 (
            .O(N__5312),
            .I(N__5281));
    IoSpan4Mux I__1103 (
            .O(N__5301),
            .I(N__5270));
    LocalMux I__1102 (
            .O(N__5298),
            .I(N__5270));
    LocalMux I__1101 (
            .O(N__5295),
            .I(N__5270));
    LocalMux I__1100 (
            .O(N__5292),
            .I(N__5270));
    LocalMux I__1099 (
            .O(N__5289),
            .I(N__5270));
    LocalMux I__1098 (
            .O(N__5286),
            .I(N__5267));
    IoInMux I__1097 (
            .O(N__5285),
            .I(N__5263));
    IoInMux I__1096 (
            .O(N__5284),
            .I(N__5260));
    Span4Mux_s3_h I__1095 (
            .O(N__5281),
            .I(N__5257));
    IoSpan4Mux I__1094 (
            .O(N__5270),
            .I(N__5252));
    IoSpan4Mux I__1093 (
            .O(N__5267),
            .I(N__5252));
    IoInMux I__1092 (
            .O(N__5266),
            .I(N__5249));
    LocalMux I__1091 (
            .O(N__5263),
            .I(N__5244));
    LocalMux I__1090 (
            .O(N__5260),
            .I(N__5244));
    Span4Mux_v I__1089 (
            .O(N__5257),
            .I(N__5239));
    Span4Mux_s3_h I__1088 (
            .O(N__5252),
            .I(N__5239));
    LocalMux I__1087 (
            .O(N__5249),
            .I(N__5236));
    Span12Mux_s4_h I__1086 (
            .O(N__5244),
            .I(N__5233));
    Sp12to4 I__1085 (
            .O(N__5239),
            .I(N__5228));
    Span12Mux_s4_h I__1084 (
            .O(N__5236),
            .I(N__5228));
    Span12Mux_h I__1083 (
            .O(N__5233),
            .I(N__5223));
    Span12Mux_h I__1082 (
            .O(N__5228),
            .I(N__5223));
    Odrv12 I__1081 (
            .O(N__5223),
            .I(U111_CYCLE_SM_OFFBOARD_EN_0));
    InMux I__1080 (
            .O(N__5220),
            .I(N__5216));
    InMux I__1079 (
            .O(N__5219),
            .I(N__5213));
    LocalMux I__1078 (
            .O(N__5216),
            .I(\U111_CYCLE_SM.TS_DELAYZ0 ));
    LocalMux I__1077 (
            .O(N__5213),
            .I(\U111_CYCLE_SM.TS_DELAYZ0 ));
    CascadeMux I__1076 (
            .O(N__5208),
            .I(\U111_CYCLE_SM.un4_TS_OUT_i_0_cascade_ ));
    IoInMux I__1075 (
            .O(N__5205),
            .I(N__5202));
    LocalMux I__1074 (
            .O(N__5202),
            .I(N__5199));
    Span4Mux_s1_v I__1073 (
            .O(N__5199),
            .I(N__5196));
    Span4Mux_h I__1072 (
            .O(N__5196),
            .I(N__5193));
    Span4Mux_v I__1071 (
            .O(N__5193),
            .I(N__5190));
    Span4Mux_v I__1070 (
            .O(N__5190),
            .I(N__5186));
    InMux I__1069 (
            .O(N__5189),
            .I(N__5183));
    Span4Mux_v I__1068 (
            .O(N__5186),
            .I(N__5176));
    LocalMux I__1067 (
            .O(N__5183),
            .I(N__5176));
    InMux I__1066 (
            .O(N__5182),
            .I(N__5173));
    InMux I__1065 (
            .O(N__5181),
            .I(N__5170));
    Span4Mux_v I__1064 (
            .O(N__5176),
            .I(N__5163));
    LocalMux I__1063 (
            .O(N__5173),
            .I(N__5163));
    LocalMux I__1062 (
            .O(N__5170),
            .I(N__5163));
    Span4Mux_v I__1061 (
            .O(N__5163),
            .I(N__5159));
    CascadeMux I__1060 (
            .O(N__5162),
            .I(N__5155));
    Sp12to4 I__1059 (
            .O(N__5159),
            .I(N__5151));
    InMux I__1058 (
            .O(N__5158),
            .I(N__5146));
    InMux I__1057 (
            .O(N__5155),
            .I(N__5146));
    InMux I__1056 (
            .O(N__5154),
            .I(N__5143));
    Span12Mux_h I__1055 (
            .O(N__5151),
            .I(N__5136));
    LocalMux I__1054 (
            .O(N__5146),
            .I(N__5136));
    LocalMux I__1053 (
            .O(N__5143),
            .I(N__5136));
    Span12Mux_v I__1052 (
            .O(N__5136),
            .I(N__5133));
    Odrv12 I__1051 (
            .O(N__5133),
            .I(TACKn_in));
    InMux I__1050 (
            .O(N__5130),
            .I(N__5123));
    InMux I__1049 (
            .O(N__5129),
            .I(N__5120));
    InMux I__1048 (
            .O(N__5128),
            .I(N__5115));
    InMux I__1047 (
            .O(N__5127),
            .I(N__5115));
    InMux I__1046 (
            .O(N__5126),
            .I(N__5112));
    LocalMux I__1045 (
            .O(N__5123),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ));
    LocalMux I__1044 (
            .O(N__5120),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ));
    LocalMux I__1043 (
            .O(N__5115),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ));
    LocalMux I__1042 (
            .O(N__5112),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ));
    CascadeMux I__1041 (
            .O(N__5103),
            .I(\U111_CYCLE_SM.N_99_cascade_ ));
    CascadeMux I__1040 (
            .O(N__5100),
            .I(N__5097));
    InMux I__1039 (
            .O(N__5097),
            .I(N__5088));
    InMux I__1038 (
            .O(N__5096),
            .I(N__5088));
    InMux I__1037 (
            .O(N__5095),
            .I(N__5085));
    InMux I__1036 (
            .O(N__5094),
            .I(N__5081));
    InMux I__1035 (
            .O(N__5093),
            .I(N__5078));
    LocalMux I__1034 (
            .O(N__5088),
            .I(N__5075));
    LocalMux I__1033 (
            .O(N__5085),
            .I(N__5072));
    InMux I__1032 (
            .O(N__5084),
            .I(N__5069));
    LocalMux I__1031 (
            .O(N__5081),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    LocalMux I__1030 (
            .O(N__5078),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    Odrv4 I__1029 (
            .O(N__5075),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    Odrv4 I__1028 (
            .O(N__5072),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    LocalMux I__1027 (
            .O(N__5069),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    InMux I__1026 (
            .O(N__5058),
            .I(N__5055));
    LocalMux I__1025 (
            .O(N__5055),
            .I(\U111_CYCLE_SM.N_51 ));
    CascadeMux I__1024 (
            .O(N__5052),
            .I(N__5045));
    InMux I__1023 (
            .O(N__5051),
            .I(N__5040));
    InMux I__1022 (
            .O(N__5050),
            .I(N__5037));
    InMux I__1021 (
            .O(N__5049),
            .I(N__5026));
    InMux I__1020 (
            .O(N__5048),
            .I(N__5026));
    InMux I__1019 (
            .O(N__5045),
            .I(N__5026));
    InMux I__1018 (
            .O(N__5044),
            .I(N__5026));
    InMux I__1017 (
            .O(N__5043),
            .I(N__5026));
    LocalMux I__1016 (
            .O(N__5040),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    LocalMux I__1015 (
            .O(N__5037),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    LocalMux I__1014 (
            .O(N__5026),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    IoInMux I__1013 (
            .O(N__5019),
            .I(N__5016));
    LocalMux I__1012 (
            .O(N__5016),
            .I(N__5013));
    Span4Mux_s3_h I__1011 (
            .O(N__5013),
            .I(N__5009));
    InMux I__1010 (
            .O(N__5012),
            .I(N__5006));
    Sp12to4 I__1009 (
            .O(N__5009),
            .I(N__5003));
    LocalMux I__1008 (
            .O(N__5006),
            .I(N__5000));
    Span12Mux_v I__1007 (
            .O(N__5003),
            .I(N__4997));
    Span12Mux_v I__1006 (
            .O(N__5000),
            .I(N__4994));
    Span12Mux_h I__1005 (
            .O(N__4997),
            .I(N__4989));
    Span12Mux_v I__1004 (
            .O(N__4994),
            .I(N__4989));
    Span12Mux_h I__1003 (
            .O(N__4989),
            .I(N__4986));
    Odrv12 I__1002 (
            .O(N__4986),
            .I(D_LM_040_in_1));
    InMux I__1001 (
            .O(N__4983),
            .I(N__4980));
    LocalMux I__1000 (
            .O(N__4980),
            .I(N__4977));
    Span12Mux_v I__999 (
            .O(N__4977),
            .I(N__4974));
    Span12Mux_h I__998 (
            .O(N__4974),
            .I(N__4971));
    Odrv12 I__997 (
            .O(N__4971),
            .I(D_UU_040_in_1));
    IoInMux I__996 (
            .O(N__4968),
            .I(N__4965));
    LocalMux I__995 (
            .O(N__4965),
            .I(N__4962));
    IoSpan4Mux I__994 (
            .O(N__4962),
            .I(N__4959));
    Span4Mux_s0_h I__993 (
            .O(N__4959),
            .I(N__4956));
    Sp12to4 I__992 (
            .O(N__4956),
            .I(N__4953));
    Span12Mux_s11_h I__991 (
            .O(N__4953),
            .I(N__4950));
    Odrv12 I__990 (
            .O(N__4950),
            .I(un1_D_UU_040_1));
    InMux I__989 (
            .O(N__4947),
            .I(N__4944));
    LocalMux I__988 (
            .O(N__4944),
            .I(N__4941));
    Span4Mux_v I__987 (
            .O(N__4941),
            .I(N__4938));
    Span4Mux_v I__986 (
            .O(N__4938),
            .I(N__4934));
    InMux I__985 (
            .O(N__4937),
            .I(N__4931));
    Odrv4 I__984 (
            .O(N__4934),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ));
    LocalMux I__983 (
            .O(N__4931),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ));
    IoInMux I__982 (
            .O(N__4926),
            .I(N__4923));
    LocalMux I__981 (
            .O(N__4923),
            .I(N__4920));
    Span4Mux_s2_v I__980 (
            .O(N__4920),
            .I(N__4917));
    Span4Mux_h I__979 (
            .O(N__4917),
            .I(N__4914));
    Span4Mux_v I__978 (
            .O(N__4914),
            .I(N__4911));
    Sp12to4 I__977 (
            .O(N__4911),
            .I(N__4908));
    Odrv12 I__976 (
            .O(N__4908),
            .I(N_115));
    CascadeMux I__975 (
            .O(N__4905),
            .I(\U111_CYCLE_SM.CYCLE_STATE_srsts_i_i_o2_0_5_cascade_ ));
    InMux I__974 (
            .O(N__4902),
            .I(N__4899));
    LocalMux I__973 (
            .O(N__4899),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ));
    CascadeMux I__972 (
            .O(N__4896),
            .I(N__4893));
    InMux I__971 (
            .O(N__4893),
            .I(N__4887));
    InMux I__970 (
            .O(N__4892),
            .I(N__4884));
    InMux I__969 (
            .O(N__4891),
            .I(N__4879));
    InMux I__968 (
            .O(N__4890),
            .I(N__4879));
    LocalMux I__967 (
            .O(N__4887),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    LocalMux I__966 (
            .O(N__4884),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    LocalMux I__965 (
            .O(N__4879),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    InMux I__964 (
            .O(N__4872),
            .I(N__4866));
    InMux I__963 (
            .O(N__4871),
            .I(N__4863));
    InMux I__962 (
            .O(N__4870),
            .I(N__4858));
    InMux I__961 (
            .O(N__4869),
            .I(N__4858));
    LocalMux I__960 (
            .O(N__4866),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    LocalMux I__959 (
            .O(N__4863),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    LocalMux I__958 (
            .O(N__4858),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    InMux I__957 (
            .O(N__4851),
            .I(N__4843));
    InMux I__956 (
            .O(N__4850),
            .I(N__4840));
    InMux I__955 (
            .O(N__4849),
            .I(N__4837));
    InMux I__954 (
            .O(N__4848),
            .I(N__4834));
    InMux I__953 (
            .O(N__4847),
            .I(N__4829));
    InMux I__952 (
            .O(N__4846),
            .I(N__4829));
    LocalMux I__951 (
            .O(N__4843),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    LocalMux I__950 (
            .O(N__4840),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    LocalMux I__949 (
            .O(N__4837),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    LocalMux I__948 (
            .O(N__4834),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    LocalMux I__947 (
            .O(N__4829),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    CascadeMux I__946 (
            .O(N__4818),
            .I(\U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_a3_2_0_0_cascade_ ));
    InMux I__945 (
            .O(N__4815),
            .I(N__4812));
    LocalMux I__944 (
            .O(N__4812),
            .I(\U111_CYCLE_SM.N_133 ));
    InMux I__943 (
            .O(N__4809),
            .I(N__4806));
    LocalMux I__942 (
            .O(N__4806),
            .I(\U111_CYCLE_SM.N_131 ));
    CascadeMux I__941 (
            .O(N__4803),
            .I(\U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_2_0_cascade_ ));
    InMux I__940 (
            .O(N__4800),
            .I(N__4797));
    LocalMux I__939 (
            .O(N__4797),
            .I(N__4794));
    Span4Mux_h I__938 (
            .O(N__4794),
            .I(N__4791));
    Sp12to4 I__937 (
            .O(N__4791),
            .I(N__4788));
    Span12Mux_v I__936 (
            .O(N__4788),
            .I(N__4785));
    Odrv12 I__935 (
            .O(N__4785),
            .I(TS_CPUn_in));
    InMux I__934 (
            .O(N__4782),
            .I(N__4779));
    LocalMux I__933 (
            .O(N__4779),
            .I(N__4776));
    Span4Mux_v I__932 (
            .O(N__4776),
            .I(N__4773));
    Sp12to4 I__931 (
            .O(N__4773),
            .I(N__4770));
    Span12Mux_h I__930 (
            .O(N__4770),
            .I(N__4767));
    Odrv12 I__929 (
            .O(N__4767),
            .I(D_LM_AMIGA_in_4));
    IoInMux I__928 (
            .O(N__4764),
            .I(N__4761));
    LocalMux I__927 (
            .O(N__4761),
            .I(N__4758));
    IoSpan4Mux I__926 (
            .O(N__4758),
            .I(N__4755));
    Span4Mux_s3_h I__925 (
            .O(N__4755),
            .I(N__4752));
    Sp12to4 I__924 (
            .O(N__4752),
            .I(N__4749));
    Span12Mux_h I__923 (
            .O(N__4749),
            .I(N__4746));
    Odrv12 I__922 (
            .O(N__4746),
            .I(N_109));
    InMux I__921 (
            .O(N__4743),
            .I(N__4740));
    LocalMux I__920 (
            .O(N__4740),
            .I(N__4737));
    Span4Mux_v I__919 (
            .O(N__4737),
            .I(N__4734));
    Sp12to4 I__918 (
            .O(N__4734),
            .I(N__4731));
    Span12Mux_h I__917 (
            .O(N__4731),
            .I(N__4728));
    Odrv12 I__916 (
            .O(N__4728),
            .I(D_UU_040_in_2));
    IoInMux I__915 (
            .O(N__4725),
            .I(N__4721));
    InMux I__914 (
            .O(N__4724),
            .I(N__4718));
    LocalMux I__913 (
            .O(N__4721),
            .I(N__4715));
    LocalMux I__912 (
            .O(N__4718),
            .I(N__4712));
    Span4Mux_s2_h I__911 (
            .O(N__4715),
            .I(N__4709));
    Span4Mux_h I__910 (
            .O(N__4712),
            .I(N__4706));
    Sp12to4 I__909 (
            .O(N__4709),
            .I(N__4703));
    Sp12to4 I__908 (
            .O(N__4706),
            .I(N__4700));
    Span12Mux_h I__907 (
            .O(N__4703),
            .I(N__4697));
    Span12Mux_v I__906 (
            .O(N__4700),
            .I(N__4694));
    Span12Mux_h I__905 (
            .O(N__4697),
            .I(N__4691));
    Span12Mux_v I__904 (
            .O(N__4694),
            .I(N__4688));
    Span12Mux_v I__903 (
            .O(N__4691),
            .I(N__4685));
    Span12Mux_h I__902 (
            .O(N__4688),
            .I(N__4682));
    Odrv12 I__901 (
            .O(N__4685),
            .I(D_LM_040_in_2));
    Odrv12 I__900 (
            .O(N__4682),
            .I(D_LM_040_in_2));
    IoInMux I__899 (
            .O(N__4677),
            .I(N__4674));
    LocalMux I__898 (
            .O(N__4674),
            .I(N__4671));
    Span4Mux_s2_v I__897 (
            .O(N__4671),
            .I(N__4668));
    Span4Mux_h I__896 (
            .O(N__4668),
            .I(N__4665));
    Span4Mux_h I__895 (
            .O(N__4665),
            .I(N__4662));
    Span4Mux_v I__894 (
            .O(N__4662),
            .I(N__4659));
    Odrv4 I__893 (
            .O(N__4659),
            .I(un1_D_UU_040_2));
    InMux I__892 (
            .O(N__4656),
            .I(N__4653));
    LocalMux I__891 (
            .O(N__4653),
            .I(N__4649));
    CascadeMux I__890 (
            .O(N__4652),
            .I(N__4645));
    Span4Mux_v I__889 (
            .O(N__4649),
            .I(N__4642));
    InMux I__888 (
            .O(N__4648),
            .I(N__4639));
    InMux I__887 (
            .O(N__4645),
            .I(N__4636));
    Span4Mux_v I__886 (
            .O(N__4642),
            .I(N__4633));
    LocalMux I__885 (
            .O(N__4639),
            .I(N__4630));
    LocalMux I__884 (
            .O(N__4636),
            .I(N__4627));
    Span4Mux_v I__883 (
            .O(N__4633),
            .I(N__4624));
    Span4Mux_v I__882 (
            .O(N__4630),
            .I(N__4621));
    Span12Mux_h I__881 (
            .O(N__4627),
            .I(N__4618));
    Sp12to4 I__880 (
            .O(N__4624),
            .I(N__4613));
    Sp12to4 I__879 (
            .O(N__4621),
            .I(N__4613));
    Span12Mux_v I__878 (
            .O(N__4618),
            .I(N__4608));
    Span12Mux_h I__877 (
            .O(N__4613),
            .I(N__4608));
    Odrv12 I__876 (
            .O(N__4608),
            .I(D_UU_AMIGA_in_2));
    InMux I__875 (
            .O(N__4605),
            .I(N__4602));
    LocalMux I__874 (
            .O(N__4602),
            .I(N__4598));
    InMux I__873 (
            .O(N__4601),
            .I(N__4595));
    Odrv12 I__872 (
            .O(N__4598),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ));
    LocalMux I__871 (
            .O(N__4595),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ));
    IoInMux I__870 (
            .O(N__4590),
            .I(N__4587));
    LocalMux I__869 (
            .O(N__4587),
            .I(N__4584));
    Span12Mux_s8_v I__868 (
            .O(N__4584),
            .I(N__4581));
    Span12Mux_h I__867 (
            .O(N__4581),
            .I(N__4578));
    Odrv12 I__866 (
            .O(N__4578),
            .I(N_118));
    InMux I__865 (
            .O(N__4575),
            .I(N__4572));
    LocalMux I__864 (
            .O(N__4572),
            .I(N__4569));
    Span12Mux_s8_v I__863 (
            .O(N__4569),
            .I(N__4565));
    InMux I__862 (
            .O(N__4568),
            .I(N__4562));
    Odrv12 I__861 (
            .O(N__4565),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ));
    LocalMux I__860 (
            .O(N__4562),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ));
    CascadeMux I__859 (
            .O(N__4557),
            .I(N__4554));
    InMux I__858 (
            .O(N__4554),
            .I(N__4551));
    LocalMux I__857 (
            .O(N__4551),
            .I(N__4547));
    InMux I__856 (
            .O(N__4550),
            .I(N__4544));
    Span4Mux_h I__855 (
            .O(N__4547),
            .I(N__4539));
    LocalMux I__854 (
            .O(N__4544),
            .I(N__4539));
    Span4Mux_v I__853 (
            .O(N__4539),
            .I(N__4535));
    InMux I__852 (
            .O(N__4538),
            .I(N__4532));
    Span4Mux_v I__851 (
            .O(N__4535),
            .I(N__4527));
    LocalMux I__850 (
            .O(N__4532),
            .I(N__4527));
    Span4Mux_v I__849 (
            .O(N__4527),
            .I(N__4524));
    IoSpan4Mux I__848 (
            .O(N__4524),
            .I(N__4521));
    IoSpan4Mux I__847 (
            .O(N__4521),
            .I(N__4518));
    Odrv4 I__846 (
            .O(N__4518),
            .I(D_UU_AMIGA_in_4));
    IoInMux I__845 (
            .O(N__4515),
            .I(N__4512));
    LocalMux I__844 (
            .O(N__4512),
            .I(N__4509));
    Span4Mux_s2_v I__843 (
            .O(N__4509),
            .I(N__4506));
    Span4Mux_h I__842 (
            .O(N__4506),
            .I(N__4503));
    Span4Mux_h I__841 (
            .O(N__4503),
            .I(N__4500));
    Span4Mux_v I__840 (
            .O(N__4500),
            .I(N__4497));
    Odrv4 I__839 (
            .O(N__4497),
            .I(N_116));
    CascadeMux I__838 (
            .O(N__4494),
            .I(N__4490));
    InMux I__837 (
            .O(N__4493),
            .I(N__4487));
    InMux I__836 (
            .O(N__4490),
            .I(N__4483));
    LocalMux I__835 (
            .O(N__4487),
            .I(N__4480));
    InMux I__834 (
            .O(N__4486),
            .I(N__4477));
    LocalMux I__833 (
            .O(N__4483),
            .I(N__4474));
    Span4Mux_v I__832 (
            .O(N__4480),
            .I(N__4469));
    LocalMux I__831 (
            .O(N__4477),
            .I(N__4469));
    Sp12to4 I__830 (
            .O(N__4474),
            .I(N__4466));
    Span4Mux_v I__829 (
            .O(N__4469),
            .I(N__4463));
    Span12Mux_v I__828 (
            .O(N__4466),
            .I(N__4458));
    Sp12to4 I__827 (
            .O(N__4463),
            .I(N__4458));
    Span12Mux_h I__826 (
            .O(N__4458),
            .I(N__4455));
    Odrv12 I__825 (
            .O(N__4455),
            .I(D_UU_AMIGA_in_7));
    InMux I__824 (
            .O(N__4452),
            .I(N__4449));
    LocalMux I__823 (
            .O(N__4449),
            .I(N__4446));
    Span12Mux_v I__822 (
            .O(N__4446),
            .I(N__4442));
    InMux I__821 (
            .O(N__4445),
            .I(N__4439));
    Odrv12 I__820 (
            .O(N__4442),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ));
    LocalMux I__819 (
            .O(N__4439),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ));
    IoInMux I__818 (
            .O(N__4434),
            .I(N__4431));
    LocalMux I__817 (
            .O(N__4431),
            .I(N__4428));
    IoSpan4Mux I__816 (
            .O(N__4428),
            .I(N__4425));
    Span4Mux_s2_v I__815 (
            .O(N__4425),
            .I(N__4422));
    Span4Mux_v I__814 (
            .O(N__4422),
            .I(N__4419));
    Sp12to4 I__813 (
            .O(N__4419),
            .I(N__4416));
    Odrv12 I__812 (
            .O(N__4416),
            .I(N_113));
    IoInMux I__811 (
            .O(N__4413),
            .I(N__4410));
    LocalMux I__810 (
            .O(N__4410),
            .I(N__4407));
    IoSpan4Mux I__809 (
            .O(N__4407),
            .I(N__4403));
    InMux I__808 (
            .O(N__4406),
            .I(N__4400));
    IoSpan4Mux I__807 (
            .O(N__4403),
            .I(N__4397));
    LocalMux I__806 (
            .O(N__4400),
            .I(N__4394));
    Span4Mux_s2_h I__805 (
            .O(N__4397),
            .I(N__4391));
    Span4Mux_v I__804 (
            .O(N__4394),
            .I(N__4388));
    Sp12to4 I__803 (
            .O(N__4391),
            .I(N__4385));
    Sp12to4 I__802 (
            .O(N__4388),
            .I(N__4382));
    Span12Mux_h I__801 (
            .O(N__4385),
            .I(N__4379));
    Span12Mux_h I__800 (
            .O(N__4382),
            .I(N__4376));
    Span12Mux_h I__799 (
            .O(N__4379),
            .I(N__4373));
    Span12Mux_v I__798 (
            .O(N__4376),
            .I(N__4370));
    Odrv12 I__797 (
            .O(N__4373),
            .I(D_LM_040_in_3));
    Odrv12 I__796 (
            .O(N__4370),
            .I(D_LM_040_in_3));
    InMux I__795 (
            .O(N__4365),
            .I(N__4362));
    LocalMux I__794 (
            .O(N__4362),
            .I(N__4359));
    Span4Mux_v I__793 (
            .O(N__4359),
            .I(N__4356));
    Span4Mux_h I__792 (
            .O(N__4356),
            .I(N__4353));
    Sp12to4 I__791 (
            .O(N__4353),
            .I(N__4350));
    Span12Mux_h I__790 (
            .O(N__4350),
            .I(N__4347));
    Odrv12 I__789 (
            .O(N__4347),
            .I(D_UU_040_in_3));
    IoInMux I__788 (
            .O(N__4344),
            .I(N__4341));
    LocalMux I__787 (
            .O(N__4341),
            .I(N__4338));
    Span12Mux_s1_v I__786 (
            .O(N__4338),
            .I(N__4335));
    Span12Mux_h I__785 (
            .O(N__4335),
            .I(N__4332));
    Odrv12 I__784 (
            .O(N__4332),
            .I(un1_D_UU_040_3));
    CascadeMux I__783 (
            .O(N__4329),
            .I(N__4326));
    InMux I__782 (
            .O(N__4326),
            .I(N__4323));
    LocalMux I__781 (
            .O(N__4323),
            .I(N__4319));
    InMux I__780 (
            .O(N__4322),
            .I(N__4316));
    Span4Mux_v I__779 (
            .O(N__4319),
            .I(N__4313));
    LocalMux I__778 (
            .O(N__4316),
            .I(N__4310));
    Span4Mux_h I__777 (
            .O(N__4313),
            .I(N__4304));
    Span4Mux_v I__776 (
            .O(N__4310),
            .I(N__4304));
    InMux I__775 (
            .O(N__4309),
            .I(N__4301));
    Span4Mux_v I__774 (
            .O(N__4304),
            .I(N__4298));
    LocalMux I__773 (
            .O(N__4301),
            .I(N__4295));
    Span4Mux_v I__772 (
            .O(N__4298),
            .I(N__4290));
    Span4Mux_h I__771 (
            .O(N__4295),
            .I(N__4290));
    Span4Mux_v I__770 (
            .O(N__4290),
            .I(N__4287));
    Span4Mux_h I__769 (
            .O(N__4287),
            .I(N__4284));
    Span4Mux_h I__768 (
            .O(N__4284),
            .I(N__4281));
    Odrv4 I__767 (
            .O(N__4281),
            .I(D_UU_AMIGA_in_5));
    InMux I__766 (
            .O(N__4278),
            .I(N__4274));
    InMux I__765 (
            .O(N__4277),
            .I(N__4271));
    LocalMux I__764 (
            .O(N__4274),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_1 ));
    LocalMux I__763 (
            .O(N__4271),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_1 ));
    InMux I__762 (
            .O(N__4266),
            .I(N__4260));
    InMux I__761 (
            .O(N__4265),
            .I(N__4260));
    LocalMux I__760 (
            .O(N__4260),
            .I(N__4257));
    Span4Mux_v I__759 (
            .O(N__4257),
            .I(N__4254));
    Sp12to4 I__758 (
            .O(N__4254),
            .I(N__4251));
    Span12Mux_h I__757 (
            .O(N__4251),
            .I(N__4248));
    Span12Mux_v I__756 (
            .O(N__4248),
            .I(N__4245));
    Odrv12 I__755 (
            .O(N__4245),
            .I(SIZ_c_0));
    CascadeMux I__754 (
            .O(N__4242),
            .I(N__4238));
    InMux I__753 (
            .O(N__4241),
            .I(N__4233));
    InMux I__752 (
            .O(N__4238),
            .I(N__4233));
    LocalMux I__751 (
            .O(N__4233),
            .I(N__4230));
    Span4Mux_v I__750 (
            .O(N__4230),
            .I(N__4227));
    Sp12to4 I__749 (
            .O(N__4227),
            .I(N__4224));
    Span12Mux_h I__748 (
            .O(N__4224),
            .I(N__4221));
    Span12Mux_v I__747 (
            .O(N__4221),
            .I(N__4218));
    Odrv12 I__746 (
            .O(N__4218),
            .I(SIZ_c_1));
    CascadeMux I__745 (
            .O(N__4215),
            .I(N__4210));
    InMux I__744 (
            .O(N__4214),
            .I(N__4205));
    InMux I__743 (
            .O(N__4213),
            .I(N__4205));
    InMux I__742 (
            .O(N__4210),
            .I(N__4202));
    LocalMux I__741 (
            .O(N__4205),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ));
    LocalMux I__740 (
            .O(N__4202),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ));
    CascadeMux I__739 (
            .O(N__4197),
            .I(N__4194));
    InMux I__738 (
            .O(N__4194),
            .I(N__4187));
    InMux I__737 (
            .O(N__4193),
            .I(N__4187));
    InMux I__736 (
            .O(N__4192),
            .I(N__4184));
    LocalMux I__735 (
            .O(N__4187),
            .I(\U111_CYCLE_SM.LW_TRANSZ0 ));
    LocalMux I__734 (
            .O(N__4184),
            .I(\U111_CYCLE_SM.LW_TRANSZ0 ));
    InMux I__733 (
            .O(N__4179),
            .I(N__4170));
    InMux I__732 (
            .O(N__4178),
            .I(N__4170));
    InMux I__731 (
            .O(N__4177),
            .I(N__4167));
    InMux I__730 (
            .O(N__4176),
            .I(N__4162));
    InMux I__729 (
            .O(N__4175),
            .I(N__4162));
    LocalMux I__728 (
            .O(N__4170),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__727 (
            .O(N__4167),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__726 (
            .O(N__4162),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    InMux I__725 (
            .O(N__4155),
            .I(N__4151));
    InMux I__724 (
            .O(N__4154),
            .I(N__4148));
    LocalMux I__723 (
            .O(N__4151),
            .I(N__4143));
    LocalMux I__722 (
            .O(N__4148),
            .I(N__4143));
    Span4Mux_v I__721 (
            .O(N__4143),
            .I(N__4139));
    InMux I__720 (
            .O(N__4142),
            .I(N__4136));
    Sp12to4 I__719 (
            .O(N__4139),
            .I(N__4131));
    LocalMux I__718 (
            .O(N__4136),
            .I(N__4131));
    Span12Mux_h I__717 (
            .O(N__4131),
            .I(N__4128));
    Span12Mux_v I__716 (
            .O(N__4128),
            .I(N__4125));
    Odrv12 I__715 (
            .O(N__4125),
            .I(PORTSIZE_c));
    InMux I__714 (
            .O(N__4122),
            .I(N__4119));
    LocalMux I__713 (
            .O(N__4119),
            .I(\U111_CYCLE_SM.N_179 ));
    CascadeMux I__712 (
            .O(N__4116),
            .I(\U111_CYCLE_SM.N_179_cascade_ ));
    CascadeMux I__711 (
            .O(N__4113),
            .I(\U111_CYCLE_SM.N_101_cascade_ ));
    CascadeMux I__710 (
            .O(N__4110),
            .I(N__4107));
    InMux I__709 (
            .O(N__4107),
            .I(N__4100));
    InMux I__708 (
            .O(N__4106),
            .I(N__4100));
    CascadeMux I__707 (
            .O(N__4105),
            .I(N__4097));
    LocalMux I__706 (
            .O(N__4100),
            .I(N__4094));
    InMux I__705 (
            .O(N__4097),
            .I(N__4091));
    Odrv12 I__704 (
            .O(N__4094),
            .I(\U111_CYCLE_SM.N_98 ));
    LocalMux I__703 (
            .O(N__4091),
            .I(\U111_CYCLE_SM.N_98 ));
    InMux I__702 (
            .O(N__4086),
            .I(N__4083));
    LocalMux I__701 (
            .O(N__4083),
            .I(\U111_CYCLE_SM.N_10 ));
    InMux I__700 (
            .O(N__4080),
            .I(N__4077));
    LocalMux I__699 (
            .O(N__4077),
            .I(\U111_CYCLE_SM.N_101 ));
    CascadeMux I__698 (
            .O(N__4074),
            .I(\U111_CYCLE_SM.N_12_i_1_cascade_ ));
    InMux I__697 (
            .O(N__4071),
            .I(N__4068));
    LocalMux I__696 (
            .O(N__4068),
            .I(\U111_CYCLE_SM.N_55 ));
    InMux I__695 (
            .O(N__4065),
            .I(N__4061));
    InMux I__694 (
            .O(N__4064),
            .I(N__4058));
    LocalMux I__693 (
            .O(N__4061),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    LocalMux I__692 (
            .O(N__4058),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    InMux I__691 (
            .O(N__4053),
            .I(N__4050));
    LocalMux I__690 (
            .O(N__4050),
            .I(N__4047));
    Span4Mux_v I__689 (
            .O(N__4047),
            .I(N__4044));
    Sp12to4 I__688 (
            .O(N__4044),
            .I(N__4041));
    Span12Mux_h I__687 (
            .O(N__4041),
            .I(N__4038));
    Odrv12 I__686 (
            .O(N__4038),
            .I(D_LM_AMIGA_in_7));
    IoInMux I__685 (
            .O(N__4035),
            .I(N__4032));
    LocalMux I__684 (
            .O(N__4032),
            .I(N__4029));
    IoSpan4Mux I__683 (
            .O(N__4029),
            .I(N__4026));
    Span4Mux_s3_h I__682 (
            .O(N__4026),
            .I(N__4023));
    Span4Mux_h I__681 (
            .O(N__4023),
            .I(N__4020));
    Sp12to4 I__680 (
            .O(N__4020),
            .I(N__4017));
    Odrv12 I__679 (
            .O(N__4017),
            .I(N_106));
    InMux I__678 (
            .O(N__4014),
            .I(N__4011));
    LocalMux I__677 (
            .O(N__4011),
            .I(N__4008));
    Span12Mux_v I__676 (
            .O(N__4008),
            .I(N__4005));
    Span12Mux_h I__675 (
            .O(N__4005),
            .I(N__4002));
    Odrv12 I__674 (
            .O(N__4002),
            .I(D_LM_AMIGA_in_6));
    IoInMux I__673 (
            .O(N__3999),
            .I(N__3996));
    LocalMux I__672 (
            .O(N__3996),
            .I(N__3993));
    IoSpan4Mux I__671 (
            .O(N__3993),
            .I(N__3990));
    Sp12to4 I__670 (
            .O(N__3990),
            .I(N__3987));
    Span12Mux_s9_h I__669 (
            .O(N__3987),
            .I(N__3984));
    Odrv12 I__668 (
            .O(N__3984),
            .I(N_107));
    InMux I__667 (
            .O(N__3981),
            .I(N__3978));
    LocalMux I__666 (
            .O(N__3978),
            .I(N__3975));
    Span12Mux_v I__665 (
            .O(N__3975),
            .I(N__3972));
    Span12Mux_h I__664 (
            .O(N__3972),
            .I(N__3969));
    Odrv12 I__663 (
            .O(N__3969),
            .I(D_UM_040_in_3));
    InMux I__662 (
            .O(N__3966),
            .I(N__3962));
    IoInMux I__661 (
            .O(N__3965),
            .I(N__3959));
    LocalMux I__660 (
            .O(N__3962),
            .I(N__3956));
    LocalMux I__659 (
            .O(N__3959),
            .I(N__3953));
    Span4Mux_v I__658 (
            .O(N__3956),
            .I(N__3950));
    Span4Mux_s3_h I__657 (
            .O(N__3953),
            .I(N__3947));
    Sp12to4 I__656 (
            .O(N__3950),
            .I(N__3944));
    Sp12to4 I__655 (
            .O(N__3947),
            .I(N__3941));
    Span12Mux_h I__654 (
            .O(N__3944),
            .I(N__3938));
    Span12Mux_v I__653 (
            .O(N__3941),
            .I(N__3935));
    Span12Mux_v I__652 (
            .O(N__3938),
            .I(N__3932));
    Span12Mux_h I__651 (
            .O(N__3935),
            .I(N__3929));
    Span12Mux_v I__650 (
            .O(N__3932),
            .I(N__3924));
    Span12Mux_h I__649 (
            .O(N__3929),
            .I(N__3924));
    Odrv12 I__648 (
            .O(N__3924),
            .I(D_LL_040_in_3));
    IoInMux I__647 (
            .O(N__3921),
            .I(N__3918));
    LocalMux I__646 (
            .O(N__3918),
            .I(N__3915));
    IoSpan4Mux I__645 (
            .O(N__3915),
            .I(N__3912));
    Span4Mux_s2_h I__644 (
            .O(N__3912),
            .I(N__3909));
    Sp12to4 I__643 (
            .O(N__3909),
            .I(N__3906));
    Odrv12 I__642 (
            .O(N__3906),
            .I(un1_D_UM_040_3));
    InMux I__641 (
            .O(N__3903),
            .I(N__3900));
    LocalMux I__640 (
            .O(N__3900),
            .I(N__3897));
    Span4Mux_v I__639 (
            .O(N__3897),
            .I(N__3894));
    Span4Mux_h I__638 (
            .O(N__3894),
            .I(N__3891));
    Sp12to4 I__637 (
            .O(N__3891),
            .I(N__3888));
    Odrv12 I__636 (
            .O(N__3888),
            .I(D_LL_AMIGA_in_3));
    IoInMux I__635 (
            .O(N__3885),
            .I(N__3882));
    LocalMux I__634 (
            .O(N__3882),
            .I(N__3879));
    Span4Mux_s2_h I__633 (
            .O(N__3879),
            .I(N__3876));
    Span4Mux_v I__632 (
            .O(N__3876),
            .I(N__3873));
    Span4Mux_h I__631 (
            .O(N__3873),
            .I(N__3870));
    Sp12to4 I__630 (
            .O(N__3870),
            .I(N__3867));
    Span12Mux_h I__629 (
            .O(N__3867),
            .I(N__3864));
    Odrv12 I__628 (
            .O(N__3864),
            .I(un2_D_LL_AMIGA_3));
    IoInMux I__627 (
            .O(N__3861),
            .I(N__3858));
    LocalMux I__626 (
            .O(N__3858),
            .I(N__3855));
    Odrv12 I__625 (
            .O(N__3855),
            .I(LBENn_c_i));
    InMux I__624 (
            .O(N__3852),
            .I(N__3849));
    LocalMux I__623 (
            .O(N__3849),
            .I(N__3846));
    Span4Mux_v I__622 (
            .O(N__3846),
            .I(N__3843));
    Sp12to4 I__621 (
            .O(N__3843),
            .I(N__3840));
    Span12Mux_h I__620 (
            .O(N__3840),
            .I(N__3837));
    Odrv12 I__619 (
            .O(N__3837),
            .I(D_LM_AMIGA_in_0));
    IoInMux I__618 (
            .O(N__3834),
            .I(N__3831));
    LocalMux I__617 (
            .O(N__3831),
            .I(N__3828));
    IoSpan4Mux I__616 (
            .O(N__3828),
            .I(N__3825));
    Span4Mux_s3_h I__615 (
            .O(N__3825),
            .I(N__3822));
    Sp12to4 I__614 (
            .O(N__3822),
            .I(N__3819));
    Span12Mux_h I__613 (
            .O(N__3819),
            .I(N__3816));
    Odrv12 I__612 (
            .O(N__3816),
            .I(un2_D_LM_AMIGA_0));
    InMux I__611 (
            .O(N__3813),
            .I(N__3807));
    InMux I__610 (
            .O(N__3812),
            .I(N__3807));
    LocalMux I__609 (
            .O(N__3807),
            .I(N__3804));
    Span4Mux_h I__608 (
            .O(N__3804),
            .I(N__3801));
    Span4Mux_v I__607 (
            .O(N__3801),
            .I(N__3798));
    Span4Mux_h I__606 (
            .O(N__3798),
            .I(N__3794));
    InMux I__605 (
            .O(N__3797),
            .I(N__3791));
    Odrv4 I__604 (
            .O(N__3794),
            .I(\U111_CYCLE_SM.A2_ENZ0 ));
    LocalMux I__603 (
            .O(N__3791),
            .I(\U111_CYCLE_SM.A2_ENZ0 ));
    InMux I__602 (
            .O(N__3786),
            .I(N__3783));
    LocalMux I__601 (
            .O(N__3783),
            .I(N__3780));
    Span4Mux_v I__600 (
            .O(N__3780),
            .I(N__3777));
    Sp12to4 I__599 (
            .O(N__3777),
            .I(N__3774));
    Span12Mux_h I__598 (
            .O(N__3774),
            .I(N__3771));
    Odrv12 I__597 (
            .O(N__3771),
            .I(D_LL_AMIGA_in_2));
    IoInMux I__596 (
            .O(N__3768),
            .I(N__3765));
    LocalMux I__595 (
            .O(N__3765),
            .I(N__3762));
    Span12Mux_s7_h I__594 (
            .O(N__3762),
            .I(N__3759));
    Span12Mux_h I__593 (
            .O(N__3759),
            .I(N__3756));
    Odrv12 I__592 (
            .O(N__3756),
            .I(un2_D_LL_AMIGA_2));
    IoInMux I__591 (
            .O(N__3753),
            .I(N__3750));
    LocalMux I__590 (
            .O(N__3750),
            .I(N__3746));
    InMux I__589 (
            .O(N__3749),
            .I(N__3743));
    IoSpan4Mux I__588 (
            .O(N__3746),
            .I(N__3740));
    LocalMux I__587 (
            .O(N__3743),
            .I(N__3737));
    Span4Mux_s2_h I__586 (
            .O(N__3740),
            .I(N__3734));
    Span4Mux_v I__585 (
            .O(N__3737),
            .I(N__3731));
    Sp12to4 I__584 (
            .O(N__3734),
            .I(N__3728));
    Sp12to4 I__583 (
            .O(N__3731),
            .I(N__3725));
    Span12Mux_h I__582 (
            .O(N__3728),
            .I(N__3720));
    Span12Mux_v I__581 (
            .O(N__3725),
            .I(N__3720));
    Span12Mux_h I__580 (
            .O(N__3720),
            .I(N__3717));
    Odrv12 I__579 (
            .O(N__3717),
            .I(D_LL_040_in_0));
    InMux I__578 (
            .O(N__3714),
            .I(N__3711));
    LocalMux I__577 (
            .O(N__3711),
            .I(N__3708));
    Span4Mux_v I__576 (
            .O(N__3708),
            .I(N__3705));
    Sp12to4 I__575 (
            .O(N__3705),
            .I(N__3702));
    Span12Mux_h I__574 (
            .O(N__3702),
            .I(N__3699));
    Span12Mux_h I__573 (
            .O(N__3699),
            .I(N__3696));
    Odrv12 I__572 (
            .O(N__3696),
            .I(D_UM_040_in_0));
    IoInMux I__571 (
            .O(N__3693),
            .I(N__3690));
    LocalMux I__570 (
            .O(N__3690),
            .I(N__3687));
    IoSpan4Mux I__569 (
            .O(N__3687),
            .I(N__3684));
    Sp12to4 I__568 (
            .O(N__3684),
            .I(N__3681));
    Span12Mux_h I__567 (
            .O(N__3681),
            .I(N__3678));
    Odrv12 I__566 (
            .O(N__3678),
            .I(un1_D_UM_040_0));
    InMux I__565 (
            .O(N__3675),
            .I(N__3672));
    LocalMux I__564 (
            .O(N__3672),
            .I(N__3669));
    Span12Mux_h I__563 (
            .O(N__3669),
            .I(N__3666));
    Odrv12 I__562 (
            .O(N__3666),
            .I(D_LM_AMIGA_in_1));
    IoInMux I__561 (
            .O(N__3663),
            .I(N__3660));
    LocalMux I__560 (
            .O(N__3660),
            .I(N__3657));
    IoSpan4Mux I__559 (
            .O(N__3657),
            .I(N__3654));
    Sp12to4 I__558 (
            .O(N__3654),
            .I(N__3651));
    Span12Mux_s7_h I__557 (
            .O(N__3651),
            .I(N__3648));
    Span12Mux_h I__556 (
            .O(N__3648),
            .I(N__3645));
    Odrv12 I__555 (
            .O(N__3645),
            .I(N_112));
    IoInMux I__554 (
            .O(N__3642),
            .I(N__3639));
    LocalMux I__553 (
            .O(N__3639),
            .I(N__3636));
    Span4Mux_s2_v I__552 (
            .O(N__3636),
            .I(N__3633));
    Span4Mux_h I__551 (
            .O(N__3633),
            .I(N__3630));
    Span4Mux_v I__550 (
            .O(N__3630),
            .I(N__3627));
    Odrv4 I__549 (
            .O(N__3627),
            .I(N_96));
    IoInMux I__548 (
            .O(N__3624),
            .I(N__3621));
    LocalMux I__547 (
            .O(N__3621),
            .I(N__3618));
    Span4Mux_s2_v I__546 (
            .O(N__3618),
            .I(N__3615));
    Span4Mux_h I__545 (
            .O(N__3615),
            .I(N__3612));
    Span4Mux_v I__544 (
            .O(N__3612),
            .I(N__3609));
    Odrv4 I__543 (
            .O(N__3609),
            .I(N_94_i));
    InMux I__542 (
            .O(N__3606),
            .I(N__3601));
    InMux I__541 (
            .O(N__3605),
            .I(N__3596));
    InMux I__540 (
            .O(N__3604),
            .I(N__3596));
    LocalMux I__539 (
            .O(N__3601),
            .I(N__3591));
    LocalMux I__538 (
            .O(N__3596),
            .I(N__3591));
    Span4Mux_h I__537 (
            .O(N__3591),
            .I(N__3588));
    Span4Mux_v I__536 (
            .O(N__3588),
            .I(N__3585));
    Odrv4 I__535 (
            .O(N__3585),
            .I(BBn_c));
    IoInMux I__534 (
            .O(N__3582),
            .I(N__3579));
    LocalMux I__533 (
            .O(N__3579),
            .I(N__3576));
    IoSpan4Mux I__532 (
            .O(N__3576),
            .I(N__3573));
    Span4Mux_s2_v I__531 (
            .O(N__3573),
            .I(N__3570));
    Span4Mux_v I__530 (
            .O(N__3570),
            .I(N__3567));
    Odrv4 I__529 (
            .O(N__3567),
            .I(BUFDIR_c));
    IoInMux I__528 (
            .O(N__3564),
            .I(N__3560));
    IoInMux I__527 (
            .O(N__3563),
            .I(N__3557));
    LocalMux I__526 (
            .O(N__3560),
            .I(N__3553));
    LocalMux I__525 (
            .O(N__3557),
            .I(N__3549));
    IoInMux I__524 (
            .O(N__3556),
            .I(N__3546));
    IoSpan4Mux I__523 (
            .O(N__3553),
            .I(N__3543));
    IoInMux I__522 (
            .O(N__3552),
            .I(N__3540));
    Span4Mux_s2_h I__521 (
            .O(N__3549),
            .I(N__3537));
    LocalMux I__520 (
            .O(N__3546),
            .I(N__3534));
    IoSpan4Mux I__519 (
            .O(N__3543),
            .I(N__3529));
    LocalMux I__518 (
            .O(N__3540),
            .I(N__3529));
    Span4Mux_h I__517 (
            .O(N__3537),
            .I(N__3526));
    Span4Mux_s1_h I__516 (
            .O(N__3534),
            .I(N__3523));
    IoSpan4Mux I__515 (
            .O(N__3529),
            .I(N__3520));
    Span4Mux_h I__514 (
            .O(N__3526),
            .I(N__3517));
    Span4Mux_h I__513 (
            .O(N__3523),
            .I(N__3514));
    Span4Mux_s3_v I__512 (
            .O(N__3520),
            .I(N__3511));
    Span4Mux_h I__511 (
            .O(N__3517),
            .I(N__3508));
    Span4Mux_h I__510 (
            .O(N__3514),
            .I(N__3505));
    Sp12to4 I__509 (
            .O(N__3511),
            .I(N__3502));
    Span4Mux_h I__508 (
            .O(N__3508),
            .I(N__3497));
    Span4Mux_h I__507 (
            .O(N__3505),
            .I(N__3497));
    Odrv12 I__506 (
            .O(N__3502),
            .I(GB_BUFFER_CLK40_THRU_CO));
    Odrv4 I__505 (
            .O(N__3497),
            .I(GB_BUFFER_CLK40_THRU_CO));
    CascadeMux I__504 (
            .O(N__3492),
            .I(N__3489));
    InMux I__503 (
            .O(N__3489),
            .I(N__3486));
    LocalMux I__502 (
            .O(N__3486),
            .I(N__3483));
    Span4Mux_v I__501 (
            .O(N__3483),
            .I(N__3480));
    Odrv4 I__500 (
            .O(N__3480),
            .I(\U111_CYCLE_SM.N_141 ));
    InMux I__499 (
            .O(N__3477),
            .I(N__3474));
    LocalMux I__498 (
            .O(N__3474),
            .I(N__3471));
    Span4Mux_v I__497 (
            .O(N__3471),
            .I(N__3468));
    Span4Mux_v I__496 (
            .O(N__3468),
            .I(N__3464));
    InMux I__495 (
            .O(N__3467),
            .I(N__3461));
    Sp12to4 I__494 (
            .O(N__3464),
            .I(N__3456));
    LocalMux I__493 (
            .O(N__3461),
            .I(N__3456));
    Span12Mux_h I__492 (
            .O(N__3456),
            .I(N__3453));
    Odrv12 I__491 (
            .O(N__3453),
            .I(A_040_c_1));
    InMux I__490 (
            .O(N__3450),
            .I(N__3447));
    LocalMux I__489 (
            .O(N__3447),
            .I(N__3444));
    Span12Mux_v I__488 (
            .O(N__3444),
            .I(N__3441));
    Odrv12 I__487 (
            .O(N__3441),
            .I(D_LM_AMIGA_in_5));
    IoInMux I__486 (
            .O(N__3438),
            .I(N__3435));
    LocalMux I__485 (
            .O(N__3435),
            .I(N__3432));
    Span12Mux_s8_h I__484 (
            .O(N__3432),
            .I(N__3429));
    Span12Mux_h I__483 (
            .O(N__3429),
            .I(N__3426));
    Odrv12 I__482 (
            .O(N__3426),
            .I(N_108));
    InMux I__481 (
            .O(N__3423),
            .I(N__3420));
    LocalMux I__480 (
            .O(N__3420),
            .I(N__3417));
    Span12Mux_h I__479 (
            .O(N__3417),
            .I(N__3414));
    Odrv12 I__478 (
            .O(N__3414),
            .I(D_LM_AMIGA_in_3));
    IoInMux I__477 (
            .O(N__3411),
            .I(N__3408));
    LocalMux I__476 (
            .O(N__3408),
            .I(N__3405));
    IoSpan4Mux I__475 (
            .O(N__3405),
            .I(N__3402));
    Span4Mux_s1_h I__474 (
            .O(N__3402),
            .I(N__3399));
    Span4Mux_v I__473 (
            .O(N__3399),
            .I(N__3396));
    Sp12to4 I__472 (
            .O(N__3396),
            .I(N__3393));
    Span12Mux_s10_h I__471 (
            .O(N__3393),
            .I(N__3390));
    Odrv12 I__470 (
            .O(N__3390),
            .I(N_110));
    InMux I__469 (
            .O(N__3387),
            .I(N__3384));
    LocalMux I__468 (
            .O(N__3384),
            .I(N__3381));
    Span12Mux_h I__467 (
            .O(N__3381),
            .I(N__3378));
    Odrv12 I__466 (
            .O(N__3378),
            .I(D_LM_AMIGA_in_2));
    IoInMux I__465 (
            .O(N__3375),
            .I(N__3372));
    LocalMux I__464 (
            .O(N__3372),
            .I(N__3369));
    Span12Mux_s3_h I__463 (
            .O(N__3369),
            .I(N__3366));
    Span12Mux_h I__462 (
            .O(N__3366),
            .I(N__3363));
    Span12Mux_v I__461 (
            .O(N__3363),
            .I(N__3360));
    Odrv12 I__460 (
            .O(N__3360),
            .I(N_111));
    InMux I__459 (
            .O(N__3357),
            .I(N__3354));
    LocalMux I__458 (
            .O(N__3354),
            .I(N__3351));
    Span4Mux_v I__457 (
            .O(N__3351),
            .I(N__3348));
    Sp12to4 I__456 (
            .O(N__3348),
            .I(N__3345));
    Span12Mux_h I__455 (
            .O(N__3345),
            .I(N__3342));
    Odrv12 I__454 (
            .O(N__3342),
            .I(D_UM_040_in_6));
    IoInMux I__453 (
            .O(N__3339),
            .I(N__3336));
    LocalMux I__452 (
            .O(N__3336),
            .I(N__3333));
    IoSpan4Mux I__451 (
            .O(N__3333),
            .I(N__3329));
    InMux I__450 (
            .O(N__3332),
            .I(N__3326));
    IoSpan4Mux I__449 (
            .O(N__3329),
            .I(N__3323));
    LocalMux I__448 (
            .O(N__3326),
            .I(N__3320));
    Span4Mux_s2_h I__447 (
            .O(N__3323),
            .I(N__3317));
    Span4Mux_v I__446 (
            .O(N__3320),
            .I(N__3314));
    Sp12to4 I__445 (
            .O(N__3317),
            .I(N__3311));
    Sp12to4 I__444 (
            .O(N__3314),
            .I(N__3308));
    Span12Mux_h I__443 (
            .O(N__3311),
            .I(N__3305));
    Span12Mux_h I__442 (
            .O(N__3308),
            .I(N__3302));
    Span12Mux_h I__441 (
            .O(N__3305),
            .I(N__3297));
    Span12Mux_v I__440 (
            .O(N__3302),
            .I(N__3297));
    Odrv12 I__439 (
            .O(N__3297),
            .I(D_LL_040_in_6));
    IoInMux I__438 (
            .O(N__3294),
            .I(N__3291));
    LocalMux I__437 (
            .O(N__3291),
            .I(N__3288));
    Span12Mux_s9_h I__436 (
            .O(N__3288),
            .I(N__3285));
    Span12Mux_v I__435 (
            .O(N__3285),
            .I(N__3282));
    Odrv12 I__434 (
            .O(N__3282),
            .I(un1_D_UM_040_6));
    InMux I__433 (
            .O(N__3279),
            .I(N__3276));
    LocalMux I__432 (
            .O(N__3276),
            .I(N__3273));
    Span4Mux_v I__431 (
            .O(N__3273),
            .I(N__3270));
    Span4Mux_h I__430 (
            .O(N__3270),
            .I(N__3267));
    Sp12to4 I__429 (
            .O(N__3267),
            .I(N__3264));
    Span12Mux_h I__428 (
            .O(N__3264),
            .I(N__3261));
    Odrv12 I__427 (
            .O(N__3261),
            .I(D_UU_040_in_0));
    IoInMux I__426 (
            .O(N__3258),
            .I(N__3254));
    InMux I__425 (
            .O(N__3257),
            .I(N__3251));
    LocalMux I__424 (
            .O(N__3254),
            .I(N__3248));
    LocalMux I__423 (
            .O(N__3251),
            .I(N__3245));
    IoSpan4Mux I__422 (
            .O(N__3248),
            .I(N__3242));
    Span4Mux_v I__421 (
            .O(N__3245),
            .I(N__3239));
    Span4Mux_s2_h I__420 (
            .O(N__3242),
            .I(N__3236));
    Sp12to4 I__419 (
            .O(N__3239),
            .I(N__3233));
    Span4Mux_v I__418 (
            .O(N__3236),
            .I(N__3230));
    Span12Mux_h I__417 (
            .O(N__3233),
            .I(N__3227));
    Sp12to4 I__416 (
            .O(N__3230),
            .I(N__3224));
    Span12Mux_v I__415 (
            .O(N__3227),
            .I(N__3221));
    Span12Mux_s9_h I__414 (
            .O(N__3224),
            .I(N__3218));
    Span12Mux_v I__413 (
            .O(N__3221),
            .I(N__3213));
    Span12Mux_h I__412 (
            .O(N__3218),
            .I(N__3213));
    Odrv12 I__411 (
            .O(N__3213),
            .I(D_LM_040_in_0));
    IoInMux I__410 (
            .O(N__3210),
            .I(N__3207));
    LocalMux I__409 (
            .O(N__3207),
            .I(N__3204));
    IoSpan4Mux I__408 (
            .O(N__3204),
            .I(N__3201));
    Span4Mux_s2_v I__407 (
            .O(N__3201),
            .I(N__3198));
    Span4Mux_v I__406 (
            .O(N__3198),
            .I(N__3195));
    Odrv4 I__405 (
            .O(N__3195),
            .I(un1_D_UU_040_0));
    InMux I__404 (
            .O(N__3192),
            .I(N__3189));
    LocalMux I__403 (
            .O(N__3189),
            .I(N__3186));
    Span4Mux_v I__402 (
            .O(N__3186),
            .I(N__3183));
    Span4Mux_h I__401 (
            .O(N__3183),
            .I(N__3180));
    Sp12to4 I__400 (
            .O(N__3180),
            .I(N__3177));
    Span12Mux_h I__399 (
            .O(N__3177),
            .I(N__3174));
    Odrv12 I__398 (
            .O(N__3174),
            .I(D_UU_040_in_6));
    IoInMux I__397 (
            .O(N__3171),
            .I(N__3168));
    LocalMux I__396 (
            .O(N__3168),
            .I(N__3164));
    InMux I__395 (
            .O(N__3167),
            .I(N__3161));
    Span4Mux_s2_h I__394 (
            .O(N__3164),
            .I(N__3158));
    LocalMux I__393 (
            .O(N__3161),
            .I(N__3155));
    Span4Mux_v I__392 (
            .O(N__3158),
            .I(N__3152));
    Span4Mux_v I__391 (
            .O(N__3155),
            .I(N__3149));
    Sp12to4 I__390 (
            .O(N__3152),
            .I(N__3146));
    Span4Mux_v I__389 (
            .O(N__3149),
            .I(N__3143));
    Span12Mux_h I__388 (
            .O(N__3146),
            .I(N__3138));
    Sp12to4 I__387 (
            .O(N__3143),
            .I(N__3138));
    Span12Mux_h I__386 (
            .O(N__3138),
            .I(N__3135));
    Odrv12 I__385 (
            .O(N__3135),
            .I(D_LM_040_in_6));
    IoInMux I__384 (
            .O(N__3132),
            .I(N__3129));
    LocalMux I__383 (
            .O(N__3129),
            .I(N__3126));
    Span4Mux_s3_v I__382 (
            .O(N__3126),
            .I(N__3123));
    Span4Mux_h I__381 (
            .O(N__3123),
            .I(N__3120));
    Span4Mux_h I__380 (
            .O(N__3120),
            .I(N__3117));
    Odrv4 I__379 (
            .O(N__3117),
            .I(un1_D_UU_040_6));
    InMux I__378 (
            .O(N__3114),
            .I(N__3111));
    LocalMux I__377 (
            .O(N__3111),
            .I(N__3108));
    Span4Mux_v I__376 (
            .O(N__3108),
            .I(N__3105));
    Sp12to4 I__375 (
            .O(N__3105),
            .I(N__3102));
    Odrv12 I__374 (
            .O(N__3102),
            .I(D_LL_AMIGA_in_4));
    IoInMux I__373 (
            .O(N__3099),
            .I(N__3096));
    LocalMux I__372 (
            .O(N__3096),
            .I(N__3093));
    Span4Mux_s2_h I__371 (
            .O(N__3093),
            .I(N__3090));
    Sp12to4 I__370 (
            .O(N__3090),
            .I(N__3087));
    Span12Mux_s8_v I__369 (
            .O(N__3087),
            .I(N__3084));
    Span12Mux_h I__368 (
            .O(N__3084),
            .I(N__3081));
    Odrv12 I__367 (
            .O(N__3081),
            .I(un2_D_LL_AMIGA_4));
    IoInMux I__366 (
            .O(N__3078),
            .I(N__3075));
    LocalMux I__365 (
            .O(N__3075),
            .I(N__3072));
    Odrv12 I__364 (
            .O(N__3072),
            .I(U111_CYCLE_SM_A_AMIGA_0_i_1));
    InMux I__363 (
            .O(N__3069),
            .I(N__3066));
    LocalMux I__362 (
            .O(N__3066),
            .I(N__3063));
    Span4Mux_h I__361 (
            .O(N__3063),
            .I(N__3060));
    Span4Mux_v I__360 (
            .O(N__3060),
            .I(N__3057));
    Odrv4 I__359 (
            .O(N__3057),
            .I(A_040_c_0));
    IoInMux I__358 (
            .O(N__3054),
            .I(N__3051));
    LocalMux I__357 (
            .O(N__3051),
            .I(N__3048));
    Span12Mux_s6_v I__356 (
            .O(N__3048),
            .I(N__3045));
    Odrv12 I__355 (
            .O(N__3045),
            .I(A_AMIGA_c_0));
    InMux I__354 (
            .O(N__3042),
            .I(N__3039));
    LocalMux I__353 (
            .O(N__3039),
            .I(N__3036));
    Span12Mux_h I__352 (
            .O(N__3036),
            .I(N__3033));
    Span12Mux_h I__351 (
            .O(N__3033),
            .I(N__3030));
    Odrv12 I__350 (
            .O(N__3030),
            .I(D_UM_040_in_2));
    IoInMux I__349 (
            .O(N__3027),
            .I(N__3023));
    InMux I__348 (
            .O(N__3026),
            .I(N__3020));
    LocalMux I__347 (
            .O(N__3023),
            .I(N__3017));
    LocalMux I__346 (
            .O(N__3020),
            .I(N__3014));
    IoSpan4Mux I__345 (
            .O(N__3017),
            .I(N__3011));
    Span4Mux_v I__344 (
            .O(N__3014),
            .I(N__3008));
    Span4Mux_s2_h I__343 (
            .O(N__3011),
            .I(N__3005));
    Sp12to4 I__342 (
            .O(N__3008),
            .I(N__3002));
    Sp12to4 I__341 (
            .O(N__3005),
            .I(N__2999));
    Span12Mux_h I__340 (
            .O(N__3002),
            .I(N__2996));
    Span12Mux_h I__339 (
            .O(N__2999),
            .I(N__2993));
    Span12Mux_v I__338 (
            .O(N__2996),
            .I(N__2990));
    Span12Mux_h I__337 (
            .O(N__2993),
            .I(N__2987));
    Odrv12 I__336 (
            .O(N__2990),
            .I(D_LL_040_in_2));
    Odrv12 I__335 (
            .O(N__2987),
            .I(D_LL_040_in_2));
    IoInMux I__334 (
            .O(N__2982),
            .I(N__2979));
    LocalMux I__333 (
            .O(N__2979),
            .I(N__2976));
    Span4Mux_s3_h I__332 (
            .O(N__2976),
            .I(N__2973));
    Span4Mux_h I__331 (
            .O(N__2973),
            .I(N__2970));
    Span4Mux_v I__330 (
            .O(N__2970),
            .I(N__2967));
    Odrv4 I__329 (
            .O(N__2967),
            .I(un1_D_UM_040_2));
    InMux I__328 (
            .O(N__2964),
            .I(N__2961));
    LocalMux I__327 (
            .O(N__2961),
            .I(N__2958));
    Span4Mux_h I__326 (
            .O(N__2958),
            .I(N__2955));
    Span4Mux_v I__325 (
            .O(N__2955),
            .I(N__2952));
    Span4Mux_h I__324 (
            .O(N__2952),
            .I(N__2949));
    Span4Mux_h I__323 (
            .O(N__2949),
            .I(N__2946));
    Span4Mux_h I__322 (
            .O(N__2946),
            .I(N__2943));
    Odrv4 I__321 (
            .O(N__2943),
            .I(D_UU_040_in_4));
    IoInMux I__320 (
            .O(N__2940),
            .I(N__2937));
    LocalMux I__319 (
            .O(N__2937),
            .I(N__2934));
    Span4Mux_s1_h I__318 (
            .O(N__2934),
            .I(N__2931));
    Span4Mux_h I__317 (
            .O(N__2931),
            .I(N__2927));
    InMux I__316 (
            .O(N__2930),
            .I(N__2924));
    Sp12to4 I__315 (
            .O(N__2927),
            .I(N__2921));
    LocalMux I__314 (
            .O(N__2924),
            .I(N__2918));
    Span12Mux_v I__313 (
            .O(N__2921),
            .I(N__2915));
    Span12Mux_h I__312 (
            .O(N__2918),
            .I(N__2912));
    Span12Mux_h I__311 (
            .O(N__2915),
            .I(N__2907));
    Span12Mux_v I__310 (
            .O(N__2912),
            .I(N__2907));
    Span12Mux_h I__309 (
            .O(N__2907),
            .I(N__2904));
    Odrv12 I__308 (
            .O(N__2904),
            .I(D_LM_040_in_4));
    IoInMux I__307 (
            .O(N__2901),
            .I(N__2898));
    LocalMux I__306 (
            .O(N__2898),
            .I(N__2895));
    Span4Mux_s3_v I__305 (
            .O(N__2895),
            .I(N__2892));
    Span4Mux_h I__304 (
            .O(N__2892),
            .I(N__2889));
    Odrv4 I__303 (
            .O(N__2889),
            .I(un1_D_UU_040_4));
    InMux I__302 (
            .O(N__2886),
            .I(N__2883));
    LocalMux I__301 (
            .O(N__2883),
            .I(N__2880));
    Span4Mux_v I__300 (
            .O(N__2880),
            .I(N__2877));
    Sp12to4 I__299 (
            .O(N__2877),
            .I(N__2874));
    Span12Mux_h I__298 (
            .O(N__2874),
            .I(N__2871));
    Span12Mux_h I__297 (
            .O(N__2871),
            .I(N__2868));
    Odrv12 I__296 (
            .O(N__2868),
            .I(D_UM_040_in_4));
    IoInMux I__295 (
            .O(N__2865),
            .I(N__2862));
    LocalMux I__294 (
            .O(N__2862),
            .I(N__2858));
    InMux I__293 (
            .O(N__2861),
            .I(N__2855));
    Span4Mux_s2_h I__292 (
            .O(N__2858),
            .I(N__2852));
    LocalMux I__291 (
            .O(N__2855),
            .I(N__2849));
    Span4Mux_v I__290 (
            .O(N__2852),
            .I(N__2846));
    Span12Mux_h I__289 (
            .O(N__2849),
            .I(N__2843));
    Sp12to4 I__288 (
            .O(N__2846),
            .I(N__2840));
    Span12Mux_v I__287 (
            .O(N__2843),
            .I(N__2837));
    Span12Mux_h I__286 (
            .O(N__2840),
            .I(N__2834));
    Span12Mux_v I__285 (
            .O(N__2837),
            .I(N__2831));
    Span12Mux_h I__284 (
            .O(N__2834),
            .I(N__2828));
    Odrv12 I__283 (
            .O(N__2831),
            .I(D_LL_040_in_4));
    Odrv12 I__282 (
            .O(N__2828),
            .I(D_LL_040_in_4));
    IoInMux I__281 (
            .O(N__2823),
            .I(N__2820));
    LocalMux I__280 (
            .O(N__2820),
            .I(N__2817));
    Span4Mux_s2_h I__279 (
            .O(N__2817),
            .I(N__2814));
    Span4Mux_h I__278 (
            .O(N__2814),
            .I(N__2811));
    Span4Mux_h I__277 (
            .O(N__2811),
            .I(N__2808));
    Odrv4 I__276 (
            .O(N__2808),
            .I(un1_D_UM_040_4));
    InMux I__275 (
            .O(N__2805),
            .I(N__2802));
    LocalMux I__274 (
            .O(N__2802),
            .I(N__2799));
    Span4Mux_v I__273 (
            .O(N__2799),
            .I(N__2796));
    Sp12to4 I__272 (
            .O(N__2796),
            .I(N__2793));
    Span12Mux_h I__271 (
            .O(N__2793),
            .I(N__2790));
    Odrv12 I__270 (
            .O(N__2790),
            .I(D_LL_AMIGA_in_1));
    IoInMux I__269 (
            .O(N__2787),
            .I(N__2784));
    LocalMux I__268 (
            .O(N__2784),
            .I(N__2781));
    IoSpan4Mux I__267 (
            .O(N__2781),
            .I(N__2778));
    Span4Mux_s3_h I__266 (
            .O(N__2778),
            .I(N__2775));
    Span4Mux_v I__265 (
            .O(N__2775),
            .I(N__2772));
    Span4Mux_h I__264 (
            .O(N__2772),
            .I(N__2769));
    Sp12to4 I__263 (
            .O(N__2769),
            .I(N__2766));
    Odrv12 I__262 (
            .O(N__2766),
            .I(un2_D_LL_AMIGA_1));
    IoInMux I__261 (
            .O(N__2763),
            .I(N__2760));
    LocalMux I__260 (
            .O(N__2760),
            .I(N__2757));
    Span12Mux_s1_v I__259 (
            .O(N__2757),
            .I(N__2754));
    Odrv12 I__258 (
            .O(N__2754),
            .I(CPUBGn_c_i_0));
    InMux I__257 (
            .O(N__2751),
            .I(N__2748));
    LocalMux I__256 (
            .O(N__2748),
            .I(N__2745));
    Span4Mux_v I__255 (
            .O(N__2745),
            .I(N__2742));
    Sp12to4 I__254 (
            .O(N__2742),
            .I(N__2739));
    Span12Mux_h I__253 (
            .O(N__2739),
            .I(N__2736));
    Odrv12 I__252 (
            .O(N__2736),
            .I(D_LL_AMIGA_in_5));
    IoInMux I__251 (
            .O(N__2733),
            .I(N__2730));
    LocalMux I__250 (
            .O(N__2730),
            .I(N__2727));
    Span12Mux_s8_h I__249 (
            .O(N__2727),
            .I(N__2724));
    Span12Mux_h I__248 (
            .O(N__2724),
            .I(N__2721));
    Odrv12 I__247 (
            .O(N__2721),
            .I(un2_D_LL_AMIGA_5));
    InMux I__246 (
            .O(N__2718),
            .I(N__2715));
    LocalMux I__245 (
            .O(N__2715),
            .I(N__2712));
    Span12Mux_v I__244 (
            .O(N__2712),
            .I(N__2709));
    Odrv12 I__243 (
            .O(N__2709),
            .I(D_LL_AMIGA_in_7));
    IoInMux I__242 (
            .O(N__2706),
            .I(N__2703));
    LocalMux I__241 (
            .O(N__2703),
            .I(N__2700));
    Span4Mux_s2_h I__240 (
            .O(N__2700),
            .I(N__2697));
    Sp12to4 I__239 (
            .O(N__2697),
            .I(N__2694));
    Span12Mux_v I__238 (
            .O(N__2694),
            .I(N__2691));
    Span12Mux_h I__237 (
            .O(N__2691),
            .I(N__2688));
    Odrv12 I__236 (
            .O(N__2688),
            .I(un2_D_LL_AMIGA_7));
    IoInMux I__235 (
            .O(N__2685),
            .I(N__2682));
    LocalMux I__234 (
            .O(N__2682),
            .I(N__2679));
    Span4Mux_s0_v I__233 (
            .O(N__2679),
            .I(N__2676));
    Sp12to4 I__232 (
            .O(N__2676),
            .I(N__2673));
    Span12Mux_h I__231 (
            .O(N__2673),
            .I(N__2670));
    Span12Mux_v I__230 (
            .O(N__2670),
            .I(N__2667));
    Span12Mux_v I__229 (
            .O(N__2667),
            .I(N__2664));
    Odrv12 I__228 (
            .O(N__2664),
            .I(TAn_in));
    IoInMux I__227 (
            .O(N__2661),
            .I(N__2658));
    LocalMux I__226 (
            .O(N__2658),
            .I(N__2655));
    Odrv12 I__225 (
            .O(N__2655),
            .I(RESETn_c_i));
    INV \INVU111_CYCLE_SM.TS_OUTC  (
            .O(\INVU111_CYCLE_SM.TS_OUTC_net ),
            .I(N__7133));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__2661),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_1_10_1.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_1_10_1.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_1_10_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_1_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6214),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_1  (
            .in0(N__3467),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3813),
            .lcout(U111_CYCLE_SM_A_AMIGA_0_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_5  (
            .in0(N__3069),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3812),
            .lcout(A_AMIGA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_7_10_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_7_10_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_7_10_3  (
            .in0(N__8134),
            .in1(N__3042),
            .in2(_gnd_net_),
            .in3(N__3026),
            .lcout(un1_D_UM_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_7_20_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_7_20_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_7_20_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_7_20_6  (
            .in0(N__8214),
            .in1(N__2964),
            .in2(_gnd_net_),
            .in3(N__2930),
            .lcout(un1_D_UU_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_7_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_7_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_7_20_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_7_20_7  (
            .in0(N__2886),
            .in1(N__2861),
            .in2(_gnd_net_),
            .in3(N__8213),
            .lcout(un1_D_UM_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_8_3_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_8_3_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_8_3_4  (
            .in0(N__7014),
            .in1(N__2805),
            .in2(_gnd_net_),
            .in3(N__8174),
            .lcout(un2_D_LL_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TSn_obuft_RNO_LC_8_3_5.C_ON=1'b0;
    defparam TSn_obuft_RNO_LC_8_3_5.SEQ_MODE=4'b0000;
    defparam TSn_obuft_RNO_LC_8_3_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 TSn_obuft_RNO_LC_8_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7791),
            .lcout(CPUBGn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_8_6_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_8_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_8_6_4  (
            .in0(N__2751),
            .in1(N__7952),
            .in2(_gnd_net_),
            .in3(N__8130),
            .lcout(un2_D_LL_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_8_7_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_8_7_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_8_7_2  (
            .in0(N__2718),
            .in1(N__8426),
            .in2(_gnd_net_),
            .in3(N__8129),
            .lcout(un2_D_LL_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_8_7_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_8_7_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_8_7_5  (
            .in0(N__4142),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3477),
            .lcout(\U111_CYCLE_SM.N_141 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_8_11_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_8_11_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_8_11_2  (
            .in0(N__3450),
            .in1(N__4322),
            .in2(_gnd_net_),
            .in3(N__8136),
            .lcout(N_108),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_8_11_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_8_11_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_8_11_6  (
            .in0(N__3423),
            .in1(N__6728),
            .in2(_gnd_net_),
            .in3(N__8135),
            .lcout(N_110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_8_12_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_8_12_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_8_12_3  (
            .in0(N__3387),
            .in1(N__4656),
            .in2(_gnd_net_),
            .in3(N__8137),
            .lcout(N_111),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_8_12_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_8_12_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_8_12_6  (
            .in0(N__8138),
            .in1(N__3357),
            .in2(_gnd_net_),
            .in3(N__3332),
            .lcout(un1_D_UM_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_8_20_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_8_20_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_8_20_4  (
            .in0(N__8211),
            .in1(N__3279),
            .in2(_gnd_net_),
            .in3(N__3257),
            .lcout(un1_D_UU_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_8_20_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_8_20_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_8_20_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_8_20_6  (
            .in0(N__8212),
            .in1(N__3192),
            .in2(_gnd_net_),
            .in3(N__3167),
            .lcout(un1_D_UU_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_9_3_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_9_3_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_9_3_3  (
            .in0(N__8168),
            .in1(N__5942),
            .in2(_gnd_net_),
            .in3(N__3114),
            .lcout(un2_D_LL_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_9_3_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_9_3_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_9_3_6  (
            .in0(N__3786),
            .in1(N__6411),
            .in2(_gnd_net_),
            .in3(N__8167),
            .lcout(un2_D_LL_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_9_10_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_9_10_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_9_10_0  (
            .in0(N__3749),
            .in1(N__3714),
            .in2(_gnd_net_),
            .in3(N__8025),
            .lcout(un1_D_UM_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_9_10_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_9_10_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_9_10_5  (
            .in0(N__8026),
            .in1(N__6038),
            .in2(_gnd_net_),
            .in3(N__3675),
            .lcout(N_112),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_BUFFERS.DMA_EN_i_0_LC_9_20_3 .C_ON=1'b0;
    defparam \U111_BUFFERS.DMA_EN_i_0_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_BUFFERS.DMA_EN_i_0_LC_9_20_3 .LUT_INIT=16'b1011101110111011;
    LogicCell40 \U111_BUFFERS.DMA_EN_i_0_LC_9_20_3  (
            .in0(N__3604),
            .in1(N__7805),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_96),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_BUFFERS.N_94_i_LC_9_20_6 .C_ON=1'b0;
    defparam \U111_BUFFERS.N_94_i_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \U111_BUFFERS.N_94_i_LC_9_20_6 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U111_BUFFERS.N_94_i_LC_9_20_6  (
            .in0(N__7806),
            .in1(N__3605),
            .in2(_gnd_net_),
            .in3(N__6875),
            .lcout(N_94_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_BUFFERS.un1_DMA_EN_0_0_LC_9_20_7 .C_ON=1'b0;
    defparam \U111_BUFFERS.un1_DMA_EN_0_0_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_BUFFERS.un1_DMA_EN_0_0_LC_9_20_7 .LUT_INIT=16'b0001000110101010;
    LogicCell40 \U111_BUFFERS.un1_DMA_EN_0_0_LC_9_20_7  (
            .in0(N__7725),
            .in1(N__3606),
            .in2(_gnd_net_),
            .in3(N__7807),
            .lcout(BUFDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_10_8_4.C_ON=1'b0;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_10_8_4.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_10_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK40_THRU_LUT4_0_LC_10_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7143),
            .lcout(GB_BUFFER_CLK40_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_LC_10_9_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_LC_10_9_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TS_EN_LC_10_9_0 .LUT_INIT=16'b1111111000110010;
    LogicCell40 \U111_CYCLE_SM.TS_EN_LC_10_9_0  (
            .in0(N__4122),
            .in1(N__4086),
            .in2(N__5100),
            .in3(N__4065),
            .lcout(\U111_CYCLE_SM.TS_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7135),
            .ce(),
            .sr(N__6294));
    defparam \U111_CYCLE_SM.FLIP_WORD_LC_10_9_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_LC_10_9_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.FLIP_WORD_LC_10_9_4 .LUT_INIT=16'b1111000011101110;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_LC_10_9_4  (
            .in0(N__5096),
            .in1(N__8024),
            .in2(N__3492),
            .in3(N__4177),
            .lcout(\U111_CYCLE_SM.FLIP_WORDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7135),
            .ce(),
            .sr(N__6294));
    defparam \U111_CYCLE_SM.TS_OUT_LC_10_10_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_OUT_LC_10_10_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TS_OUT_LC_10_10_3 .LUT_INIT=16'b0111011101010111;
    LogicCell40 \U111_CYCLE_SM.TS_OUT_LC_10_10_3  (
            .in0(N__6263),
            .in1(N__4064),
            .in2(N__6876),
            .in3(N__5220),
            .lcout(TS_OUT),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.TS_OUTC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_10_16_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_10_16_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_10_16_4  (
            .in0(N__8149),
            .in1(N__4493),
            .in2(_gnd_net_),
            .in3(N__4053),
            .lcout(N_106),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_10_16_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_10_16_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_10_16_7  (
            .in0(N__4014),
            .in1(N__5613),
            .in2(_gnd_net_),
            .in3(N__8148),
            .lcout(N_107),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_10_18_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_10_18_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_10_18_7  (
            .in0(N__3981),
            .in1(N__3966),
            .in2(_gnd_net_),
            .in3(N__8186),
            .lcout(un1_D_UM_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_11_1_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_11_1_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_11_1_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_11_1_2  (
            .in0(N__3903),
            .in1(N__8206),
            .in2(_gnd_net_),
            .in3(N__8616),
            .lcout(un2_D_LL_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LBENn_c_sbtinv_LC_11_1_5.C_ON=1'b0;
    defparam LBENn_c_sbtinv_LC_11_1_5.SEQ_MODE=4'b0000;
    defparam LBENn_c_sbtinv_LC_11_1_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 LBENn_c_sbtinv_LC_11_1_5 (
            .in0(N__6835),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(LBENn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_11_7_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_11_7_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_11_7_3  (
            .in0(N__8067),
            .in1(N__5811),
            .in2(_gnd_net_),
            .in3(N__3852),
            .lcout(un2_D_LM_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.un1_CYCLE_STATE_1_i_i_o2_LC_11_7_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.un1_CYCLE_STATE_1_i_i_o2_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.un1_CYCLE_STATE_1_i_i_o2_LC_11_7_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U111_CYCLE_SM.un1_CYCLE_STATE_1_i_i_o2_LC_11_7_6  (
            .in0(N__6484),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5154),
            .lcout(\U111_CYCLE_SM.N_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A2_EN_LC_11_8_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A2_EN_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.A2_EN_LC_11_8_1 .LUT_INIT=16'b1110110011101110;
    LogicCell40 \U111_CYCLE_SM.A2_EN_LC_11_8_1  (
            .in0(N__3797),
            .in1(N__5093),
            .in2(N__4105),
            .in3(N__4851),
            .lcout(\U111_CYCLE_SM.A2_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7136),
            .ce(),
            .sr(N__6297));
    defparam \U111_CYCLE_SM.BURST_RNILNBJ_LC_11_9_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_RNILNBJ_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.BURST_RNILNBJ_LC_11_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U111_CYCLE_SM.BURST_RNILNBJ_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__4870),
            .in2(_gnd_net_),
            .in3(N__4848),
            .lcout(\U111_CYCLE_SM.N_179 ),
            .ltout(\U111_CYCLE_SM.N_179_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_11_9_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_11_9_1 .LUT_INIT=16'b1100110001000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_1_LC_11_9_1  (
            .in0(N__4106),
            .in1(N__6252),
            .in2(N__4116),
            .in3(N__5051),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7134),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_DIS_RNO_0_LC_11_9_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_RNO_0_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_DIS_RNO_0_LC_11_9_2 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_RNO_0_LC_11_9_2  (
            .in0(N__4154),
            .in1(N__4192),
            .in2(_gnd_net_),
            .in3(N__4175),
            .lcout(\U111_CYCLE_SM.N_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_11_9_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_11_9_3 .LUT_INIT=16'b1111011101110111;
    LogicCell40 \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_11_9_3  (
            .in0(N__4869),
            .in1(N__6618),
            .in2(N__4215),
            .in3(N__4277),
            .lcout(\U111_CYCLE_SM.N_101 ),
            .ltout(\U111_CYCLE_SM.N_101_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_11_9_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_11_9_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_11_9_4  (
            .in0(N__5158),
            .in1(N__4890),
            .in2(N__4113),
            .in3(N__5127),
            .lcout(\U111_CYCLE_SM.N_133 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_9_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_9_5 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_9_5  (
            .in0(N__5128),
            .in1(N__4849),
            .in2(N__4110),
            .in3(N__6335),
            .lcout(\U111_CYCLE_SM.N_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_11_9_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_11_9_6 .LUT_INIT=16'b0101111101011101;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_11_9_6  (
            .in0(N__6498),
            .in1(N__4080),
            .in2(N__5162),
            .in3(N__4891),
            .lcout(),
            .ltout(\U111_CYCLE_SM.N_12_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_2_LC_11_9_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_2_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_2_LC_11_9_7 .LUT_INIT=16'b1010111000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_2_LC_11_9_7  (
            .in0(N__4176),
            .in1(N__5130),
            .in2(N__4074),
            .in3(N__6253),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7134),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_DIS_LC_11_10_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TA_DIS_LC_11_10_0 .LUT_INIT=16'b0001000011111110;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_LC_11_10_0  (
            .in0(N__5094),
            .in1(N__4179),
            .in2(N__6940),
            .in3(N__4071),
            .lcout(\U111_CYCLE_SM.TA_DISZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7129),
            .ce(),
            .sr(N__6293));
    defparam \U111_CYCLE_SM.BURST_LC_11_10_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.BURST_LC_11_10_1 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U111_CYCLE_SM.BURST_LC_11_10_1  (
            .in0(N__5048),
            .in1(N__4265),
            .in2(N__4242),
            .in3(N__4872),
            .lcout(\U111_CYCLE_SM.BURSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7129),
            .ce(),
            .sr(N__6293));
    defparam \U111_CYCLE_SM.BURST_COUNT_1_LC_11_10_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_COUNT_1_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.BURST_COUNT_1_LC_11_10_3 .LUT_INIT=16'b0000100100001100;
    LogicCell40 \U111_CYCLE_SM.BURST_COUNT_1_LC_11_10_3  (
            .in0(N__6185),
            .in1(N__4278),
            .in2(N__5052),
            .in3(N__4214),
            .lcout(\U111_CYCLE_SM.BURST_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7129),
            .ce(),
            .sr(N__6293));
    defparam \U111_CYCLE_SM.LW_TRANS_LC_11_10_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_TRANS_LC_11_10_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LW_TRANS_LC_11_10_4 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \U111_CYCLE_SM.LW_TRANS_LC_11_10_4  (
            .in0(N__4266),
            .in1(N__4241),
            .in2(N__4197),
            .in3(N__5049),
            .lcout(\U111_CYCLE_SM.LW_TRANSZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7129),
            .ce(),
            .sr(N__6293));
    defparam \U111_CYCLE_SM.BURST_COUNT_0_LC_11_10_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_COUNT_0_LC_11_10_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.BURST_COUNT_0_LC_11_10_5 .LUT_INIT=16'b0100010000010001;
    LogicCell40 \U111_CYCLE_SM.BURST_COUNT_0_LC_11_10_5  (
            .in0(N__5043),
            .in1(N__6184),
            .in2(_gnd_net_),
            .in3(N__4213),
            .lcout(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7129),
            .ce(),
            .sr(N__6293));
    defparam \U111_CYCLE_SM.PORT_MISMATCH_LC_11_10_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.PORT_MISMATCH_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.PORT_MISMATCH_LC_11_10_6 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \U111_CYCLE_SM.PORT_MISMATCH_LC_11_10_6  (
            .in0(N__4193),
            .in1(N__4178),
            .in2(N__4896),
            .in3(N__4155),
            .lcout(\U111_CYCLE_SM.PORT_MISMATCHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7129),
            .ce(),
            .sr(N__6293));
    defparam \U111_CYCLE_SM.CYCLE_EN_LC_11_10_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_EN_LC_11_10_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_EN_LC_11_10_7 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \U111_CYCLE_SM.CYCLE_EN_LC_11_10_7  (
            .in0(N__5044),
            .in1(N__5503),
            .in2(_gnd_net_),
            .in3(N__6337),
            .lcout(\U111_CYCLE_SM.CYCLE_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7129),
            .ce(),
            .sr(N__6293));
    defparam \U111_CYCLE_SM.UU_LATCHED_5_LC_11_11_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_5_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_5_LC_11_11_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_5_LC_11_11_0  (
            .in0(N__7882),
            .in1(N__4937),
            .in2(N__4329),
            .in3(N__6157),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7125),
            .ce(),
            .sr(N__6295));
    defparam \U111_CYCLE_SM.UU_LATCHED_2_LC_11_11_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_2_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_2_LC_11_11_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_2_LC_11_11_2  (
            .in0(N__7880),
            .in1(N__4601),
            .in2(N__4652),
            .in3(N__6155),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7125),
            .ce(),
            .sr(N__6295));
    defparam \U111_CYCLE_SM.UU_LATCHED_7_LC_11_11_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_7_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_7_LC_11_11_4 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_7_LC_11_11_4  (
            .in0(N__7883),
            .in1(N__4445),
            .in2(N__4494),
            .in3(N__6158),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7125),
            .ce(),
            .sr(N__6295));
    defparam \U111_CYCLE_SM.TS_DELAY_LC_11_11_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_DELAY_LC_11_11_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.TS_DELAY_LC_11_11_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.TS_DELAY_LC_11_11_6  (
            .in0(N__4800),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.TS_DELAYZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7125),
            .ce(),
            .sr(N__6295));
    defparam \U111_CYCLE_SM.UU_LATCHED_4_LC_11_11_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_4_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_4_LC_11_11_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_4_LC_11_11_7  (
            .in0(N__6156),
            .in1(N__4568),
            .in2(N__4557),
            .in3(N__7881),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7125),
            .ce(),
            .sr(N__6295));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_11_13_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_11_13_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_11_13_1  (
            .in0(N__4782),
            .in1(N__4550),
            .in2(_gnd_net_),
            .in3(N__8139),
            .lcout(N_109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_11_20_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_11_20_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_11_20_0  (
            .in0(N__8208),
            .in1(N__4743),
            .in2(_gnd_net_),
            .in3(N__4724),
            .lcout(un1_D_UU_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_RNINJKT_2_LC_11_20_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNINJKT_2_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNINJKT_2_LC_11_20_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_RNINJKT_2_LC_11_20_2  (
            .in0(N__7340),
            .in1(N__4648),
            .in2(_gnd_net_),
            .in3(N__4605),
            .lcout(N_118),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIRNKT_4_LC_11_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIRNKT_4_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIRNKT_4_LC_11_20_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_RNIRNKT_4_LC_11_20_3  (
            .in0(N__4575),
            .in1(N__4538),
            .in2(_gnd_net_),
            .in3(N__7341),
            .lcout(N_116),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_RNI1UKT_7_LC_11_20_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNI1UKT_7_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNI1UKT_7_LC_11_20_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_RNI1UKT_7_LC_11_20_4  (
            .in0(N__7339),
            .in1(N__4486),
            .in2(_gnd_net_),
            .in3(N__4452),
            .lcout(N_113),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_11_20_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_11_20_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_11_20_5  (
            .in0(N__4406),
            .in1(N__4365),
            .in2(_gnd_net_),
            .in3(N__8209),
            .lcout(un1_D_UU_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_RNITPKT_5_LC_11_20_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNITPKT_5_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNITPKT_5_LC_11_20_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_RNITPKT_5_LC_11_20_6  (
            .in0(N__7342),
            .in1(N__4309),
            .in2(_gnd_net_),
            .in3(N__4947),
            .lcout(N_115),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_12_8_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_12_8_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(N__6491),
            .in2(_gnd_net_),
            .in3(N__5181),
            .lcout(),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_srsts_i_i_o2_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_5_LC_12_8_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_5_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_5_LC_12_8_2 .LUT_INIT=16'b1000101010001000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_5_LC_12_8_2  (
            .in0(N__6255),
            .in1(N__4902),
            .in2(N__4905),
            .in3(N__4850),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7132),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_8_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_8_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_8_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_8_6  (
            .in0(N__6254),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5084),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7132),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_3_LC_12_9_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_3_LC_12_9_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_3_LC_12_9_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_3_LC_12_9_0  (
            .in0(N__6269),
            .in1(N__4892),
            .in2(_gnd_net_),
            .in3(N__6186),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7128),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_9_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_9_2 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_9_2  (
            .in0(N__6502),
            .in1(N__4846),
            .in2(_gnd_net_),
            .in3(N__5129),
            .lcout(\U111_CYCLE_SM.N_131 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_12_9_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_12_9_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_12_9_4  (
            .in0(N__5182),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4871),
            .lcout(),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_a3_2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_9_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_9_5 .LUT_INIT=16'b1111111110110011;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_9_5  (
            .in0(N__4847),
            .in1(N__6270),
            .in2(N__4818),
            .in3(N__4815),
            .lcout(),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_9_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_9_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_9_6 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_9_6  (
            .in0(N__6361),
            .in1(N__4809),
            .in2(N__4803),
            .in3(N__6336),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7128),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_DELAY_RNIDR7G_LC_12_10_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_DELAY_RNIDR7G_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_DELAY_RNIDR7G_LC_12_10_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U111_CYCLE_SM.TS_DELAY_RNIDR7G_LC_12_10_0  (
            .in0(N__6839),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5219),
            .lcout(\U111_CYCLE_SM.un4_TS_OUT_i_0 ),
            .ltout(\U111_CYCLE_SM.un4_TS_OUT_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI9UTM_0_LC_12_10_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI9UTM_0_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI9UTM_0_LC_12_10_1 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNI9UTM_0_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5208),
            .in3(N__6334),
            .lcout(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_10_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_10_3 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_10_3  (
            .in0(N__5189),
            .in1(N__6503),
            .in2(_gnd_net_),
            .in3(N__5126),
            .lcout(\U111_CYCLE_SM.N_99 ),
            .ltout(\U111_CYCLE_SM.N_99_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_0_2_LC_12_10_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_0_2_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_0_2_LC_12_10_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_0_2_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5103),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.N_99_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LATCH_EN_RNO_0_LC_12_10_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LATCH_EN_RNO_0_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LATCH_EN_RNO_0_LC_12_10_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \U111_CYCLE_SM.LATCH_EN_RNO_0_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(N__6333),
            .in2(_gnd_net_),
            .in3(N__7863),
            .lcout(\U111_CYCLE_SM.N_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LATCH_EN_LC_12_11_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LATCH_EN_LC_12_11_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LATCH_EN_LC_12_11_3 .LUT_INIT=16'b0011001101110010;
    LogicCell40 \U111_CYCLE_SM.LATCH_EN_LC_12_11_3  (
            .in0(N__5095),
            .in1(N__5058),
            .in2(N__7280),
            .in3(N__5050),
            .lcout(\U111_CYCLE_SM.LATCH_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7123),
            .ce(),
            .sr(N__6298));
    defparam \U111_CYCLE_SM.CYCLE_EN_RNI26B3_LC_12_11_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_EN_RNI26B3_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_EN_RNI26B3_LC_12_11_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U111_CYCLE_SM.CYCLE_EN_RNI26B3_LC_12_11_6  (
            .in0(N__5538),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5504),
            .lcout(CPUBGn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_LC_12_12_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_LC_12_12_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_LC_12_12_2 .LUT_INIT=16'b0010001000101110;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_LC_12_12_2  (
            .in0(N__5486),
            .in1(N__6344),
            .in2(N__7720),
            .in3(N__6366),
            .lcout(\U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7122),
            .ce(),
            .sr(N__6299));
    defparam \U111_CYCLE_SM.UU_LATCHED_6_LC_12_12_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_6_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_6_LC_12_12_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_6_LC_12_12_7  (
            .in0(N__5624),
            .in1(N__7876),
            .in2(N__5609),
            .in3(N__6159),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7122),
            .ce(),
            .sr(N__6299));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_12_18_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_12_18_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_12_18_0  (
            .in0(N__5012),
            .in1(N__4983),
            .in2(_gnd_net_),
            .in3(N__8207),
            .lcout(un1_D_UU_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TS_CPUn_iobuf_RNO_LC_12_18_7.C_ON=1'b0;
    defparam TS_CPUn_iobuf_RNO_LC_12_18_7.SEQ_MODE=4'b0000;
    defparam TS_CPUn_iobuf_RNO_LC_12_18_7.LUT_INIT=16'b0101010100000000;
    LogicCell40 TS_CPUn_iobuf_RNO_LC_12_18_7 (
            .in0(N__7775),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5753),
            .lcout(TSnz),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_12_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_12_20_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_12_20_1  (
            .in0(N__5699),
            .in1(N__5664),
            .in2(_gnd_net_),
            .in3(N__8210),
            .lcout(un1_D_UU_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIVRKT_6_LC_12_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIVRKT_6_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIVRKT_6_LC_12_20_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_RNIVRKT_6_LC_12_20_3  (
            .in0(N__5631),
            .in1(N__5602),
            .in2(_gnd_net_),
            .in3(N__7309),
            .lcout(N_114),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_20_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_20_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_20_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_1_LC_13_10_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_1_LC_13_10_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_1_LC_13_10_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_1_LC_13_10_1  (
            .in0(N__5987),
            .in1(N__7865),
            .in2(N__6039),
            .in3(N__6150),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7130),
            .ce(),
            .sr(N__6296));
    defparam \U111_CYCLE_SM.UU_LATCHED_3_LC_13_10_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_3_LC_13_10_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_3_LC_13_10_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_3_LC_13_10_3  (
            .in0(N__6743),
            .in1(N__7866),
            .in2(N__6732),
            .in3(N__6151),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7130),
            .ce(),
            .sr(N__6296));
    defparam \U111_CYCLE_SM.UU_LATCHED_0_LC_13_10_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_0_LC_13_10_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_0_LC_13_10_5 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_0_LC_13_10_5  (
            .in0(N__5822),
            .in1(N__7864),
            .in2(N__5810),
            .in3(N__6149),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7130),
            .ce(),
            .sr(N__6296));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_RNINRNR_LC_13_11_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_RNINRNR_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_RNINRNR_LC_13_11_0 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_RNINRNR_LC_13_11_0  (
            .in0(N__7719),
            .in1(N__5537),
            .in2(N__5514),
            .in3(N__5487),
            .lcout(U111_CYCLE_SM_OFFBOARD_EN_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_13_11_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_13_11_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_13_11_2 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_13_11_2  (
            .in0(N__7862),
            .in1(N__6365),
            .in2(N__7724),
            .in3(N__6345),
            .lcout(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7126),
            .ce(),
            .sr(N__6300));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTO81_LC_13_11_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTO81_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTO81_LC_13_11_3 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTO81_LC_13_11_3  (
            .in0(N__6262),
            .in1(N__7861),
            .in2(_gnd_net_),
            .in3(N__6183),
            .lcout(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81 ),
            .ltout(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNI0BVS1_LC_13_11_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNI0BVS1_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNI0BVS1_LC_13_11_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNI0BVS1_LC_13_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6162),
            .in3(N__6148),
            .lcout(\U111_CYCLE_SM.N_99_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_13_12_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_13_12_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_13_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5943),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7124),
            .ce(N__7085),
            .sr(N__7039));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_13_15_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_13_15_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_13_15_1  (
            .in0(N__6117),
            .in1(N__6098),
            .in2(_gnd_net_),
            .in3(N__8197),
            .lcout(un1_D_UM_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_RNILHKT_1_LC_13_15_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNILHKT_1_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNILHKT_1_LC_13_15_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_RNILHKT_1_LC_13_15_3  (
            .in0(N__7343),
            .in1(N__6028),
            .in2(_gnd_net_),
            .in3(N__5991),
            .lcout(N_119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_13_18_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_13_18_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_13_18_0  (
            .in0(N__7333),
            .in1(N__5955),
            .in2(_gnd_net_),
            .in3(N__5932),
            .lcout(un1_D_UM_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_13_18_5.C_ON=1'b0;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_13_18_5.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_13_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK80_THRU_LUT4_0_LC_13_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5868),
            .lcout(GB_BUFFER_CLK80_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIJFKT_0_LC_13_20_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIJFKT_0_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIJFKT_0_LC_13_20_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_RNIJFKT_0_LC_13_20_0  (
            .in0(N__5829),
            .in1(N__5797),
            .in2(_gnd_net_),
            .in3(N__7348),
            .lcout(un1_D_UU_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIPLKT_3_LC_13_20_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIPLKT_3_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIPLKT_3_LC_13_20_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_RNIPLKT_3_LC_13_20_2  (
            .in0(N__6747),
            .in1(N__6718),
            .in2(_gnd_net_),
            .in3(N__7349),
            .lcout(N_117),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_14_1_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_14_1_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_14_1_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_14_1_0  (
            .in0(N__6654),
            .in1(N__7185),
            .in2(_gnd_net_),
            .in3(N__8173),
            .lcout(un2_D_LL_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TBI_CPUn_0_i_LC_14_1_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TBI_CPUn_0_i_LC_14_1_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TBI_CPUn_0_i_LC_14_1_5 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U111_CYCLE_SM.TBI_CPUn_0_i_LC_14_1_5  (
            .in0(N__6608),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6849),
            .lcout(U111_CYCLE_SM_TBI_CPUn_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_14_6_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_14_6_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_14_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_14_6_7  (
            .in0(N__6576),
            .in1(N__7221),
            .in2(_gnd_net_),
            .in3(N__8172),
            .lcout(un2_D_LL_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_14_10_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_14_10_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_14_10_5  (
            .in0(N__7320),
            .in1(N__6372),
            .in2(_gnd_net_),
            .in3(N__6401),
            .lcout(un1_D_UM_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_14_10_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_14_10_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_14_10_6  (
            .in0(N__7178),
            .in1(N__7149),
            .in2(_gnd_net_),
            .in3(N__7319),
            .lcout(un1_D_UM_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_DIS_RNI576J_LC_14_10_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_RNI576J_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_DIS_RNI576J_LC_14_10_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_RNI576J_LC_14_10_7  (
            .in0(_gnd_net_),
            .in1(N__6504),
            .in2(_gnd_net_),
            .in3(N__6941),
            .lcout(U111_CYCLE_SM_TEA_CPUn_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_14_11_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_14_11_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_14_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6400),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7131),
            .ce(N__7075),
            .sr(N__7046));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_14_11_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_14_11_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_14_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_14_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7177),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7131),
            .ce(N__7075),
            .sr(N__7046));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_14_12_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_14_12_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_14_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_14_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8615),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7127),
            .ce(N__7086),
            .sr(N__7047));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_14_12_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_14_12_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_14_12_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_14_12_3  (
            .in0(N__7007),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7127),
            .ce(N__7086),
            .sr(N__7047));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_14_12_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_14_12_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_14_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7210),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7127),
            .ce(N__7086),
            .sr(N__7047));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_14_12_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_14_12_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_14_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_14_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8430),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7127),
            .ce(N__7086),
            .sr(N__7047));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_14_12_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_14_12_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_14_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_14_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7953),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7127),
            .ce(N__7086),
            .sr(N__7047));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_14_13_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_14_13_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_14_13_2  (
            .in0(N__7006),
            .in1(N__6972),
            .in2(_gnd_net_),
            .in3(N__7321),
            .lcout(un1_D_UM_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_14_13_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_14_13_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_14_13_4  (
            .in0(N__6861),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6945),
            .lcout(N_64),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TCI_CPUn_0_i_LC_14_13_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TCI_CPUn_0_i_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TCI_CPUn_0_i_LC_14_13_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \U111_CYCLE_SM.TCI_CPUn_0_i_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(N__6897),
            .in2(_gnd_net_),
            .in3(N__6862),
            .lcout(U111_CYCLE_SM_TCI_CPUn_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_14_14_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_14_14_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_14_14_7  (
            .in0(N__8608),
            .in1(N__8565),
            .in2(_gnd_net_),
            .in3(N__7323),
            .lcout(un1_D_UM_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_14_19_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_14_19_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_14_19_2  (
            .in0(N__8531),
            .in1(N__8484),
            .in2(_gnd_net_),
            .in3(N__8215),
            .lcout(un1_D_UM_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_14_19_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_14_19_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_14_19_7  (
            .in0(N__8442),
            .in1(N__8422),
            .in2(_gnd_net_),
            .in3(N__7344),
            .lcout(un1_D_UM_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_14_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_14_20_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_14_20_3  (
            .in0(N__8348),
            .in1(N__8319),
            .in2(_gnd_net_),
            .in3(N__8217),
            .lcout(un1_D_UU_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_14_20_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_14_20_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_14_20_5  (
            .in0(N__8283),
            .in1(N__8264),
            .in2(_gnd_net_),
            .in3(N__8216),
            .lcout(un1_D_UM_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_14_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_14_20_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_14_20_7  (
            .in0(N__7350),
            .in1(N__7965),
            .in2(_gnd_net_),
            .in3(N__7942),
            .lcout(un1_D_UM_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNI8QUM_LC_15_12_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNI8QUM_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNI8QUM_LC_15_12_3 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNI8QUM_LC_15_12_3  (
            .in0(N__7887),
            .in1(N__7769),
            .in2(_gnd_net_),
            .in3(N__7704),
            .lcout(N_60_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_15_12_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_15_12_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_15_12_5  (
            .in0(N__7322),
            .in1(N__7227),
            .in2(_gnd_net_),
            .in3(N__7211),
            .lcout(un1_D_UM_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U111_TOP

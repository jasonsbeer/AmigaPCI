// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Dec 16 2024 18:13:15

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    CMA,
    DRA,
    A,
    TSn,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    VBENn,
    CUMBEn,
    CLKRAM,
    C3,
    ASn,
    LDSn,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CASLn,
    RAMSPACEn,
    WEn,
    REGENn,
    DBRn,
    CLK40C,
    CLK40_IN,
    REGSPACEn,
    RAMENn,
    RASn,
    TACKn,
    C1);

    input [1:0] SIZ;
    output [10:0] CMA;
    input [9:0] DRA;
    input [20:0] A;
    input TSn;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    input C3;
    output ASn;
    output LDSn;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    input CASLn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    input DBRn;
    output CLK40C;
    input CLK40_IN;
    input REGSPACEn;
    output RAMENn;
    output RASn;
    output TACKn;
    input C1;

    wire N__9911;
    wire N__9910;
    wire N__9909;
    wire N__9902;
    wire N__9901;
    wire N__9900;
    wire N__9893;
    wire N__9892;
    wire N__9891;
    wire N__9884;
    wire N__9883;
    wire N__9882;
    wire N__9875;
    wire N__9874;
    wire N__9873;
    wire N__9866;
    wire N__9865;
    wire N__9864;
    wire N__9857;
    wire N__9856;
    wire N__9855;
    wire N__9848;
    wire N__9847;
    wire N__9846;
    wire N__9839;
    wire N__9838;
    wire N__9837;
    wire N__9830;
    wire N__9829;
    wire N__9828;
    wire N__9821;
    wire N__9820;
    wire N__9819;
    wire N__9812;
    wire N__9811;
    wire N__9810;
    wire N__9803;
    wire N__9802;
    wire N__9801;
    wire N__9794;
    wire N__9793;
    wire N__9792;
    wire N__9785;
    wire N__9784;
    wire N__9783;
    wire N__9776;
    wire N__9775;
    wire N__9774;
    wire N__9767;
    wire N__9766;
    wire N__9765;
    wire N__9758;
    wire N__9757;
    wire N__9756;
    wire N__9749;
    wire N__9748;
    wire N__9747;
    wire N__9740;
    wire N__9739;
    wire N__9738;
    wire N__9731;
    wire N__9730;
    wire N__9729;
    wire N__9722;
    wire N__9721;
    wire N__9720;
    wire N__9713;
    wire N__9712;
    wire N__9711;
    wire N__9704;
    wire N__9703;
    wire N__9702;
    wire N__9695;
    wire N__9694;
    wire N__9693;
    wire N__9686;
    wire N__9685;
    wire N__9684;
    wire N__9677;
    wire N__9676;
    wire N__9675;
    wire N__9668;
    wire N__9667;
    wire N__9666;
    wire N__9659;
    wire N__9658;
    wire N__9657;
    wire N__9650;
    wire N__9649;
    wire N__9648;
    wire N__9641;
    wire N__9640;
    wire N__9639;
    wire N__9632;
    wire N__9631;
    wire N__9630;
    wire N__9623;
    wire N__9622;
    wire N__9621;
    wire N__9614;
    wire N__9613;
    wire N__9612;
    wire N__9605;
    wire N__9604;
    wire N__9603;
    wire N__9596;
    wire N__9595;
    wire N__9594;
    wire N__9587;
    wire N__9586;
    wire N__9585;
    wire N__9578;
    wire N__9577;
    wire N__9576;
    wire N__9569;
    wire N__9568;
    wire N__9567;
    wire N__9560;
    wire N__9559;
    wire N__9558;
    wire N__9551;
    wire N__9550;
    wire N__9549;
    wire N__9542;
    wire N__9541;
    wire N__9540;
    wire N__9533;
    wire N__9532;
    wire N__9531;
    wire N__9524;
    wire N__9523;
    wire N__9522;
    wire N__9515;
    wire N__9514;
    wire N__9513;
    wire N__9506;
    wire N__9505;
    wire N__9504;
    wire N__9497;
    wire N__9496;
    wire N__9495;
    wire N__9488;
    wire N__9487;
    wire N__9486;
    wire N__9479;
    wire N__9478;
    wire N__9477;
    wire N__9470;
    wire N__9469;
    wire N__9468;
    wire N__9461;
    wire N__9460;
    wire N__9459;
    wire N__9452;
    wire N__9451;
    wire N__9450;
    wire N__9443;
    wire N__9442;
    wire N__9441;
    wire N__9434;
    wire N__9433;
    wire N__9432;
    wire N__9425;
    wire N__9424;
    wire N__9423;
    wire N__9416;
    wire N__9415;
    wire N__9414;
    wire N__9407;
    wire N__9406;
    wire N__9405;
    wire N__9398;
    wire N__9397;
    wire N__9396;
    wire N__9389;
    wire N__9388;
    wire N__9387;
    wire N__9380;
    wire N__9379;
    wire N__9378;
    wire N__9371;
    wire N__9370;
    wire N__9369;
    wire N__9362;
    wire N__9361;
    wire N__9360;
    wire N__9353;
    wire N__9352;
    wire N__9351;
    wire N__9344;
    wire N__9343;
    wire N__9342;
    wire N__9335;
    wire N__9334;
    wire N__9333;
    wire N__9326;
    wire N__9325;
    wire N__9324;
    wire N__9317;
    wire N__9316;
    wire N__9315;
    wire N__9308;
    wire N__9307;
    wire N__9306;
    wire N__9299;
    wire N__9298;
    wire N__9297;
    wire N__9290;
    wire N__9289;
    wire N__9288;
    wire N__9281;
    wire N__9280;
    wire N__9279;
    wire N__9272;
    wire N__9271;
    wire N__9270;
    wire N__9263;
    wire N__9262;
    wire N__9261;
    wire N__9254;
    wire N__9253;
    wire N__9252;
    wire N__9245;
    wire N__9244;
    wire N__9243;
    wire N__9236;
    wire N__9235;
    wire N__9234;
    wire N__9227;
    wire N__9226;
    wire N__9225;
    wire N__9218;
    wire N__9217;
    wire N__9216;
    wire N__9209;
    wire N__9208;
    wire N__9207;
    wire N__9200;
    wire N__9199;
    wire N__9198;
    wire N__9181;
    wire N__9180;
    wire N__9177;
    wire N__9174;
    wire N__9169;
    wire N__9166;
    wire N__9163;
    wire N__9160;
    wire N__9159;
    wire N__9158;
    wire N__9157;
    wire N__9156;
    wire N__9155;
    wire N__9154;
    wire N__9153;
    wire N__9152;
    wire N__9151;
    wire N__9150;
    wire N__9149;
    wire N__9148;
    wire N__9147;
    wire N__9146;
    wire N__9145;
    wire N__9144;
    wire N__9143;
    wire N__9142;
    wire N__9141;
    wire N__9140;
    wire N__9139;
    wire N__9136;
    wire N__9135;
    wire N__9134;
    wire N__9133;
    wire N__9132;
    wire N__9131;
    wire N__9130;
    wire N__9129;
    wire N__9128;
    wire N__9127;
    wire N__9126;
    wire N__9125;
    wire N__9124;
    wire N__9123;
    wire N__9122;
    wire N__9121;
    wire N__9120;
    wire N__9119;
    wire N__9118;
    wire N__9117;
    wire N__9034;
    wire N__9031;
    wire N__9030;
    wire N__9029;
    wire N__9028;
    wire N__9027;
    wire N__9024;
    wire N__9023;
    wire N__9022;
    wire N__9021;
    wire N__9020;
    wire N__9019;
    wire N__9018;
    wire N__9013;
    wire N__9010;
    wire N__9005;
    wire N__9002;
    wire N__8997;
    wire N__8994;
    wire N__8991;
    wire N__8988;
    wire N__8987;
    wire N__8986;
    wire N__8985;
    wire N__8984;
    wire N__8983;
    wire N__8982;
    wire N__8981;
    wire N__8980;
    wire N__8979;
    wire N__8978;
    wire N__8977;
    wire N__8976;
    wire N__8973;
    wire N__8970;
    wire N__8969;
    wire N__8968;
    wire N__8967;
    wire N__8966;
    wire N__8965;
    wire N__8962;
    wire N__8959;
    wire N__8958;
    wire N__8957;
    wire N__8956;
    wire N__8953;
    wire N__8952;
    wire N__8951;
    wire N__8948;
    wire N__8947;
    wire N__8946;
    wire N__8945;
    wire N__8944;
    wire N__8943;
    wire N__8940;
    wire N__8939;
    wire N__8938;
    wire N__8937;
    wire N__8936;
    wire N__8935;
    wire N__8934;
    wire N__8933;
    wire N__8930;
    wire N__8929;
    wire N__8842;
    wire N__8839;
    wire N__8836;
    wire N__8833;
    wire N__8830;
    wire N__8829;
    wire N__8826;
    wire N__8823;
    wire N__8820;
    wire N__8817;
    wire N__8814;
    wire N__8811;
    wire N__8808;
    wire N__8805;
    wire N__8800;
    wire N__8797;
    wire N__8796;
    wire N__8793;
    wire N__8790;
    wire N__8787;
    wire N__8784;
    wire N__8781;
    wire N__8778;
    wire N__8775;
    wire N__8772;
    wire N__8767;
    wire N__8764;
    wire N__8761;
    wire N__8758;
    wire N__8757;
    wire N__8754;
    wire N__8751;
    wire N__8746;
    wire N__8743;
    wire N__8740;
    wire N__8737;
    wire N__8734;
    wire N__8731;
    wire N__8728;
    wire N__8727;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8692;
    wire N__8689;
    wire N__8688;
    wire N__8685;
    wire N__8682;
    wire N__8679;
    wire N__8676;
    wire N__8673;
    wire N__8670;
    wire N__8667;
    wire N__8664;
    wire N__8661;
    wire N__8658;
    wire N__8653;
    wire N__8650;
    wire N__8647;
    wire N__8644;
    wire N__8641;
    wire N__8640;
    wire N__8637;
    wire N__8636;
    wire N__8635;
    wire N__8632;
    wire N__8629;
    wire N__8626;
    wire N__8623;
    wire N__8622;
    wire N__8619;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8596;
    wire N__8595;
    wire N__8592;
    wire N__8589;
    wire N__8588;
    wire N__8587;
    wire N__8586;
    wire N__8585;
    wire N__8584;
    wire N__8583;
    wire N__8580;
    wire N__8577;
    wire N__8576;
    wire N__8575;
    wire N__8572;
    wire N__8569;
    wire N__8566;
    wire N__8563;
    wire N__8562;
    wire N__8561;
    wire N__8556;
    wire N__8551;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8539;
    wire N__8538;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8524;
    wire N__8521;
    wire N__8518;
    wire N__8513;
    wire N__8510;
    wire N__8503;
    wire N__8498;
    wire N__8493;
    wire N__8490;
    wire N__8487;
    wire N__8484;
    wire N__8475;
    wire N__8472;
    wire N__8461;
    wire N__8458;
    wire N__8455;
    wire N__8452;
    wire N__8449;
    wire N__8446;
    wire N__8443;
    wire N__8442;
    wire N__8441;
    wire N__8438;
    wire N__8437;
    wire N__8436;
    wire N__8435;
    wire N__8432;
    wire N__8431;
    wire N__8430;
    wire N__8427;
    wire N__8426;
    wire N__8425;
    wire N__8420;
    wire N__8419;
    wire N__8416;
    wire N__8413;
    wire N__8410;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8398;
    wire N__8397;
    wire N__8394;
    wire N__8391;
    wire N__8386;
    wire N__8377;
    wire N__8370;
    wire N__8367;
    wire N__8364;
    wire N__8357;
    wire N__8350;
    wire N__8347;
    wire N__8344;
    wire N__8341;
    wire N__8338;
    wire N__8335;
    wire N__8332;
    wire N__8329;
    wire N__8328;
    wire N__8325;
    wire N__8322;
    wire N__8321;
    wire N__8318;
    wire N__8315;
    wire N__8312;
    wire N__8311;
    wire N__8304;
    wire N__8301;
    wire N__8296;
    wire N__8293;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8281;
    wire N__8278;
    wire N__8277;
    wire N__8274;
    wire N__8271;
    wire N__8268;
    wire N__8265;
    wire N__8262;
    wire N__8259;
    wire N__8254;
    wire N__8251;
    wire N__8248;
    wire N__8245;
    wire N__8242;
    wire N__8239;
    wire N__8236;
    wire N__8235;
    wire N__8232;
    wire N__8231;
    wire N__8230;
    wire N__8227;
    wire N__8226;
    wire N__8225;
    wire N__8224;
    wire N__8221;
    wire N__8218;
    wire N__8215;
    wire N__8212;
    wire N__8209;
    wire N__8206;
    wire N__8203;
    wire N__8198;
    wire N__8195;
    wire N__8192;
    wire N__8189;
    wire N__8184;
    wire N__8179;
    wire N__8172;
    wire N__8169;
    wire N__8166;
    wire N__8163;
    wire N__8160;
    wire N__8155;
    wire N__8152;
    wire N__8149;
    wire N__8148;
    wire N__8145;
    wire N__8142;
    wire N__8141;
    wire N__8138;
    wire N__8135;
    wire N__8132;
    wire N__8125;
    wire N__8122;
    wire N__8119;
    wire N__8116;
    wire N__8115;
    wire N__8114;
    wire N__8113;
    wire N__8112;
    wire N__8109;
    wire N__8106;
    wire N__8103;
    wire N__8100;
    wire N__8099;
    wire N__8098;
    wire N__8095;
    wire N__8090;
    wire N__8089;
    wire N__8088;
    wire N__8087;
    wire N__8086;
    wire N__8083;
    wire N__8080;
    wire N__8075;
    wire N__8072;
    wire N__8069;
    wire N__8066;
    wire N__8063;
    wire N__8060;
    wire N__8057;
    wire N__8038;
    wire N__8037;
    wire N__8036;
    wire N__8035;
    wire N__8034;
    wire N__8031;
    wire N__8028;
    wire N__8021;
    wire N__8018;
    wire N__8017;
    wire N__8016;
    wire N__8013;
    wire N__8008;
    wire N__8005;
    wire N__8002;
    wire N__7993;
    wire N__7992;
    wire N__7991;
    wire N__7990;
    wire N__7989;
    wire N__7988;
    wire N__7985;
    wire N__7982;
    wire N__7979;
    wire N__7978;
    wire N__7977;
    wire N__7976;
    wire N__7975;
    wire N__7974;
    wire N__7973;
    wire N__7970;
    wire N__7965;
    wire N__7962;
    wire N__7959;
    wire N__7956;
    wire N__7951;
    wire N__7948;
    wire N__7945;
    wire N__7940;
    wire N__7921;
    wire N__7920;
    wire N__7917;
    wire N__7916;
    wire N__7915;
    wire N__7910;
    wire N__7905;
    wire N__7900;
    wire N__7899;
    wire N__7898;
    wire N__7897;
    wire N__7894;
    wire N__7891;
    wire N__7886;
    wire N__7883;
    wire N__7876;
    wire N__7873;
    wire N__7870;
    wire N__7869;
    wire N__7866;
    wire N__7863;
    wire N__7862;
    wire N__7857;
    wire N__7854;
    wire N__7849;
    wire N__7848;
    wire N__7847;
    wire N__7846;
    wire N__7843;
    wire N__7840;
    wire N__7839;
    wire N__7838;
    wire N__7833;
    wire N__7828;
    wire N__7827;
    wire N__7824;
    wire N__7823;
    wire N__7820;
    wire N__7819;
    wire N__7814;
    wire N__7813;
    wire N__7810;
    wire N__7809;
    wire N__7808;
    wire N__7807;
    wire N__7804;
    wire N__7801;
    wire N__7796;
    wire N__7793;
    wire N__7788;
    wire N__7785;
    wire N__7780;
    wire N__7765;
    wire N__7762;
    wire N__7761;
    wire N__7758;
    wire N__7757;
    wire N__7754;
    wire N__7751;
    wire N__7748;
    wire N__7741;
    wire N__7740;
    wire N__7739;
    wire N__7736;
    wire N__7735;
    wire N__7734;
    wire N__7733;
    wire N__7732;
    wire N__7731;
    wire N__7730;
    wire N__7727;
    wire N__7726;
    wire N__7723;
    wire N__7722;
    wire N__7721;
    wire N__7720;
    wire N__7717;
    wire N__7716;
    wire N__7713;
    wire N__7710;
    wire N__7703;
    wire N__7702;
    wire N__7701;
    wire N__7700;
    wire N__7699;
    wire N__7698;
    wire N__7697;
    wire N__7696;
    wire N__7695;
    wire N__7694;
    wire N__7691;
    wire N__7688;
    wire N__7685;
    wire N__7682;
    wire N__7679;
    wire N__7674;
    wire N__7671;
    wire N__7668;
    wire N__7665;
    wire N__7662;
    wire N__7659;
    wire N__7652;
    wire N__7649;
    wire N__7644;
    wire N__7641;
    wire N__7636;
    wire N__7633;
    wire N__7600;
    wire N__7599;
    wire N__7596;
    wire N__7593;
    wire N__7590;
    wire N__7585;
    wire N__7584;
    wire N__7583;
    wire N__7582;
    wire N__7581;
    wire N__7580;
    wire N__7579;
    wire N__7576;
    wire N__7573;
    wire N__7572;
    wire N__7567;
    wire N__7564;
    wire N__7561;
    wire N__7558;
    wire N__7555;
    wire N__7552;
    wire N__7549;
    wire N__7546;
    wire N__7545;
    wire N__7538;
    wire N__7531;
    wire N__7528;
    wire N__7525;
    wire N__7520;
    wire N__7513;
    wire N__7512;
    wire N__7509;
    wire N__7506;
    wire N__7503;
    wire N__7500;
    wire N__7497;
    wire N__7496;
    wire N__7493;
    wire N__7490;
    wire N__7487;
    wire N__7486;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7468;
    wire N__7465;
    wire N__7462;
    wire N__7459;
    wire N__7456;
    wire N__7453;
    wire N__7450;
    wire N__7447;
    wire N__7444;
    wire N__7441;
    wire N__7438;
    wire N__7435;
    wire N__7432;
    wire N__7429;
    wire N__7426;
    wire N__7423;
    wire N__7420;
    wire N__7417;
    wire N__7414;
    wire N__7413;
    wire N__7412;
    wire N__7411;
    wire N__7410;
    wire N__7409;
    wire N__7408;
    wire N__7407;
    wire N__7400;
    wire N__7393;
    wire N__7390;
    wire N__7389;
    wire N__7388;
    wire N__7385;
    wire N__7384;
    wire N__7383;
    wire N__7382;
    wire N__7381;
    wire N__7378;
    wire N__7375;
    wire N__7374;
    wire N__7373;
    wire N__7372;
    wire N__7371;
    wire N__7370;
    wire N__7367;
    wire N__7362;
    wire N__7361;
    wire N__7360;
    wire N__7359;
    wire N__7358;
    wire N__7355;
    wire N__7352;
    wire N__7345;
    wire N__7342;
    wire N__7339;
    wire N__7330;
    wire N__7327;
    wire N__7322;
    wire N__7317;
    wire N__7314;
    wire N__7311;
    wire N__7288;
    wire N__7285;
    wire N__7282;
    wire N__7279;
    wire N__7276;
    wire N__7273;
    wire N__7272;
    wire N__7271;
    wire N__7268;
    wire N__7263;
    wire N__7258;
    wire N__7257;
    wire N__7254;
    wire N__7249;
    wire N__7246;
    wire N__7245;
    wire N__7244;
    wire N__7241;
    wire N__7240;
    wire N__7239;
    wire N__7238;
    wire N__7237;
    wire N__7236;
    wire N__7231;
    wire N__7228;
    wire N__7225;
    wire N__7222;
    wire N__7221;
    wire N__7218;
    wire N__7215;
    wire N__7212;
    wire N__7209;
    wire N__7204;
    wire N__7201;
    wire N__7198;
    wire N__7183;
    wire N__7180;
    wire N__7177;
    wire N__7174;
    wire N__7171;
    wire N__7168;
    wire N__7165;
    wire N__7162;
    wire N__7159;
    wire N__7156;
    wire N__7153;
    wire N__7150;
    wire N__7147;
    wire N__7144;
    wire N__7141;
    wire N__7138;
    wire N__7135;
    wire N__7132;
    wire N__7129;
    wire N__7126;
    wire N__7123;
    wire N__7120;
    wire N__7117;
    wire N__7114;
    wire N__7111;
    wire N__7108;
    wire N__7107;
    wire N__7104;
    wire N__7103;
    wire N__7102;
    wire N__7101;
    wire N__7100;
    wire N__7099;
    wire N__7096;
    wire N__7095;
    wire N__7094;
    wire N__7089;
    wire N__7084;
    wire N__7081;
    wire N__7078;
    wire N__7077;
    wire N__7076;
    wire N__7075;
    wire N__7074;
    wire N__7073;
    wire N__7070;
    wire N__7065;
    wire N__7060;
    wire N__7055;
    wire N__7052;
    wire N__7045;
    wire N__7042;
    wire N__7039;
    wire N__7028;
    wire N__7021;
    wire N__7018;
    wire N__7015;
    wire N__7012;
    wire N__7009;
    wire N__7006;
    wire N__7003;
    wire N__7000;
    wire N__6997;
    wire N__6994;
    wire N__6993;
    wire N__6990;
    wire N__6989;
    wire N__6986;
    wire N__6985;
    wire N__6982;
    wire N__6979;
    wire N__6978;
    wire N__6975;
    wire N__6972;
    wire N__6971;
    wire N__6968;
    wire N__6965;
    wire N__6962;
    wire N__6957;
    wire N__6954;
    wire N__6951;
    wire N__6948;
    wire N__6945;
    wire N__6942;
    wire N__6939;
    wire N__6928;
    wire N__6927;
    wire N__6924;
    wire N__6921;
    wire N__6918;
    wire N__6915;
    wire N__6912;
    wire N__6909;
    wire N__6906;
    wire N__6903;
    wire N__6900;
    wire N__6897;
    wire N__6894;
    wire N__6889;
    wire N__6886;
    wire N__6883;
    wire N__6880;
    wire N__6879;
    wire N__6878;
    wire N__6875;
    wire N__6874;
    wire N__6871;
    wire N__6868;
    wire N__6865;
    wire N__6862;
    wire N__6859;
    wire N__6856;
    wire N__6853;
    wire N__6850;
    wire N__6847;
    wire N__6844;
    wire N__6835;
    wire N__6832;
    wire N__6829;
    wire N__6826;
    wire N__6825;
    wire N__6824;
    wire N__6823;
    wire N__6822;
    wire N__6821;
    wire N__6820;
    wire N__6817;
    wire N__6816;
    wire N__6815;
    wire N__6814;
    wire N__6813;
    wire N__6812;
    wire N__6811;
    wire N__6810;
    wire N__6809;
    wire N__6806;
    wire N__6801;
    wire N__6798;
    wire N__6793;
    wire N__6792;
    wire N__6791;
    wire N__6790;
    wire N__6787;
    wire N__6782;
    wire N__6781;
    wire N__6780;
    wire N__6777;
    wire N__6776;
    wire N__6775;
    wire N__6774;
    wire N__6773;
    wire N__6770;
    wire N__6767;
    wire N__6764;
    wire N__6759;
    wire N__6754;
    wire N__6749;
    wire N__6748;
    wire N__6747;
    wire N__6744;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6732;
    wire N__6723;
    wire N__6720;
    wire N__6717;
    wire N__6714;
    wire N__6711;
    wire N__6706;
    wire N__6701;
    wire N__6698;
    wire N__6695;
    wire N__6692;
    wire N__6689;
    wire N__6686;
    wire N__6683;
    wire N__6676;
    wire N__6669;
    wire N__6662;
    wire N__6643;
    wire N__6640;
    wire N__6637;
    wire N__6634;
    wire N__6631;
    wire N__6630;
    wire N__6629;
    wire N__6626;
    wire N__6625;
    wire N__6624;
    wire N__6621;
    wire N__6620;
    wire N__6619;
    wire N__6616;
    wire N__6613;
    wire N__6608;
    wire N__6601;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6577;
    wire N__6574;
    wire N__6571;
    wire N__6568;
    wire N__6565;
    wire N__6562;
    wire N__6559;
    wire N__6556;
    wire N__6553;
    wire N__6550;
    wire N__6547;
    wire N__6546;
    wire N__6545;
    wire N__6542;
    wire N__6539;
    wire N__6536;
    wire N__6529;
    wire N__6528;
    wire N__6525;
    wire N__6522;
    wire N__6517;
    wire N__6514;
    wire N__6511;
    wire N__6510;
    wire N__6507;
    wire N__6504;
    wire N__6501;
    wire N__6496;
    wire N__6495;
    wire N__6494;
    wire N__6493;
    wire N__6492;
    wire N__6491;
    wire N__6488;
    wire N__6487;
    wire N__6486;
    wire N__6479;
    wire N__6478;
    wire N__6475;
    wire N__6472;
    wire N__6469;
    wire N__6464;
    wire N__6461;
    wire N__6458;
    wire N__6445;
    wire N__6442;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6430;
    wire N__6427;
    wire N__6426;
    wire N__6423;
    wire N__6420;
    wire N__6417;
    wire N__6414;
    wire N__6413;
    wire N__6410;
    wire N__6407;
    wire N__6404;
    wire N__6397;
    wire N__6394;
    wire N__6391;
    wire N__6388;
    wire N__6385;
    wire N__6382;
    wire N__6379;
    wire N__6376;
    wire N__6373;
    wire N__6370;
    wire N__6367;
    wire N__6364;
    wire N__6361;
    wire N__6358;
    wire N__6355;
    wire N__6352;
    wire N__6349;
    wire N__6346;
    wire N__6343;
    wire N__6340;
    wire N__6337;
    wire N__6334;
    wire N__6331;
    wire N__6328;
    wire N__6325;
    wire N__6322;
    wire N__6319;
    wire N__6316;
    wire N__6313;
    wire N__6310;
    wire N__6307;
    wire N__6304;
    wire N__6301;
    wire N__6298;
    wire N__6297;
    wire N__6296;
    wire N__6289;
    wire N__6286;
    wire N__6285;
    wire N__6284;
    wire N__6281;
    wire N__6278;
    wire N__6273;
    wire N__6268;
    wire N__6265;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6253;
    wire N__6250;
    wire N__6247;
    wire N__6246;
    wire N__6245;
    wire N__6242;
    wire N__6237;
    wire N__6232;
    wire N__6231;
    wire N__6228;
    wire N__6225;
    wire N__6222;
    wire N__6217;
    wire N__6214;
    wire N__6211;
    wire N__6208;
    wire N__6205;
    wire N__6202;
    wire N__6201;
    wire N__6198;
    wire N__6195;
    wire N__6190;
    wire N__6187;
    wire N__6184;
    wire N__6181;
    wire N__6180;
    wire N__6179;
    wire N__6178;
    wire N__6177;
    wire N__6174;
    wire N__6171;
    wire N__6168;
    wire N__6163;
    wire N__6160;
    wire N__6155;
    wire N__6152;
    wire N__6151;
    wire N__6148;
    wire N__6145;
    wire N__6142;
    wire N__6139;
    wire N__6130;
    wire N__6127;
    wire N__6124;
    wire N__6121;
    wire N__6118;
    wire N__6115;
    wire N__6112;
    wire N__6109;
    wire N__6106;
    wire N__6103;
    wire N__6100;
    wire N__6099;
    wire N__6096;
    wire N__6093;
    wire N__6090;
    wire N__6087;
    wire N__6082;
    wire N__6079;
    wire N__6076;
    wire N__6073;
    wire N__6070;
    wire N__6067;
    wire N__6064;
    wire N__6061;
    wire N__6058;
    wire N__6055;
    wire N__6052;
    wire N__6049;
    wire N__6046;
    wire N__6043;
    wire N__6040;
    wire N__6037;
    wire N__6034;
    wire N__6031;
    wire N__6028;
    wire N__6025;
    wire N__6022;
    wire N__6019;
    wire N__6016;
    wire N__6013;
    wire N__6010;
    wire N__6007;
    wire N__6004;
    wire N__6001;
    wire N__5998;
    wire N__5995;
    wire N__5992;
    wire N__5989;
    wire N__5986;
    wire N__5983;
    wire N__5980;
    wire N__5979;
    wire N__5976;
    wire N__5973;
    wire N__5970;
    wire N__5965;
    wire N__5962;
    wire N__5959;
    wire N__5956;
    wire N__5955;
    wire N__5952;
    wire N__5949;
    wire N__5944;
    wire N__5941;
    wire N__5940;
    wire N__5939;
    wire N__5936;
    wire N__5933;
    wire N__5930;
    wire N__5923;
    wire N__5920;
    wire N__5919;
    wire N__5916;
    wire N__5913;
    wire N__5908;
    wire N__5905;
    wire N__5902;
    wire N__5899;
    wire N__5896;
    wire N__5893;
    wire N__5890;
    wire N__5887;
    wire N__5884;
    wire N__5881;
    wire N__5878;
    wire N__5875;
    wire N__5872;
    wire N__5869;
    wire N__5866;
    wire N__5863;
    wire N__5860;
    wire N__5857;
    wire N__5854;
    wire N__5851;
    wire N__5848;
    wire N__5845;
    wire N__5842;
    wire N__5839;
    wire N__5836;
    wire N__5833;
    wire N__5830;
    wire N__5827;
    wire N__5824;
    wire N__5821;
    wire N__5818;
    wire N__5815;
    wire N__5812;
    wire N__5809;
    wire N__5806;
    wire N__5803;
    wire N__5800;
    wire N__5797;
    wire N__5794;
    wire N__5793;
    wire N__5790;
    wire N__5787;
    wire N__5782;
    wire N__5779;
    wire N__5776;
    wire N__5775;
    wire N__5772;
    wire N__5771;
    wire N__5768;
    wire N__5765;
    wire N__5762;
    wire N__5755;
    wire N__5752;
    wire N__5749;
    wire N__5748;
    wire N__5745;
    wire N__5742;
    wire N__5737;
    wire N__5734;
    wire N__5731;
    wire N__5728;
    wire N__5725;
    wire N__5722;
    wire N__5719;
    wire N__5716;
    wire N__5713;
    wire N__5710;
    wire N__5707;
    wire N__5704;
    wire N__5701;
    wire N__5698;
    wire N__5695;
    wire N__5692;
    wire N__5689;
    wire N__5686;
    wire N__5685;
    wire N__5680;
    wire N__5677;
    wire N__5676;
    wire N__5675;
    wire N__5672;
    wire N__5667;
    wire N__5662;
    wire N__5659;
    wire N__5656;
    wire N__5653;
    wire N__5650;
    wire N__5647;
    wire N__5644;
    wire N__5641;
    wire N__5638;
    wire N__5635;
    wire N__5632;
    wire N__5629;
    wire N__5626;
    wire N__5623;
    wire N__5622;
    wire N__5619;
    wire N__5616;
    wire N__5611;
    wire N__5608;
    wire N__5605;
    wire N__5602;
    wire N__5599;
    wire N__5596;
    wire N__5593;
    wire N__5590;
    wire N__5587;
    wire N__5584;
    wire N__5581;
    wire N__5580;
    wire N__5577;
    wire N__5574;
    wire N__5571;
    wire N__5568;
    wire N__5565;
    wire N__5562;
    wire N__5557;
    wire N__5554;
    wire N__5551;
    wire N__5548;
    wire N__5545;
    wire N__5542;
    wire N__5539;
    wire N__5536;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5518;
    wire N__5515;
    wire N__5512;
    wire N__5509;
    wire N__5506;
    wire N__5503;
    wire N__5500;
    wire N__5497;
    wire N__5494;
    wire N__5491;
    wire N__5488;
    wire N__5485;
    wire N__5482;
    wire N__5479;
    wire N__5476;
    wire N__5473;
    wire N__5470;
    wire N__5467;
    wire N__5464;
    wire N__5461;
    wire N__5458;
    wire N__5455;
    wire N__5452;
    wire N__5449;
    wire N__5446;
    wire N__5443;
    wire N__5440;
    wire N__5437;
    wire N__5434;
    wire N__5431;
    wire N__5428;
    wire N__5425;
    wire N__5422;
    wire N__5419;
    wire N__5416;
    wire N__5413;
    wire N__5410;
    wire N__5407;
    wire N__5404;
    wire N__5401;
    wire N__5398;
    wire N__5395;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5332;
    wire N__5329;
    wire N__5326;
    wire N__5323;
    wire N__5320;
    wire N__5317;
    wire N__5314;
    wire N__5311;
    wire N__5308;
    wire N__5305;
    wire N__5302;
    wire N__5299;
    wire N__5296;
    wire N__5293;
    wire N__5290;
    wire N__5287;
    wire N__5284;
    wire N__5281;
    wire N__5278;
    wire N__5275;
    wire N__5272;
    wire N__5269;
    wire N__5266;
    wire N__5263;
    wire N__5260;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5248;
    wire N__5247;
    wire N__5246;
    wire N__5243;
    wire N__5240;
    wire N__5237;
    wire N__5234;
    wire N__5229;
    wire N__5226;
    wire N__5223;
    wire N__5220;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5208;
    wire N__5203;
    wire N__5202;
    wire N__5199;
    wire N__5198;
    wire N__5191;
    wire N__5188;
    wire N__5185;
    wire N__5182;
    wire N__5179;
    wire N__5176;
    wire N__5173;
    wire N__5170;
    wire N__5167;
    wire N__5166;
    wire N__5163;
    wire N__5160;
    wire N__5157;
    wire N__5154;
    wire N__5151;
    wire N__5148;
    wire N__5143;
    wire N__5140;
    wire N__5139;
    wire N__5136;
    wire N__5133;
    wire N__5130;
    wire N__5127;
    wire N__5124;
    wire N__5121;
    wire N__5116;
    wire N__5113;
    wire N__5110;
    wire N__5107;
    wire N__5106;
    wire N__5103;
    wire N__5100;
    wire N__5095;
    wire N__5094;
    wire N__5091;
    wire N__5088;
    wire N__5087;
    wire N__5084;
    wire N__5081;
    wire N__5078;
    wire N__5071;
    wire N__5070;
    wire N__5065;
    wire N__5064;
    wire N__5061;
    wire N__5060;
    wire N__5057;
    wire N__5054;
    wire N__5051;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5035;
    wire N__5032;
    wire N__5029;
    wire N__5026;
    wire N__5023;
    wire N__5020;
    wire N__5017;
    wire N__5014;
    wire N__5011;
    wire N__5008;
    wire N__5005;
    wire N__5002;
    wire N__4999;
    wire N__4996;
    wire N__4993;
    wire N__4990;
    wire N__4987;
    wire N__4984;
    wire N__4981;
    wire N__4978;
    wire N__4975;
    wire N__4972;
    wire N__4971;
    wire N__4968;
    wire N__4965;
    wire N__4962;
    wire N__4959;
    wire N__4954;
    wire N__4951;
    wire N__4948;
    wire N__4945;
    wire N__4942;
    wire N__4939;
    wire N__4936;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4924;
    wire N__4921;
    wire N__4918;
    wire N__4915;
    wire N__4912;
    wire N__4909;
    wire N__4908;
    wire N__4905;
    wire N__4902;
    wire N__4897;
    wire N__4896;
    wire N__4893;
    wire N__4890;
    wire N__4885;
    wire N__4884;
    wire N__4881;
    wire N__4878;
    wire N__4875;
    wire N__4870;
    wire N__4869;
    wire N__4866;
    wire N__4863;
    wire N__4858;
    wire N__4857;
    wire N__4854;
    wire N__4851;
    wire N__4846;
    wire N__4845;
    wire N__4842;
    wire N__4839;
    wire N__4834;
    wire N__4831;
    wire N__4828;
    wire N__4825;
    wire N__4824;
    wire N__4821;
    wire N__4818;
    wire N__4815;
    wire N__4812;
    wire N__4807;
    wire N__4804;
    wire N__4803;
    wire N__4800;
    wire N__4797;
    wire N__4792;
    wire N__4789;
    wire N__4786;
    wire N__4783;
    wire N__4780;
    wire N__4777;
    wire N__4774;
    wire N__4771;
    wire N__4770;
    wire N__4767;
    wire N__4764;
    wire N__4761;
    wire N__4758;
    wire N__4753;
    wire N__4750;
    wire N__4747;
    wire N__4744;
    wire N__4741;
    wire N__4738;
    wire N__4735;
    wire N__4732;
    wire N__4731;
    wire N__4728;
    wire N__4725;
    wire N__4720;
    wire N__4717;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4705;
    wire N__4702;
    wire N__4699;
    wire N__4696;
    wire N__4693;
    wire N__4690;
    wire N__4689;
    wire N__4686;
    wire N__4683;
    wire N__4678;
    wire N__4675;
    wire N__4674;
    wire N__4673;
    wire N__4672;
    wire N__4669;
    wire N__4666;
    wire N__4661;
    wire N__4658;
    wire N__4651;
    wire N__4650;
    wire N__4649;
    wire N__4646;
    wire N__4641;
    wire N__4636;
    wire N__4633;
    wire N__4632;
    wire N__4629;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4612;
    wire N__4611;
    wire N__4608;
    wire N__4605;
    wire N__4602;
    wire N__4599;
    wire N__4594;
    wire N__4591;
    wire N__4588;
    wire N__4585;
    wire N__4582;
    wire N__4579;
    wire N__4578;
    wire N__4577;
    wire N__4576;
    wire N__4567;
    wire N__4564;
    wire N__4563;
    wire N__4560;
    wire N__4559;
    wire N__4554;
    wire N__4551;
    wire N__4546;
    wire N__4545;
    wire N__4542;
    wire N__4539;
    wire N__4534;
    wire N__4531;
    wire N__4528;
    wire N__4525;
    wire N__4522;
    wire N__4519;
    wire N__4516;
    wire N__4513;
    wire N__4510;
    wire N__4507;
    wire N__4504;
    wire N__4501;
    wire N__4498;
    wire N__4495;
    wire N__4492;
    wire N__4489;
    wire N__4486;
    wire N__4483;
    wire N__4480;
    wire N__4477;
    wire N__4474;
    wire N__4471;
    wire N__4468;
    wire N__4465;
    wire N__4462;
    wire N__4461;
    wire N__4460;
    wire N__4459;
    wire N__4456;
    wire N__4453;
    wire N__4448;
    wire N__4441;
    wire N__4440;
    wire N__4437;
    wire N__4436;
    wire N__4435;
    wire N__4434;
    wire N__4431;
    wire N__4428;
    wire N__4425;
    wire N__4420;
    wire N__4411;
    wire N__4410;
    wire N__4407;
    wire N__4404;
    wire N__4399;
    wire N__4396;
    wire N__4395;
    wire N__4392;
    wire N__4389;
    wire N__4384;
    wire N__4383;
    wire N__4382;
    wire N__4381;
    wire N__4380;
    wire N__4379;
    wire N__4378;
    wire N__4375;
    wire N__4368;
    wire N__4361;
    wire N__4354;
    wire N__4351;
    wire N__4350;
    wire N__4349;
    wire N__4348;
    wire N__4347;
    wire N__4346;
    wire N__4341;
    wire N__4340;
    wire N__4339;
    wire N__4336;
    wire N__4331;
    wire N__4328;
    wire N__4325;
    wire N__4320;
    wire N__4309;
    wire N__4308;
    wire N__4303;
    wire N__4300;
    wire N__4299;
    wire N__4296;
    wire N__4295;
    wire N__4294;
    wire N__4293;
    wire N__4288;
    wire N__4281;
    wire N__4276;
    wire N__4273;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4261;
    wire N__4258;
    wire N__4255;
    wire N__4252;
    wire N__4249;
    wire N__4246;
    wire N__4243;
    wire N__4240;
    wire N__4237;
    wire N__4236;
    wire N__4233;
    wire N__4230;
    wire N__4225;
    wire N__4222;
    wire N__4221;
    wire N__4220;
    wire N__4219;
    wire N__4216;
    wire N__4209;
    wire N__4204;
    wire N__4201;
    wire N__4198;
    wire N__4195;
    wire N__4192;
    wire N__4189;
    wire N__4186;
    wire N__4183;
    wire N__4180;
    wire N__4177;
    wire N__4174;
    wire N__4171;
    wire N__4168;
    wire N__4165;
    wire N__4162;
    wire N__4161;
    wire N__4160;
    wire N__4153;
    wire N__4150;
    wire N__4149;
    wire N__4148;
    wire N__4147;
    wire N__4140;
    wire N__4137;
    wire N__4132;
    wire N__4129;
    wire N__4126;
    wire N__4123;
    wire N__4120;
    wire N__4117;
    wire N__4116;
    wire N__4111;
    wire N__4108;
    wire N__4105;
    wire N__4102;
    wire N__4099;
    wire N__4096;
    wire N__4093;
    wire N__4090;
    wire N__4087;
    wire N__4084;
    wire N__4083;
    wire N__4080;
    wire N__4077;
    wire N__4072;
    wire N__4071;
    wire N__4068;
    wire N__4067;
    wire N__4060;
    wire N__4057;
    wire N__4056;
    wire N__4055;
    wire N__4048;
    wire N__4045;
    wire N__4044;
    wire N__4043;
    wire N__4040;
    wire N__4037;
    wire N__4034;
    wire N__4027;
    wire N__4024;
    wire N__4021;
    wire N__4020;
    wire N__4019;
    wire N__4014;
    wire N__4011;
    wire N__4006;
    wire N__4003;
    wire N__4002;
    wire N__3999;
    wire N__3996;
    wire N__3991;
    wire N__3988;
    wire N__3985;
    wire N__3982;
    wire N__3979;
    wire N__3976;
    wire N__3973;
    wire N__3972;
    wire N__3969;
    wire N__3966;
    wire N__3963;
    wire N__3960;
    wire N__3957;
    wire N__3952;
    wire N__3949;
    wire N__3946;
    wire N__3945;
    wire N__3944;
    wire N__3943;
    wire N__3940;
    wire N__3933;
    wire N__3928;
    wire N__3927;
    wire N__3924;
    wire N__3921;
    wire N__3916;
    wire N__3913;
    wire N__3910;
    wire N__3907;
    wire N__3904;
    wire N__3901;
    wire N__3898;
    wire N__3895;
    wire N__3892;
    wire N__3891;
    wire N__3886;
    wire N__3883;
    wire N__3882;
    wire N__3877;
    wire N__3874;
    wire N__3873;
    wire N__3870;
    wire N__3867;
    wire N__3864;
    wire N__3861;
    wire N__3858;
    wire N__3855;
    wire N__3852;
    wire N__3849;
    wire N__3846;
    wire N__3843;
    wire N__3842;
    wire N__3839;
    wire N__3836;
    wire N__3833;
    wire N__3828;
    wire N__3825;
    wire N__3820;
    wire N__3819;
    wire N__3818;
    wire N__3815;
    wire N__3810;
    wire N__3805;
    wire N__3802;
    wire N__3801;
    wire N__3800;
    wire N__3795;
    wire N__3792;
    wire N__3787;
    wire N__3784;
    wire N__3781;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire N__3773;
    wire N__3772;
    wire N__3769;
    wire N__3766;
    wire N__3761;
    wire N__3754;
    wire N__3753;
    wire N__3748;
    wire N__3745;
    wire N__3742;
    wire N__3739;
    wire N__3738;
    wire N__3735;
    wire N__3732;
    wire N__3727;
    wire N__3724;
    wire N__3721;
    wire N__3718;
    wire N__3715;
    wire N__3712;
    wire N__3709;
    wire N__3706;
    wire N__3703;
    wire N__3700;
    wire N__3697;
    wire N__3694;
    wire N__3693;
    wire N__3690;
    wire N__3687;
    wire N__3682;
    wire N__3681;
    wire N__3680;
    wire N__3677;
    wire N__3672;
    wire N__3669;
    wire N__3666;
    wire N__3661;
    wire N__3658;
    wire N__3655;
    wire N__3654;
    wire N__3651;
    wire N__3648;
    wire N__3643;
    wire N__3640;
    wire N__3637;
    wire N__3634;
    wire N__3631;
    wire N__3628;
    wire N__3625;
    wire N__3622;
    wire N__3619;
    wire N__3616;
    wire N__3613;
    wire N__3610;
    wire N__3607;
    wire N__3604;
    wire N__3601;
    wire N__3598;
    wire N__3595;
    wire N__3592;
    wire N__3589;
    wire N__3586;
    wire N__3583;
    wire N__3582;
    wire N__3579;
    wire N__3574;
    wire N__3571;
    wire N__3568;
    wire N__3565;
    wire N__3562;
    wire N__3559;
    wire N__3556;
    wire N__3553;
    wire N__3550;
    wire N__3547;
    wire N__3544;
    wire N__3541;
    wire N__3538;
    wire N__3535;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire CLK80_OUT_i_i;
    wire CLK40_OUT_i_i;
    wire \U712_REG_SM.LDS_OUT_2_0_a2Z0Z_0 ;
    wire VBENn_c;
    wire SIZ_c_0;
    wire \U712_BYTE_ENABLE.N_387_cascade_ ;
    wire N_73_i;
    wire A_c_0;
    wire SIZ_c_1;
    wire REGSPACEn_c;
    wire \U712_REG_SM.N_301 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_0 ;
    wire ASn_c;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_2 ;
    wire \U712_REG_SM.N_281_cascade_ ;
    wire \U712_REG_SM.N_280_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_1 ;
    wire \U712_REG_SM.N_308 ;
    wire \U712_REG_SM.N_288_cascade_ ;
    wire \U712_REG_SM.N_307 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_2 ;
    wire C3_c;
    wire C1_c;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2Z0Z_0 ;
    wire N_75_i;
    wire \U712_BYTE_ENABLE.N_395 ;
    wire N_74_i;
    wire \U712_BYTE_ENABLE.N_387 ;
    wire A_c_1;
    wire \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_0_0 ;
    wire N_76_i;
    wire \U712_BYTE_ENABLE.N_391 ;
    wire \U712_REG_SM.N_304 ;
    wire \U712_REG_SM.N_299 ;
    wire \U712_REG_SM.N_281 ;
    wire \U712_REG_SM.N_280 ;
    wire \U712_REG_SM.N_373_cascade_ ;
    wire \U712_REG_SM.C3_SYNCZ0Z_2 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.N_289 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_6 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire \U712_REG_SM.N_289_cascade_ ;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_REG_SM.N_494 ;
    wire \U712_REG_SM.N_288 ;
    wire \U712_REG_SM.N_494_cascade_ ;
    wire \U712_REG_SM.N_424 ;
    wire \U712_REG_SM.N_369 ;
    wire \U712_REG_SM.DS_EN_RNOZ0Z_2_cascade_ ;
    wire \U712_REG_SM.N_123 ;
    wire TACK_OUTn;
    wire CLK40_OUT_i;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_2 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ;
    wire N_886_i;
    wire A_c_4;
    wire \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_2_cascade_ ;
    wire A_c_11;
    wire bfn_11_9_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire C1_c_g;
    wire \U712_REG_SM.N_306 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_5 ;
    wire \U712_REG_SM.N_298 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire \U712_REG_SM.UDS_OUTZ0 ;
    wire U712_REG_SM_un1_UDSn_i;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.N_305_i_0_en_cascade_ ;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire DRA_c_1;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.N_341_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_1_1_cascade_ ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_0_cascade_ ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ;
    wire \U712_BYTE_ENABLE.N_392 ;
    wire \U712_BYTE_ENABLE.N_388 ;
    wire CASLn_c;
    wire CASUn_c;
    wire RAMENn_c;
    wire TSn_c;
    wire REG_TACK;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire TACK_EN_i_ess;
    wire \U712_CYCLE_TERM.N_305_i_0_en_0 ;
    wire RESETn_c_i;
    wire A_c_7;
    wire A_c_14;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire A_c_9;
    wire A_c_2;
    wire \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_0_cascade_ ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire A_c_10;
    wire A_c_3;
    wire \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_1_cascade_ ;
    wire CMA_c_10;
    wire \U712_CHIP_RAM.N_313 ;
    wire CMA_c_2;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire A_c_5;
    wire \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_3_cascade_ ;
    wire A_c_12;
    wire \U712_CHIP_RAM.N_314_cascade_ ;
    wire CMA_c_3;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_5 ;
    wire DRA_c_6;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire A_c_8;
    wire \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_6_cascade_ ;
    wire A_c_15;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire DBRn_c;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_2_cascade_ ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire U712_REG_SM_DBR_SYNC_0;
    wire U712_REG_SM_DBR_SYNC_1;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_3_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_2_1_cascade_ ;
    wire \U712_CHIP_RAM.N_421_cascade_ ;
    wire \U712_CHIP_RAM.N_293_cascade_ ;
    wire \U712_CHIP_RAM.N_309_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0_a2_0_a2_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0 ;
    wire CPU_TACKm;
    wire \U712_REG_SM.DS_ENZ0 ;
    wire \U712_REG_SM.LDS_OUTZ0 ;
    wire U712_REG_SM_un1_LDSn_i;
    wire \U712_CHIP_RAM.N_311 ;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.N_312 ;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.N_316 ;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.un1_CMA31_0_i_cascade_ ;
    wire A_c_6;
    wire \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_4 ;
    wire A_c_13;
    wire \U712_CHIP_RAM.N_493_cascade_ ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_cascade_ ;
    wire \U712_CHIP_RAM.N_317 ;
    wire CMA_c_6;
    wire A_c_19;
    wire \U712_CHIP_RAM.CMA_5_i_0_8_cascade_ ;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_cascade_ ;
    wire \U712_CHIP_RAM.N_285 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_7_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0 ;
    wire DBENn_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_0_a2_0_0 ;
    wire \U712_CHIP_RAM.N_427 ;
    wire \U712_CHIP_RAM.N_421 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_ ;
    wire \U712_CHIP_RAM.N_296 ;
    wire \U712_CHIP_RAM.N_296_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_a2_0_0_0 ;
    wire \U712_CHIP_RAM.N_403 ;
    wire \U712_CHIP_RAM.N_309 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0 ;
    wire \U712_CHIP_RAM.REFRESH_CYCLEZ0 ;
    wire \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER46_cascade_ ;
    wire \U712_CHIP_RAM.N_420 ;
    wire \U712_CHIP_RAM.N_282 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_a5_i_0_cascade_ ;
    wire \U712_CHIP_RAM.N_49 ;
    wire DBDIR_c;
    wire N_218;
    wire RASn_c;
    wire A_c_18;
    wire \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_7_cascade_ ;
    wire A_c_16;
    wire A_c_17;
    wire \U712_CHIP_RAM.CMA_5_i_0_8 ;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.N_318 ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire \U712_CHIP_RAM.N_315 ;
    wire CMA_c_4;
    wire \U712_CHIP_RAM.un1_CMA31_0_i_0 ;
    wire AWEn_c;
    wire RnW_c;
    wire CPU_CYCLEm;
    wire \U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_0 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_i_a2_1_0_a2_1_0 ;
    wire \U712_CHIP_RAM.N_284 ;
    wire \U712_CHIP_RAM.N_284_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_1_2 ;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_1_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c6_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_0_3 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.N_274 ;
    wire RESETn_c;
    wire \U712_CHIP_RAM.N_274_cascade_ ;
    wire \U712_CHIP_RAM.N_337 ;
    wire \U712_CHIP_RAM.N_337_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_2_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.N_271 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER46 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.N_303 ;
    wire DMA_CYCLEm;
    wire REG_CYCLEm;
    wire DRDENn_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire CASn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire WEn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CRCSn_c;
    wire RAS0n_c;
    wire RAS1n_c;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_1 ;
    wire CLK80_OUT;
    wire RESETn_c_i_g;
    wire CONSTANT_ONE_NET;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_OUT_i),
            .REFERENCECLK(N__3553),
            .RESETB(N__8836),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_OUT),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__9911),
            .DIN(N__9910),
            .DOUT(N__9909),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__9911),
            .PADOUT(N__9910),
            .PADIN(N__9909),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6190),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__9902),
            .DIN(N__9901),
            .DOUT(N__9900),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__9902),
            .PADOUT(N__9901),
            .PADIN(N__9900),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__9893),
            .DIN(N__9892),
            .DOUT(N__9891),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__9893),
            .PADOUT(N__9892),
            .PADIN(N__9891),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8461),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__9884),
            .DIN(N__9883),
            .DOUT(N__9882),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__9884),
            .PADOUT(N__9883),
            .PADIN(N__9882),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6397),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__9875),
            .DIN(N__9874),
            .DOUT(N__9873),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__9875),
            .PADOUT(N__9874),
            .PADIN(N__9873),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__9866),
            .DIN(N__9865),
            .DOUT(N__9864),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__9866),
            .PADOUT(N__9865),
            .PADIN(N__9864),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__9857),
            .DIN(N__9856),
            .DOUT(N__9855),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__9857),
            .PADOUT(N__9856),
            .PADIN(N__9855),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__9848),
            .DIN(N__9847),
            .DOUT(N__9846),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__9848),
            .PADOUT(N__9847),
            .PADIN(N__9846),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS1n_ibuf_iopad (
            .OE(N__9839),
            .DIN(N__9838),
            .DOUT(N__9837),
            .PACKAGEPIN(RAS1n));
    defparam RAS1n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS1n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS1n_ibuf_preio (
            .PADOEN(N__9839),
            .PADOUT(N__9838),
            .PADIN(N__9837),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS1n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__9830),
            .DIN(N__9829),
            .DOUT(N__9828),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__9830),
            .PADOUT(N__9829),
            .PADIN(N__9828),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__9821),
            .DIN(N__9820),
            .DOUT(N__9819),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__9821),
            .PADOUT(N__9820),
            .PADIN(N__9819),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7129),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuf_iopad (
            .OE(N__9812),
            .DIN(N__9811),
            .DOUT(N__9810),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMENn_obuf_preio (
            .PADOEN(N__9812),
            .PADOUT(N__9811),
            .PADIN(N__9810),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5166),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__9803),
            .DIN(N__9802),
            .DOUT(N__9801),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__9803),
            .PADOUT(N__9802),
            .PADIN(N__9801),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__9794),
            .DIN(N__9793),
            .DOUT(N__9792),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__9794),
            .PADOUT(N__9793),
            .PADIN(N__9792),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__9785),
            .DIN(N__9784),
            .DOUT(N__9783),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__9785),
            .PADOUT(N__9784),
            .PADIN(N__9783),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3571),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__9776),
            .DIN(N__9775),
            .DOUT(N__9774),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__9776),
            .PADOUT(N__9775),
            .PADIN(N__9774),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__9767),
            .DIN(N__9766),
            .DOUT(N__9765),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__9767),
            .PADOUT(N__9766),
            .PADIN(N__9765),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__9758),
            .DIN(N__9757),
            .DOUT(N__9756),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__9758),
            .PADOUT(N__9757),
            .PADIN(N__9756),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5881),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__9749),
            .DIN(N__9748),
            .DOUT(N__9747),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__9749),
            .PADOUT(N__9748),
            .PADIN(N__9747),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__9740),
            .DIN(N__9739),
            .DOUT(N__9738),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__9740),
            .PADOUT(N__9739),
            .PADIN(N__9738),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8296),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__9731),
            .DIN(N__9730),
            .DOUT(N__9729),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__9731),
            .PADOUT(N__9730),
            .PADIN(N__9729),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__9722),
            .DIN(N__9721),
            .DOUT(N__9720),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__9722),
            .PADOUT(N__9721),
            .PADIN(N__9720),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__9713),
            .DIN(N__9712),
            .DOUT(N__9711),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__9713),
            .PADOUT(N__9712),
            .PADIN(N__9711),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__9704),
            .DIN(N__9703),
            .DOUT(N__9702),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__9704),
            .PADOUT(N__9703),
            .PADIN(N__9702),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__9695),
            .DIN(N__9694),
            .DOUT(N__9693),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__9695),
            .PADOUT(N__9694),
            .PADIN(N__9693),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__9686),
            .DIN(N__9685),
            .DOUT(N__9684),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__9686),
            .PADOUT(N__9685),
            .PADIN(N__9684),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8829),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__9677),
            .DIN(N__9676),
            .DOUT(N__9675),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__9677),
            .PADOUT(N__9676),
            .PADIN(N__9675),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__9668),
            .DIN(N__9667),
            .DOUT(N__9666),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__9668),
            .PADOUT(N__9667),
            .PADIN(N__9666),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__9659),
            .DIN(N__9658),
            .DOUT(N__9657),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__9659),
            .PADOUT(N__9658),
            .PADIN(N__9657),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__9650),
            .DIN(N__9649),
            .DOUT(N__9648),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__9650),
            .PADOUT(N__9649),
            .PADIN(N__9648),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__9641),
            .DIN(N__9640),
            .DOUT(N__9639),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__9641),
            .PADOUT(N__9640),
            .PADIN(N__9639),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__9632),
            .DIN(N__9631),
            .DOUT(N__9630),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__9632),
            .PADOUT(N__9631),
            .PADIN(N__9630),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6043),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__9623),
            .DIN(N__9622),
            .DOUT(N__9621),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__9623),
            .PADOUT(N__9622),
            .PADIN(N__9621),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__9614),
            .DIN(N__9613),
            .DOUT(N__9612),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__9614),
            .PADOUT(N__9613),
            .PADIN(N__9612),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__9605),
            .DIN(N__9604),
            .DOUT(N__9603),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__9605),
            .PADOUT(N__9604),
            .PADIN(N__9603),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__9596),
            .DIN(N__9595),
            .DOUT(N__9594),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__9596),
            .PADOUT(N__9595),
            .PADIN(N__9594),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_obuf_iopad (
            .OE(N__9587),
            .DIN(N__9586),
            .DOUT(N__9585),
            .PACKAGEPIN(CLK40C));
    defparam CLK40C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_obuf_preio (
            .PADOEN(N__9587),
            .PADOUT(N__9586),
            .PADIN(N__9585),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3595),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__9578),
            .DIN(N__9577),
            .DOUT(N__9576),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__9578),
            .PADOUT(N__9577),
            .PADIN(N__9576),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5908),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__9569),
            .DIN(N__9568),
            .DOUT(N__9567),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__9569),
            .PADOUT(N__9568),
            .PADIN(N__9567),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__9560),
            .DIN(N__9559),
            .DOUT(N__9558),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__9560),
            .PADOUT(N__9559),
            .PADIN(N__9558),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6382),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__9551),
            .DIN(N__9550),
            .DOUT(N__9549),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__9551),
            .PADOUT(N__9550),
            .PADIN(N__9549),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__9542),
            .DIN(N__9541),
            .DOUT(N__9540),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__9542),
            .PADOUT(N__9541),
            .PADIN(N__9540),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__9533),
            .DIN(N__9532),
            .DOUT(N__9531),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__9533),
            .PADOUT(N__9532),
            .PADIN(N__9531),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3610),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__9524),
            .DIN(N__9523),
            .DOUT(N__9522),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__9524),
            .PADOUT(N__9523),
            .PADIN(N__9522),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__9515),
            .DIN(N__9514),
            .DOUT(N__9513),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__9515),
            .PADOUT(N__9514),
            .PADIN(N__9513),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3874),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__9506),
            .DIN(N__9505),
            .DOUT(N__9504),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__9506),
            .PADOUT(N__9505),
            .PADIN(N__9504),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5659),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__9497),
            .DIN(N__9496),
            .DOUT(N__9495),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__9497),
            .PADOUT(N__9496),
            .PADIN(N__9495),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__9488),
            .DIN(N__9487),
            .DOUT(N__9486),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__9488),
            .PADOUT(N__9487),
            .PADIN(N__9486),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_0_iopad (
            .OE(N__9479),
            .DIN(N__9478),
            .DOUT(N__9477),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__9479),
            .PADOUT(N__9478),
            .PADIN(N__9477),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__9470),
            .DIN(N__9469),
            .DOUT(N__9468),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__9470),
            .PADOUT(N__9469),
            .PADIN(N__9468),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5371),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__9461),
            .DIN(N__9460),
            .DOUT(N__9459),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__9461),
            .PADOUT(N__9460),
            .PADIN(N__9459),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__9452),
            .DIN(N__9451),
            .DOUT(N__9450),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__9452),
            .PADOUT(N__9451),
            .PADIN(N__9450),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7012),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__9443),
            .DIN(N__9442),
            .DOUT(N__9441),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__9443),
            .PADOUT(N__9442),
            .PADIN(N__9441),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7468),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__9434),
            .DIN(N__9433),
            .DOUT(N__9432),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__9434),
            .PADOUT(N__9433),
            .PADIN(N__9432),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3715),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__9425),
            .DIN(N__9424),
            .DOUT(N__9423),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__9425),
            .PADOUT(N__9424),
            .PADIN(N__9423),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6004),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__9416),
            .DIN(N__9415),
            .DOUT(N__9414),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__9416),
            .PADOUT(N__9415),
            .PADIN(N__9414),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3873),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__9407),
            .DIN(N__9406),
            .DOUT(N__9405),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__9407),
            .PADOUT(N__9406),
            .PADIN(N__9405),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__9398),
            .DIN(N__9397),
            .DOUT(N__9396),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__9398),
            .PADOUT(N__9397),
            .PADIN(N__9396),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__9389),
            .DIN(N__9388),
            .DOUT(N__9387),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__9389),
            .PADOUT(N__9388),
            .PADIN(N__9387),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4186),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__9380),
            .DIN(N__9379),
            .DOUT(N__9378),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__9380),
            .PADOUT(N__9379),
            .PADIN(N__9378),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8350),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__9371),
            .DIN(N__9370),
            .DOUT(N__9369),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__9371),
            .PADOUT(N__9370),
            .PADIN(N__9369),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6436),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__9362),
            .DIN(N__9361),
            .DOUT(N__9360),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__9362),
            .PADOUT(N__9361),
            .PADIN(N__9360),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3916),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__9353),
            .DIN(N__9352),
            .DOUT(N__9351),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__9353),
            .PADOUT(N__9352),
            .PADIN(N__9351),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__9344),
            .DIN(N__9343),
            .DOUT(N__9342),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__9344),
            .PADOUT(N__9343),
            .PADIN(N__9342),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__9335),
            .DIN(N__9334),
            .DOUT(N__9333),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__9335),
            .PADOUT(N__9334),
            .PADIN(N__9333),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__9326),
            .DIN(N__9325),
            .DOUT(N__9324),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__9326),
            .PADOUT(N__9325),
            .PADIN(N__9324),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__9317),
            .DIN(N__9316),
            .DOUT(N__9315),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__9317),
            .PADOUT(N__9316),
            .PADIN(N__9315),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5857),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__9308),
            .DIN(N__9307),
            .DOUT(N__9306),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__9308),
            .PADOUT(N__9307),
            .PADIN(N__9306),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__9299),
            .DIN(N__9298),
            .DOUT(N__9297),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__9299),
            .PADOUT(N__9298),
            .PADIN(N__9297),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4108),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__9290),
            .DIN(N__9289),
            .DOUT(N__9288),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__9290),
            .PADOUT(N__9289),
            .PADIN(N__9288),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4528),
            .DIN0(),
            .DOUT0(N__4246),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__9281),
            .DIN(N__9280),
            .DOUT(N__9279),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__9281),
            .PADOUT(N__9280),
            .PADIN(N__9279),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5341),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__9272),
            .DIN(N__9271),
            .DOUT(N__9270),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__9272),
            .PADOUT(N__9271),
            .PADIN(N__9270),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__9263),
            .DIN(N__9262),
            .DOUT(N__9261),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__9263),
            .PADOUT(N__9262),
            .PADIN(N__9261),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__9254),
            .DIN(N__9253),
            .DOUT(N__9252),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__9254),
            .PADOUT(N__9253),
            .PADIN(N__9252),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7156),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__9245),
            .DIN(N__9244),
            .DOUT(N__9243),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__9245),
            .PADOUT(N__9244),
            .PADIN(N__9243),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__9236),
            .DIN(N__9235),
            .DOUT(N__9234),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__9236),
            .PADOUT(N__9235),
            .PADIN(N__9234),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__9227),
            .DIN(N__9226),
            .DOUT(N__9225),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__9227),
            .PADOUT(N__9226),
            .PADIN(N__9225),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__9218),
            .DIN(N__9217),
            .DOUT(N__9216),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__9218),
            .PADOUT(N__9217),
            .PADIN(N__9216),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__9209),
            .DIN(N__9208),
            .DOUT(N__9207),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__9209),
            .PADOUT(N__9208),
            .PADIN(N__9207),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5833),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__9200),
            .DIN(N__9199),
            .DOUT(N__9198),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__9200),
            .PADOUT(N__9199),
            .PADIN(N__9198),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4594),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2181 (
            .O(N__9181),
            .I(N__9177));
    InMux I__2180 (
            .O(N__9180),
            .I(N__9174));
    LocalMux I__2179 (
            .O(N__9177),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    LocalMux I__2178 (
            .O(N__9174),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    InMux I__2177 (
            .O(N__9169),
            .I(N__9166));
    LocalMux I__2176 (
            .O(N__9166),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ));
    InMux I__2175 (
            .O(N__9163),
            .I(N__9160));
    LocalMux I__2174 (
            .O(N__9160),
            .I(N__9136));
    ClkMux I__2173 (
            .O(N__9159),
            .I(N__9034));
    ClkMux I__2172 (
            .O(N__9158),
            .I(N__9034));
    ClkMux I__2171 (
            .O(N__9157),
            .I(N__9034));
    ClkMux I__2170 (
            .O(N__9156),
            .I(N__9034));
    ClkMux I__2169 (
            .O(N__9155),
            .I(N__9034));
    ClkMux I__2168 (
            .O(N__9154),
            .I(N__9034));
    ClkMux I__2167 (
            .O(N__9153),
            .I(N__9034));
    ClkMux I__2166 (
            .O(N__9152),
            .I(N__9034));
    ClkMux I__2165 (
            .O(N__9151),
            .I(N__9034));
    ClkMux I__2164 (
            .O(N__9150),
            .I(N__9034));
    ClkMux I__2163 (
            .O(N__9149),
            .I(N__9034));
    ClkMux I__2162 (
            .O(N__9148),
            .I(N__9034));
    ClkMux I__2161 (
            .O(N__9147),
            .I(N__9034));
    ClkMux I__2160 (
            .O(N__9146),
            .I(N__9034));
    ClkMux I__2159 (
            .O(N__9145),
            .I(N__9034));
    ClkMux I__2158 (
            .O(N__9144),
            .I(N__9034));
    ClkMux I__2157 (
            .O(N__9143),
            .I(N__9034));
    ClkMux I__2156 (
            .O(N__9142),
            .I(N__9034));
    ClkMux I__2155 (
            .O(N__9141),
            .I(N__9034));
    ClkMux I__2154 (
            .O(N__9140),
            .I(N__9034));
    ClkMux I__2153 (
            .O(N__9139),
            .I(N__9034));
    Glb2LocalMux I__2152 (
            .O(N__9136),
            .I(N__9034));
    ClkMux I__2151 (
            .O(N__9135),
            .I(N__9034));
    ClkMux I__2150 (
            .O(N__9134),
            .I(N__9034));
    ClkMux I__2149 (
            .O(N__9133),
            .I(N__9034));
    ClkMux I__2148 (
            .O(N__9132),
            .I(N__9034));
    ClkMux I__2147 (
            .O(N__9131),
            .I(N__9034));
    ClkMux I__2146 (
            .O(N__9130),
            .I(N__9034));
    ClkMux I__2145 (
            .O(N__9129),
            .I(N__9034));
    ClkMux I__2144 (
            .O(N__9128),
            .I(N__9034));
    ClkMux I__2143 (
            .O(N__9127),
            .I(N__9034));
    ClkMux I__2142 (
            .O(N__9126),
            .I(N__9034));
    ClkMux I__2141 (
            .O(N__9125),
            .I(N__9034));
    ClkMux I__2140 (
            .O(N__9124),
            .I(N__9034));
    ClkMux I__2139 (
            .O(N__9123),
            .I(N__9034));
    ClkMux I__2138 (
            .O(N__9122),
            .I(N__9034));
    ClkMux I__2137 (
            .O(N__9121),
            .I(N__9034));
    ClkMux I__2136 (
            .O(N__9120),
            .I(N__9034));
    ClkMux I__2135 (
            .O(N__9119),
            .I(N__9034));
    ClkMux I__2134 (
            .O(N__9118),
            .I(N__9034));
    ClkMux I__2133 (
            .O(N__9117),
            .I(N__9034));
    GlobalMux I__2132 (
            .O(N__9034),
            .I(CLK80_OUT));
    CascadeMux I__2131 (
            .O(N__9031),
            .I(N__9024));
    InMux I__2130 (
            .O(N__9030),
            .I(N__9013));
    InMux I__2129 (
            .O(N__9029),
            .I(N__9013));
    InMux I__2128 (
            .O(N__9028),
            .I(N__9010));
    InMux I__2127 (
            .O(N__9027),
            .I(N__9005));
    InMux I__2126 (
            .O(N__9024),
            .I(N__9005));
    InMux I__2125 (
            .O(N__9023),
            .I(N__9002));
    InMux I__2124 (
            .O(N__9022),
            .I(N__8997));
    InMux I__2123 (
            .O(N__9021),
            .I(N__8997));
    InMux I__2122 (
            .O(N__9020),
            .I(N__8994));
    InMux I__2121 (
            .O(N__9019),
            .I(N__8991));
    InMux I__2120 (
            .O(N__9018),
            .I(N__8988));
    LocalMux I__2119 (
            .O(N__9013),
            .I(N__8973));
    LocalMux I__2118 (
            .O(N__9010),
            .I(N__8970));
    LocalMux I__2117 (
            .O(N__9005),
            .I(N__8962));
    LocalMux I__2116 (
            .O(N__9002),
            .I(N__8959));
    LocalMux I__2115 (
            .O(N__8997),
            .I(N__8953));
    LocalMux I__2114 (
            .O(N__8994),
            .I(N__8948));
    LocalMux I__2113 (
            .O(N__8991),
            .I(N__8940));
    LocalMux I__2112 (
            .O(N__8988),
            .I(N__8930));
    SRMux I__2111 (
            .O(N__8987),
            .I(N__8842));
    SRMux I__2110 (
            .O(N__8986),
            .I(N__8842));
    SRMux I__2109 (
            .O(N__8985),
            .I(N__8842));
    SRMux I__2108 (
            .O(N__8984),
            .I(N__8842));
    SRMux I__2107 (
            .O(N__8983),
            .I(N__8842));
    SRMux I__2106 (
            .O(N__8982),
            .I(N__8842));
    SRMux I__2105 (
            .O(N__8981),
            .I(N__8842));
    SRMux I__2104 (
            .O(N__8980),
            .I(N__8842));
    SRMux I__2103 (
            .O(N__8979),
            .I(N__8842));
    SRMux I__2102 (
            .O(N__8978),
            .I(N__8842));
    SRMux I__2101 (
            .O(N__8977),
            .I(N__8842));
    SRMux I__2100 (
            .O(N__8976),
            .I(N__8842));
    Glb2LocalMux I__2099 (
            .O(N__8973),
            .I(N__8842));
    Glb2LocalMux I__2098 (
            .O(N__8970),
            .I(N__8842));
    SRMux I__2097 (
            .O(N__8969),
            .I(N__8842));
    SRMux I__2096 (
            .O(N__8968),
            .I(N__8842));
    SRMux I__2095 (
            .O(N__8967),
            .I(N__8842));
    SRMux I__2094 (
            .O(N__8966),
            .I(N__8842));
    SRMux I__2093 (
            .O(N__8965),
            .I(N__8842));
    Glb2LocalMux I__2092 (
            .O(N__8962),
            .I(N__8842));
    Glb2LocalMux I__2091 (
            .O(N__8959),
            .I(N__8842));
    SRMux I__2090 (
            .O(N__8958),
            .I(N__8842));
    SRMux I__2089 (
            .O(N__8957),
            .I(N__8842));
    SRMux I__2088 (
            .O(N__8956),
            .I(N__8842));
    Glb2LocalMux I__2087 (
            .O(N__8953),
            .I(N__8842));
    SRMux I__2086 (
            .O(N__8952),
            .I(N__8842));
    SRMux I__2085 (
            .O(N__8951),
            .I(N__8842));
    Glb2LocalMux I__2084 (
            .O(N__8948),
            .I(N__8842));
    SRMux I__2083 (
            .O(N__8947),
            .I(N__8842));
    SRMux I__2082 (
            .O(N__8946),
            .I(N__8842));
    SRMux I__2081 (
            .O(N__8945),
            .I(N__8842));
    SRMux I__2080 (
            .O(N__8944),
            .I(N__8842));
    SRMux I__2079 (
            .O(N__8943),
            .I(N__8842));
    Glb2LocalMux I__2078 (
            .O(N__8940),
            .I(N__8842));
    SRMux I__2077 (
            .O(N__8939),
            .I(N__8842));
    SRMux I__2076 (
            .O(N__8938),
            .I(N__8842));
    SRMux I__2075 (
            .O(N__8937),
            .I(N__8842));
    SRMux I__2074 (
            .O(N__8936),
            .I(N__8842));
    SRMux I__2073 (
            .O(N__8935),
            .I(N__8842));
    SRMux I__2072 (
            .O(N__8934),
            .I(N__8842));
    SRMux I__2071 (
            .O(N__8933),
            .I(N__8842));
    Glb2LocalMux I__2070 (
            .O(N__8930),
            .I(N__8842));
    SRMux I__2069 (
            .O(N__8929),
            .I(N__8842));
    GlobalMux I__2068 (
            .O(N__8842),
            .I(N__8839));
    gio2CtrlBuf I__2067 (
            .O(N__8839),
            .I(RESETn_c_i_g));
    IoInMux I__2066 (
            .O(N__8836),
            .I(N__8833));
    LocalMux I__2065 (
            .O(N__8833),
            .I(N__8830));
    Span4Mux_s1_v I__2064 (
            .O(N__8830),
            .I(N__8826));
    IoInMux I__2063 (
            .O(N__8829),
            .I(N__8823));
    Span4Mux_v I__2062 (
            .O(N__8826),
            .I(N__8820));
    LocalMux I__2061 (
            .O(N__8823),
            .I(N__8817));
    Span4Mux_v I__2060 (
            .O(N__8820),
            .I(N__8814));
    Span4Mux_s3_h I__2059 (
            .O(N__8817),
            .I(N__8811));
    Span4Mux_h I__2058 (
            .O(N__8814),
            .I(N__8808));
    Span4Mux_v I__2057 (
            .O(N__8811),
            .I(N__8805));
    Odrv4 I__2056 (
            .O(N__8808),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2055 (
            .O(N__8805),
            .I(CONSTANT_ONE_NET));
    InMux I__2054 (
            .O(N__8800),
            .I(N__8797));
    LocalMux I__2053 (
            .O(N__8797),
            .I(N__8793));
    InMux I__2052 (
            .O(N__8796),
            .I(N__8790));
    Span4Mux_v I__2051 (
            .O(N__8793),
            .I(N__8787));
    LocalMux I__2050 (
            .O(N__8790),
            .I(N__8784));
    Sp12to4 I__2049 (
            .O(N__8787),
            .I(N__8781));
    Span12Mux_v I__2048 (
            .O(N__8784),
            .I(N__8778));
    Span12Mux_h I__2047 (
            .O(N__8781),
            .I(N__8775));
    Span12Mux_h I__2046 (
            .O(N__8778),
            .I(N__8772));
    Odrv12 I__2045 (
            .O(N__8775),
            .I(DRA_c_7));
    Odrv12 I__2044 (
            .O(N__8772),
            .I(DRA_c_7));
    InMux I__2043 (
            .O(N__8767),
            .I(N__8764));
    LocalMux I__2042 (
            .O(N__8764),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2041 (
            .O(N__8761),
            .I(N__8758));
    LocalMux I__2040 (
            .O(N__8758),
            .I(N__8754));
    InMux I__2039 (
            .O(N__8757),
            .I(N__8751));
    Span4Mux_h I__2038 (
            .O(N__8754),
            .I(N__8746));
    LocalMux I__2037 (
            .O(N__8751),
            .I(N__8746));
    Span4Mux_v I__2036 (
            .O(N__8746),
            .I(N__8743));
    Sp12to4 I__2035 (
            .O(N__8743),
            .I(N__8740));
    Odrv12 I__2034 (
            .O(N__8740),
            .I(DRA_c_8));
    InMux I__2033 (
            .O(N__8737),
            .I(N__8734));
    LocalMux I__2032 (
            .O(N__8734),
            .I(N__8731));
    Odrv4 I__2031 (
            .O(N__8731),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    CEMux I__2030 (
            .O(N__8728),
            .I(N__8723));
    CEMux I__2029 (
            .O(N__8727),
            .I(N__8720));
    CEMux I__2028 (
            .O(N__8726),
            .I(N__8717));
    LocalMux I__2027 (
            .O(N__8723),
            .I(N__8714));
    LocalMux I__2026 (
            .O(N__8720),
            .I(N__8711));
    LocalMux I__2025 (
            .O(N__8717),
            .I(N__8708));
    Span4Mux_v I__2024 (
            .O(N__8714),
            .I(N__8705));
    Span4Mux_h I__2023 (
            .O(N__8711),
            .I(N__8702));
    Span4Mux_v I__2022 (
            .O(N__8708),
            .I(N__8699));
    Odrv4 I__2021 (
            .O(N__8705),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    Odrv4 I__2020 (
            .O(N__8702),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    Odrv4 I__2019 (
            .O(N__8699),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    InMux I__2018 (
            .O(N__8692),
            .I(N__8689));
    LocalMux I__2017 (
            .O(N__8689),
            .I(N__8685));
    InMux I__2016 (
            .O(N__8688),
            .I(N__8682));
    Span4Mux_v I__2015 (
            .O(N__8685),
            .I(N__8679));
    LocalMux I__2014 (
            .O(N__8682),
            .I(N__8676));
    Sp12to4 I__2013 (
            .O(N__8679),
            .I(N__8673));
    Span4Mux_h I__2012 (
            .O(N__8676),
            .I(N__8670));
    Span12Mux_h I__2011 (
            .O(N__8673),
            .I(N__8667));
    Sp12to4 I__2010 (
            .O(N__8670),
            .I(N__8664));
    Span12Mux_v I__2009 (
            .O(N__8667),
            .I(N__8661));
    Span12Mux_v I__2008 (
            .O(N__8664),
            .I(N__8658));
    Odrv12 I__2007 (
            .O(N__8661),
            .I(DRA_c_3));
    Odrv12 I__2006 (
            .O(N__8658),
            .I(DRA_c_3));
    InMux I__2005 (
            .O(N__8653),
            .I(N__8650));
    LocalMux I__2004 (
            .O(N__8650),
            .I(N__8647));
    Span4Mux_h I__2003 (
            .O(N__8647),
            .I(N__8644));
    Odrv4 I__2002 (
            .O(N__8644),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    CEMux I__2001 (
            .O(N__8641),
            .I(N__8637));
    CEMux I__2000 (
            .O(N__8640),
            .I(N__8632));
    LocalMux I__1999 (
            .O(N__8637),
            .I(N__8629));
    CEMux I__1998 (
            .O(N__8636),
            .I(N__8626));
    CEMux I__1997 (
            .O(N__8635),
            .I(N__8623));
    LocalMux I__1996 (
            .O(N__8632),
            .I(N__8619));
    Span4Mux_h I__1995 (
            .O(N__8629),
            .I(N__8612));
    LocalMux I__1994 (
            .O(N__8626),
            .I(N__8612));
    LocalMux I__1993 (
            .O(N__8623),
            .I(N__8612));
    CEMux I__1992 (
            .O(N__8622),
            .I(N__8609));
    Span4Mux_h I__1991 (
            .O(N__8619),
            .I(N__8606));
    Span4Mux_v I__1990 (
            .O(N__8612),
            .I(N__8603));
    LocalMux I__1989 (
            .O(N__8609),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    Odrv4 I__1988 (
            .O(N__8606),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    Odrv4 I__1987 (
            .O(N__8603),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    InMux I__1986 (
            .O(N__8596),
            .I(N__8592));
    CascadeMux I__1985 (
            .O(N__8595),
            .I(N__8589));
    LocalMux I__1984 (
            .O(N__8592),
            .I(N__8580));
    InMux I__1983 (
            .O(N__8589),
            .I(N__8577));
    CascadeMux I__1982 (
            .O(N__8588),
            .I(N__8572));
    CascadeMux I__1981 (
            .O(N__8587),
            .I(N__8569));
    CascadeMux I__1980 (
            .O(N__8586),
            .I(N__8566));
    CascadeMux I__1979 (
            .O(N__8585),
            .I(N__8563));
    InMux I__1978 (
            .O(N__8584),
            .I(N__8556));
    InMux I__1977 (
            .O(N__8583),
            .I(N__8556));
    Span4Mux_h I__1976 (
            .O(N__8580),
            .I(N__8551));
    LocalMux I__1975 (
            .O(N__8577),
            .I(N__8551));
    InMux I__1974 (
            .O(N__8576),
            .I(N__8546));
    InMux I__1973 (
            .O(N__8575),
            .I(N__8546));
    InMux I__1972 (
            .O(N__8572),
            .I(N__8543));
    InMux I__1971 (
            .O(N__8569),
            .I(N__8540));
    InMux I__1970 (
            .O(N__8566),
            .I(N__8534));
    InMux I__1969 (
            .O(N__8563),
            .I(N__8531));
    CascadeMux I__1968 (
            .O(N__8562),
            .I(N__8528));
    CascadeMux I__1967 (
            .O(N__8561),
            .I(N__8525));
    LocalMux I__1966 (
            .O(N__8556),
            .I(N__8521));
    Span4Mux_v I__1965 (
            .O(N__8551),
            .I(N__8518));
    LocalMux I__1964 (
            .O(N__8546),
            .I(N__8513));
    LocalMux I__1963 (
            .O(N__8543),
            .I(N__8513));
    LocalMux I__1962 (
            .O(N__8540),
            .I(N__8510));
    InMux I__1961 (
            .O(N__8539),
            .I(N__8503));
    InMux I__1960 (
            .O(N__8538),
            .I(N__8503));
    InMux I__1959 (
            .O(N__8537),
            .I(N__8503));
    LocalMux I__1958 (
            .O(N__8534),
            .I(N__8498));
    LocalMux I__1957 (
            .O(N__8531),
            .I(N__8498));
    InMux I__1956 (
            .O(N__8528),
            .I(N__8493));
    InMux I__1955 (
            .O(N__8525),
            .I(N__8493));
    InMux I__1954 (
            .O(N__8524),
            .I(N__8490));
    Span4Mux_v I__1953 (
            .O(N__8521),
            .I(N__8487));
    Span4Mux_v I__1952 (
            .O(N__8518),
            .I(N__8484));
    Span4Mux_v I__1951 (
            .O(N__8513),
            .I(N__8475));
    Span4Mux_h I__1950 (
            .O(N__8510),
            .I(N__8475));
    LocalMux I__1949 (
            .O(N__8503),
            .I(N__8475));
    Span4Mux_h I__1948 (
            .O(N__8498),
            .I(N__8475));
    LocalMux I__1947 (
            .O(N__8493),
            .I(N__8472));
    LocalMux I__1946 (
            .O(N__8490),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1945 (
            .O(N__8487),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1944 (
            .O(N__8484),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1943 (
            .O(N__8475),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1942 (
            .O(N__8472),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    IoInMux I__1941 (
            .O(N__8461),
            .I(N__8458));
    LocalMux I__1940 (
            .O(N__8458),
            .I(N__8455));
    Span4Mux_s3_v I__1939 (
            .O(N__8455),
            .I(N__8452));
    Span4Mux_v I__1938 (
            .O(N__8452),
            .I(N__8449));
    Span4Mux_h I__1937 (
            .O(N__8449),
            .I(N__8446));
    Odrv4 I__1936 (
            .O(N__8446),
            .I(CASn_c));
    CascadeMux I__1935 (
            .O(N__8443),
            .I(N__8438));
    CascadeMux I__1934 (
            .O(N__8442),
            .I(N__8432));
    InMux I__1933 (
            .O(N__8441),
            .I(N__8427));
    InMux I__1932 (
            .O(N__8438),
            .I(N__8420));
    InMux I__1931 (
            .O(N__8437),
            .I(N__8420));
    CascadeMux I__1930 (
            .O(N__8436),
            .I(N__8416));
    InMux I__1929 (
            .O(N__8435),
            .I(N__8413));
    InMux I__1928 (
            .O(N__8432),
            .I(N__8410));
    InMux I__1927 (
            .O(N__8431),
            .I(N__8405));
    InMux I__1926 (
            .O(N__8430),
            .I(N__8405));
    LocalMux I__1925 (
            .O(N__8427),
            .I(N__8402));
    CascadeMux I__1924 (
            .O(N__8426),
            .I(N__8399));
    CascadeMux I__1923 (
            .O(N__8425),
            .I(N__8394));
    LocalMux I__1922 (
            .O(N__8420),
            .I(N__8391));
    InMux I__1921 (
            .O(N__8419),
            .I(N__8386));
    InMux I__1920 (
            .O(N__8416),
            .I(N__8386));
    LocalMux I__1919 (
            .O(N__8413),
            .I(N__8377));
    LocalMux I__1918 (
            .O(N__8410),
            .I(N__8377));
    LocalMux I__1917 (
            .O(N__8405),
            .I(N__8377));
    Span4Mux_h I__1916 (
            .O(N__8402),
            .I(N__8377));
    InMux I__1915 (
            .O(N__8399),
            .I(N__8370));
    InMux I__1914 (
            .O(N__8398),
            .I(N__8370));
    InMux I__1913 (
            .O(N__8397),
            .I(N__8370));
    InMux I__1912 (
            .O(N__8394),
            .I(N__8367));
    Span4Mux_v I__1911 (
            .O(N__8391),
            .I(N__8364));
    LocalMux I__1910 (
            .O(N__8386),
            .I(N__8357));
    Sp12to4 I__1909 (
            .O(N__8377),
            .I(N__8357));
    LocalMux I__1908 (
            .O(N__8370),
            .I(N__8357));
    LocalMux I__1907 (
            .O(N__8367),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1906 (
            .O(N__8364),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv12 I__1905 (
            .O(N__8357),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__1904 (
            .O(N__8350),
            .I(N__8347));
    LocalMux I__1903 (
            .O(N__8347),
            .I(N__8344));
    Span4Mux_s3_h I__1902 (
            .O(N__8344),
            .I(N__8341));
    Span4Mux_v I__1901 (
            .O(N__8341),
            .I(N__8338));
    Span4Mux_v I__1900 (
            .O(N__8338),
            .I(N__8335));
    Span4Mux_h I__1899 (
            .O(N__8335),
            .I(N__8332));
    Odrv4 I__1898 (
            .O(N__8332),
            .I(WEn_c));
    InMux I__1897 (
            .O(N__8329),
            .I(N__8325));
    InMux I__1896 (
            .O(N__8328),
            .I(N__8322));
    LocalMux I__1895 (
            .O(N__8325),
            .I(N__8318));
    LocalMux I__1894 (
            .O(N__8322),
            .I(N__8315));
    InMux I__1893 (
            .O(N__8321),
            .I(N__8312));
    Span4Mux_h I__1892 (
            .O(N__8318),
            .I(N__8304));
    Span4Mux_h I__1891 (
            .O(N__8315),
            .I(N__8304));
    LocalMux I__1890 (
            .O(N__8312),
            .I(N__8304));
    InMux I__1889 (
            .O(N__8311),
            .I(N__8301));
    Odrv4 I__1888 (
            .O(N__8304),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1887 (
            .O(N__8301),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__1886 (
            .O(N__8296),
            .I(N__8293));
    LocalMux I__1885 (
            .O(N__8293),
            .I(N__8290));
    Span4Mux_s2_v I__1884 (
            .O(N__8290),
            .I(N__8287));
    Span4Mux_v I__1883 (
            .O(N__8287),
            .I(N__8284));
    Span4Mux_v I__1882 (
            .O(N__8284),
            .I(N__8281));
    Odrv4 I__1881 (
            .O(N__8281),
            .I(CRCSn_c));
    InMux I__1880 (
            .O(N__8278),
            .I(N__8274));
    InMux I__1879 (
            .O(N__8277),
            .I(N__8271));
    LocalMux I__1878 (
            .O(N__8274),
            .I(N__8268));
    LocalMux I__1877 (
            .O(N__8271),
            .I(N__8265));
    Span4Mux_v I__1876 (
            .O(N__8268),
            .I(N__8262));
    Span4Mux_v I__1875 (
            .O(N__8265),
            .I(N__8259));
    Sp12to4 I__1874 (
            .O(N__8262),
            .I(N__8254));
    Sp12to4 I__1873 (
            .O(N__8259),
            .I(N__8254));
    Span12Mux_h I__1872 (
            .O(N__8254),
            .I(N__8251));
    Odrv12 I__1871 (
            .O(N__8251),
            .I(RAS0n_c));
    InMux I__1870 (
            .O(N__8248),
            .I(N__8245));
    LocalMux I__1869 (
            .O(N__8245),
            .I(N__8242));
    Span12Mux_h I__1868 (
            .O(N__8242),
            .I(N__8239));
    Odrv12 I__1867 (
            .O(N__8239),
            .I(RAS1n_c));
    InMux I__1866 (
            .O(N__8236),
            .I(N__8232));
    InMux I__1865 (
            .O(N__8235),
            .I(N__8227));
    LocalMux I__1864 (
            .O(N__8232),
            .I(N__8221));
    InMux I__1863 (
            .O(N__8231),
            .I(N__8218));
    InMux I__1862 (
            .O(N__8230),
            .I(N__8215));
    LocalMux I__1861 (
            .O(N__8227),
            .I(N__8212));
    InMux I__1860 (
            .O(N__8226),
            .I(N__8209));
    InMux I__1859 (
            .O(N__8225),
            .I(N__8206));
    InMux I__1858 (
            .O(N__8224),
            .I(N__8203));
    Span4Mux_v I__1857 (
            .O(N__8221),
            .I(N__8198));
    LocalMux I__1856 (
            .O(N__8218),
            .I(N__8198));
    LocalMux I__1855 (
            .O(N__8215),
            .I(N__8195));
    Span4Mux_v I__1854 (
            .O(N__8212),
            .I(N__8192));
    LocalMux I__1853 (
            .O(N__8209),
            .I(N__8189));
    LocalMux I__1852 (
            .O(N__8206),
            .I(N__8184));
    LocalMux I__1851 (
            .O(N__8203),
            .I(N__8184));
    Span4Mux_v I__1850 (
            .O(N__8198),
            .I(N__8179));
    Span4Mux_v I__1849 (
            .O(N__8195),
            .I(N__8179));
    Span4Mux_h I__1848 (
            .O(N__8192),
            .I(N__8172));
    Span4Mux_v I__1847 (
            .O(N__8189),
            .I(N__8172));
    Span4Mux_v I__1846 (
            .O(N__8184),
            .I(N__8172));
    Sp12to4 I__1845 (
            .O(N__8179),
            .I(N__8169));
    Sp12to4 I__1844 (
            .O(N__8172),
            .I(N__8166));
    Span12Mux_h I__1843 (
            .O(N__8169),
            .I(N__8163));
    Span12Mux_h I__1842 (
            .O(N__8166),
            .I(N__8160));
    Odrv12 I__1841 (
            .O(N__8163),
            .I(RESETn_c));
    Odrv12 I__1840 (
            .O(N__8160),
            .I(RESETn_c));
    CascadeMux I__1839 (
            .O(N__8155),
            .I(\U712_CHIP_RAM.N_274_cascade_ ));
    CascadeMux I__1838 (
            .O(N__8152),
            .I(N__8149));
    InMux I__1837 (
            .O(N__8149),
            .I(N__8145));
    InMux I__1836 (
            .O(N__8148),
            .I(N__8142));
    LocalMux I__1835 (
            .O(N__8145),
            .I(N__8138));
    LocalMux I__1834 (
            .O(N__8142),
            .I(N__8135));
    InMux I__1833 (
            .O(N__8141),
            .I(N__8132));
    Odrv4 I__1832 (
            .O(N__8138),
            .I(\U712_CHIP_RAM.N_337 ));
    Odrv4 I__1831 (
            .O(N__8135),
            .I(\U712_CHIP_RAM.N_337 ));
    LocalMux I__1830 (
            .O(N__8132),
            .I(\U712_CHIP_RAM.N_337 ));
    CascadeMux I__1829 (
            .O(N__8125),
            .I(\U712_CHIP_RAM.N_337_cascade_ ));
    InMux I__1828 (
            .O(N__8122),
            .I(N__8119));
    LocalMux I__1827 (
            .O(N__8119),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_2_0 ));
    CascadeMux I__1826 (
            .O(N__8116),
            .I(N__8109));
    CascadeMux I__1825 (
            .O(N__8115),
            .I(N__8106));
    CascadeMux I__1824 (
            .O(N__8114),
            .I(N__8103));
    InMux I__1823 (
            .O(N__8113),
            .I(N__8100));
    InMux I__1822 (
            .O(N__8112),
            .I(N__8095));
    InMux I__1821 (
            .O(N__8109),
            .I(N__8090));
    InMux I__1820 (
            .O(N__8106),
            .I(N__8090));
    InMux I__1819 (
            .O(N__8103),
            .I(N__8083));
    LocalMux I__1818 (
            .O(N__8100),
            .I(N__8080));
    InMux I__1817 (
            .O(N__8099),
            .I(N__8075));
    InMux I__1816 (
            .O(N__8098),
            .I(N__8075));
    LocalMux I__1815 (
            .O(N__8095),
            .I(N__8072));
    LocalMux I__1814 (
            .O(N__8090),
            .I(N__8069));
    InMux I__1813 (
            .O(N__8089),
            .I(N__8066));
    InMux I__1812 (
            .O(N__8088),
            .I(N__8063));
    InMux I__1811 (
            .O(N__8087),
            .I(N__8060));
    InMux I__1810 (
            .O(N__8086),
            .I(N__8057));
    LocalMux I__1809 (
            .O(N__8083),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1808 (
            .O(N__8080),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1807 (
            .O(N__8075),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1806 (
            .O(N__8072),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1805 (
            .O(N__8069),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1804 (
            .O(N__8066),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1803 (
            .O(N__8063),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1802 (
            .O(N__8060),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1801 (
            .O(N__8057),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__1800 (
            .O(N__8038),
            .I(N__8031));
    InMux I__1799 (
            .O(N__8037),
            .I(N__8028));
    InMux I__1798 (
            .O(N__8036),
            .I(N__8021));
    InMux I__1797 (
            .O(N__8035),
            .I(N__8021));
    InMux I__1796 (
            .O(N__8034),
            .I(N__8021));
    LocalMux I__1795 (
            .O(N__8031),
            .I(N__8018));
    LocalMux I__1794 (
            .O(N__8028),
            .I(N__8013));
    LocalMux I__1793 (
            .O(N__8021),
            .I(N__8008));
    Span4Mux_h I__1792 (
            .O(N__8018),
            .I(N__8008));
    InMux I__1791 (
            .O(N__8017),
            .I(N__8005));
    InMux I__1790 (
            .O(N__8016),
            .I(N__8002));
    Odrv4 I__1789 (
            .O(N__8013),
            .I(\U712_CHIP_RAM.N_271 ));
    Odrv4 I__1788 (
            .O(N__8008),
            .I(\U712_CHIP_RAM.N_271 ));
    LocalMux I__1787 (
            .O(N__8005),
            .I(\U712_CHIP_RAM.N_271 ));
    LocalMux I__1786 (
            .O(N__8002),
            .I(\U712_CHIP_RAM.N_271 ));
    CascadeMux I__1785 (
            .O(N__7993),
            .I(N__7985));
    InMux I__1784 (
            .O(N__7992),
            .I(N__7982));
    InMux I__1783 (
            .O(N__7991),
            .I(N__7979));
    InMux I__1782 (
            .O(N__7990),
            .I(N__7970));
    InMux I__1781 (
            .O(N__7989),
            .I(N__7965));
    InMux I__1780 (
            .O(N__7988),
            .I(N__7965));
    InMux I__1779 (
            .O(N__7985),
            .I(N__7962));
    LocalMux I__1778 (
            .O(N__7982),
            .I(N__7959));
    LocalMux I__1777 (
            .O(N__7979),
            .I(N__7956));
    InMux I__1776 (
            .O(N__7978),
            .I(N__7951));
    InMux I__1775 (
            .O(N__7977),
            .I(N__7951));
    InMux I__1774 (
            .O(N__7976),
            .I(N__7948));
    InMux I__1773 (
            .O(N__7975),
            .I(N__7945));
    InMux I__1772 (
            .O(N__7974),
            .I(N__7940));
    InMux I__1771 (
            .O(N__7973),
            .I(N__7940));
    LocalMux I__1770 (
            .O(N__7970),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1769 (
            .O(N__7965),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1768 (
            .O(N__7962),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv12 I__1767 (
            .O(N__7959),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv12 I__1766 (
            .O(N__7956),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1765 (
            .O(N__7951),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1764 (
            .O(N__7948),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1763 (
            .O(N__7945),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1762 (
            .O(N__7940),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    CascadeMux I__1761 (
            .O(N__7921),
            .I(N__7917));
    InMux I__1760 (
            .O(N__7920),
            .I(N__7910));
    InMux I__1759 (
            .O(N__7917),
            .I(N__7910));
    InMux I__1758 (
            .O(N__7916),
            .I(N__7905));
    InMux I__1757 (
            .O(N__7915),
            .I(N__7905));
    LocalMux I__1756 (
            .O(N__7910),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1755 (
            .O(N__7905),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__1754 (
            .O(N__7900),
            .I(N__7894));
    InMux I__1753 (
            .O(N__7899),
            .I(N__7891));
    InMux I__1752 (
            .O(N__7898),
            .I(N__7886));
    InMux I__1751 (
            .O(N__7897),
            .I(N__7886));
    LocalMux I__1750 (
            .O(N__7894),
            .I(N__7883));
    LocalMux I__1749 (
            .O(N__7891),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c3 ));
    LocalMux I__1748 (
            .O(N__7886),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c3 ));
    Odrv4 I__1747 (
            .O(N__7883),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c3 ));
    CascadeMux I__1746 (
            .O(N__7876),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_ ));
    CascadeMux I__1745 (
            .O(N__7873),
            .I(N__7870));
    InMux I__1744 (
            .O(N__7870),
            .I(N__7866));
    InMux I__1743 (
            .O(N__7869),
            .I(N__7863));
    LocalMux I__1742 (
            .O(N__7866),
            .I(N__7857));
    LocalMux I__1741 (
            .O(N__7863),
            .I(N__7857));
    InMux I__1740 (
            .O(N__7862),
            .I(N__7854));
    Odrv4 I__1739 (
            .O(N__7857),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__1738 (
            .O(N__7854),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__1737 (
            .O(N__7849),
            .I(N__7843));
    CascadeMux I__1736 (
            .O(N__7848),
            .I(N__7840));
    InMux I__1735 (
            .O(N__7847),
            .I(N__7833));
    InMux I__1734 (
            .O(N__7846),
            .I(N__7833));
    InMux I__1733 (
            .O(N__7843),
            .I(N__7828));
    InMux I__1732 (
            .O(N__7840),
            .I(N__7828));
    CascadeMux I__1731 (
            .O(N__7839),
            .I(N__7824));
    CascadeMux I__1730 (
            .O(N__7838),
            .I(N__7820));
    LocalMux I__1729 (
            .O(N__7833),
            .I(N__7814));
    LocalMux I__1728 (
            .O(N__7828),
            .I(N__7814));
    CascadeMux I__1727 (
            .O(N__7827),
            .I(N__7810));
    InMux I__1726 (
            .O(N__7824),
            .I(N__7804));
    InMux I__1725 (
            .O(N__7823),
            .I(N__7801));
    InMux I__1724 (
            .O(N__7820),
            .I(N__7796));
    InMux I__1723 (
            .O(N__7819),
            .I(N__7796));
    Span4Mux_h I__1722 (
            .O(N__7814),
            .I(N__7793));
    InMux I__1721 (
            .O(N__7813),
            .I(N__7788));
    InMux I__1720 (
            .O(N__7810),
            .I(N__7788));
    InMux I__1719 (
            .O(N__7809),
            .I(N__7785));
    InMux I__1718 (
            .O(N__7808),
            .I(N__7780));
    InMux I__1717 (
            .O(N__7807),
            .I(N__7780));
    LocalMux I__1716 (
            .O(N__7804),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1715 (
            .O(N__7801),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1714 (
            .O(N__7796),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1713 (
            .O(N__7793),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1712 (
            .O(N__7788),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1711 (
            .O(N__7785),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1710 (
            .O(N__7780),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__1709 (
            .O(N__7765),
            .I(N__7762));
    LocalMux I__1708 (
            .O(N__7762),
            .I(N__7758));
    InMux I__1707 (
            .O(N__7761),
            .I(N__7754));
    Span4Mux_v I__1706 (
            .O(N__7758),
            .I(N__7751));
    InMux I__1705 (
            .O(N__7757),
            .I(N__7748));
    LocalMux I__1704 (
            .O(N__7754),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER46 ));
    Odrv4 I__1703 (
            .O(N__7751),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER46 ));
    LocalMux I__1702 (
            .O(N__7748),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER46 ));
    CascadeMux I__1701 (
            .O(N__7741),
            .I(N__7736));
    CascadeMux I__1700 (
            .O(N__7740),
            .I(N__7727));
    InMux I__1699 (
            .O(N__7739),
            .I(N__7723));
    InMux I__1698 (
            .O(N__7736),
            .I(N__7717));
    CascadeMux I__1697 (
            .O(N__7735),
            .I(N__7713));
    InMux I__1696 (
            .O(N__7734),
            .I(N__7710));
    InMux I__1695 (
            .O(N__7733),
            .I(N__7703));
    InMux I__1694 (
            .O(N__7732),
            .I(N__7703));
    InMux I__1693 (
            .O(N__7731),
            .I(N__7703));
    CascadeMux I__1692 (
            .O(N__7730),
            .I(N__7691));
    InMux I__1691 (
            .O(N__7727),
            .I(N__7688));
    InMux I__1690 (
            .O(N__7726),
            .I(N__7685));
    LocalMux I__1689 (
            .O(N__7723),
            .I(N__7682));
    InMux I__1688 (
            .O(N__7722),
            .I(N__7679));
    InMux I__1687 (
            .O(N__7721),
            .I(N__7674));
    InMux I__1686 (
            .O(N__7720),
            .I(N__7674));
    LocalMux I__1685 (
            .O(N__7717),
            .I(N__7671));
    InMux I__1684 (
            .O(N__7716),
            .I(N__7668));
    InMux I__1683 (
            .O(N__7713),
            .I(N__7665));
    LocalMux I__1682 (
            .O(N__7710),
            .I(N__7662));
    LocalMux I__1681 (
            .O(N__7703),
            .I(N__7659));
    InMux I__1680 (
            .O(N__7702),
            .I(N__7652));
    InMux I__1679 (
            .O(N__7701),
            .I(N__7652));
    InMux I__1678 (
            .O(N__7700),
            .I(N__7652));
    InMux I__1677 (
            .O(N__7699),
            .I(N__7649));
    InMux I__1676 (
            .O(N__7698),
            .I(N__7644));
    InMux I__1675 (
            .O(N__7697),
            .I(N__7644));
    InMux I__1674 (
            .O(N__7696),
            .I(N__7641));
    InMux I__1673 (
            .O(N__7695),
            .I(N__7636));
    InMux I__1672 (
            .O(N__7694),
            .I(N__7636));
    InMux I__1671 (
            .O(N__7691),
            .I(N__7633));
    LocalMux I__1670 (
            .O(N__7688),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1669 (
            .O(N__7685),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1668 (
            .O(N__7682),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1667 (
            .O(N__7679),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1666 (
            .O(N__7674),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1665 (
            .O(N__7671),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1664 (
            .O(N__7668),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1663 (
            .O(N__7665),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1662 (
            .O(N__7662),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1661 (
            .O(N__7659),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1660 (
            .O(N__7652),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1659 (
            .O(N__7649),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1658 (
            .O(N__7644),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1657 (
            .O(N__7641),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1656 (
            .O(N__7636),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1655 (
            .O(N__7633),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__1654 (
            .O(N__7600),
            .I(N__7596));
    InMux I__1653 (
            .O(N__7599),
            .I(N__7593));
    LocalMux I__1652 (
            .O(N__7596),
            .I(N__7590));
    LocalMux I__1651 (
            .O(N__7593),
            .I(\U712_CHIP_RAM.N_303 ));
    Odrv4 I__1650 (
            .O(N__7590),
            .I(\U712_CHIP_RAM.N_303 ));
    InMux I__1649 (
            .O(N__7585),
            .I(N__7576));
    InMux I__1648 (
            .O(N__7584),
            .I(N__7573));
    InMux I__1647 (
            .O(N__7583),
            .I(N__7567));
    InMux I__1646 (
            .O(N__7582),
            .I(N__7567));
    InMux I__1645 (
            .O(N__7581),
            .I(N__7564));
    InMux I__1644 (
            .O(N__7580),
            .I(N__7561));
    InMux I__1643 (
            .O(N__7579),
            .I(N__7558));
    LocalMux I__1642 (
            .O(N__7576),
            .I(N__7555));
    LocalMux I__1641 (
            .O(N__7573),
            .I(N__7552));
    InMux I__1640 (
            .O(N__7572),
            .I(N__7549));
    LocalMux I__1639 (
            .O(N__7567),
            .I(N__7546));
    LocalMux I__1638 (
            .O(N__7564),
            .I(N__7538));
    LocalMux I__1637 (
            .O(N__7561),
            .I(N__7538));
    LocalMux I__1636 (
            .O(N__7558),
            .I(N__7538));
    Span4Mux_v I__1635 (
            .O(N__7555),
            .I(N__7531));
    Span4Mux_v I__1634 (
            .O(N__7552),
            .I(N__7531));
    LocalMux I__1633 (
            .O(N__7549),
            .I(N__7531));
    Span4Mux_v I__1632 (
            .O(N__7546),
            .I(N__7528));
    InMux I__1631 (
            .O(N__7545),
            .I(N__7525));
    Span4Mux_v I__1630 (
            .O(N__7538),
            .I(N__7520));
    Span4Mux_h I__1629 (
            .O(N__7531),
            .I(N__7520));
    Odrv4 I__1628 (
            .O(N__7528),
            .I(DMA_CYCLEm));
    LocalMux I__1627 (
            .O(N__7525),
            .I(DMA_CYCLEm));
    Odrv4 I__1626 (
            .O(N__7520),
            .I(DMA_CYCLEm));
    CascadeMux I__1625 (
            .O(N__7513),
            .I(N__7509));
    InMux I__1624 (
            .O(N__7512),
            .I(N__7506));
    InMux I__1623 (
            .O(N__7509),
            .I(N__7503));
    LocalMux I__1622 (
            .O(N__7506),
            .I(N__7500));
    LocalMux I__1621 (
            .O(N__7503),
            .I(N__7497));
    Span4Mux_v I__1620 (
            .O(N__7500),
            .I(N__7493));
    Span4Mux_v I__1619 (
            .O(N__7497),
            .I(N__7490));
    InMux I__1618 (
            .O(N__7496),
            .I(N__7487));
    Sp12to4 I__1617 (
            .O(N__7493),
            .I(N__7481));
    Sp12to4 I__1616 (
            .O(N__7490),
            .I(N__7481));
    LocalMux I__1615 (
            .O(N__7487),
            .I(N__7478));
    InMux I__1614 (
            .O(N__7486),
            .I(N__7475));
    Odrv12 I__1613 (
            .O(N__7481),
            .I(REG_CYCLEm));
    Odrv12 I__1612 (
            .O(N__7478),
            .I(REG_CYCLEm));
    LocalMux I__1611 (
            .O(N__7475),
            .I(REG_CYCLEm));
    IoInMux I__1610 (
            .O(N__7468),
            .I(N__7465));
    LocalMux I__1609 (
            .O(N__7465),
            .I(N__7462));
    Span12Mux_s4_v I__1608 (
            .O(N__7462),
            .I(N__7459));
    Span12Mux_h I__1607 (
            .O(N__7459),
            .I(N__7456));
    Odrv12 I__1606 (
            .O(N__7456),
            .I(DRDENn_c));
    CascadeMux I__1605 (
            .O(N__7453),
            .I(N__7450));
    InMux I__1604 (
            .O(N__7450),
            .I(N__7447));
    LocalMux I__1603 (
            .O(N__7447),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    CascadeMux I__1602 (
            .O(N__7444),
            .I(\U712_CHIP_RAM.N_284_cascade_ ));
    InMux I__1601 (
            .O(N__7441),
            .I(N__7438));
    LocalMux I__1600 (
            .O(N__7438),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_1_2 ));
    InMux I__1599 (
            .O(N__7435),
            .I(N__7432));
    LocalMux I__1598 (
            .O(N__7432),
            .I(N__7429));
    Odrv12 I__1597 (
            .O(N__7429),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    CascadeMux I__1596 (
            .O(N__7426),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_1_0_cascade_ ));
    InMux I__1595 (
            .O(N__7423),
            .I(N__7420));
    LocalMux I__1594 (
            .O(N__7420),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_0 ));
    CascadeMux I__1593 (
            .O(N__7417),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c6_cascade_ ));
    InMux I__1592 (
            .O(N__7414),
            .I(N__7400));
    InMux I__1591 (
            .O(N__7413),
            .I(N__7400));
    InMux I__1590 (
            .O(N__7412),
            .I(N__7400));
    InMux I__1589 (
            .O(N__7411),
            .I(N__7393));
    InMux I__1588 (
            .O(N__7410),
            .I(N__7393));
    InMux I__1587 (
            .O(N__7409),
            .I(N__7393));
    InMux I__1586 (
            .O(N__7408),
            .I(N__7390));
    CascadeMux I__1585 (
            .O(N__7407),
            .I(N__7385));
    LocalMux I__1584 (
            .O(N__7400),
            .I(N__7378));
    LocalMux I__1583 (
            .O(N__7393),
            .I(N__7375));
    LocalMux I__1582 (
            .O(N__7390),
            .I(N__7367));
    InMux I__1581 (
            .O(N__7389),
            .I(N__7362));
    InMux I__1580 (
            .O(N__7388),
            .I(N__7362));
    InMux I__1579 (
            .O(N__7385),
            .I(N__7355));
    InMux I__1578 (
            .O(N__7384),
            .I(N__7352));
    InMux I__1577 (
            .O(N__7383),
            .I(N__7345));
    InMux I__1576 (
            .O(N__7382),
            .I(N__7345));
    InMux I__1575 (
            .O(N__7381),
            .I(N__7345));
    Span4Mux_h I__1574 (
            .O(N__7378),
            .I(N__7342));
    Span4Mux_h I__1573 (
            .O(N__7375),
            .I(N__7339));
    InMux I__1572 (
            .O(N__7374),
            .I(N__7330));
    InMux I__1571 (
            .O(N__7373),
            .I(N__7330));
    InMux I__1570 (
            .O(N__7372),
            .I(N__7330));
    InMux I__1569 (
            .O(N__7371),
            .I(N__7330));
    InMux I__1568 (
            .O(N__7370),
            .I(N__7327));
    Span4Mux_h I__1567 (
            .O(N__7367),
            .I(N__7322));
    LocalMux I__1566 (
            .O(N__7362),
            .I(N__7322));
    InMux I__1565 (
            .O(N__7361),
            .I(N__7317));
    InMux I__1564 (
            .O(N__7360),
            .I(N__7317));
    InMux I__1563 (
            .O(N__7359),
            .I(N__7314));
    InMux I__1562 (
            .O(N__7358),
            .I(N__7311));
    LocalMux I__1561 (
            .O(N__7355),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1560 (
            .O(N__7352),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1559 (
            .O(N__7345),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1558 (
            .O(N__7342),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1557 (
            .O(N__7339),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1556 (
            .O(N__7330),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1555 (
            .O(N__7327),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1554 (
            .O(N__7322),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1553 (
            .O(N__7317),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1552 (
            .O(N__7314),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1551 (
            .O(N__7311),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__1550 (
            .O(N__7288),
            .I(N__7285));
    LocalMux I__1549 (
            .O(N__7285),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_0_3 ));
    CascadeMux I__1548 (
            .O(N__7282),
            .I(N__7279));
    InMux I__1547 (
            .O(N__7279),
            .I(N__7276));
    LocalMux I__1546 (
            .O(N__7276),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c6 ));
    InMux I__1545 (
            .O(N__7273),
            .I(N__7268));
    InMux I__1544 (
            .O(N__7272),
            .I(N__7263));
    InMux I__1543 (
            .O(N__7271),
            .I(N__7263));
    LocalMux I__1542 (
            .O(N__7268),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__1541 (
            .O(N__7263),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    CascadeMux I__1540 (
            .O(N__7258),
            .I(N__7254));
    InMux I__1539 (
            .O(N__7257),
            .I(N__7249));
    InMux I__1538 (
            .O(N__7254),
            .I(N__7249));
    LocalMux I__1537 (
            .O(N__7249),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__1536 (
            .O(N__7246),
            .I(N__7241));
    InMux I__1535 (
            .O(N__7245),
            .I(N__7231));
    InMux I__1534 (
            .O(N__7244),
            .I(N__7231));
    LocalMux I__1533 (
            .O(N__7241),
            .I(N__7228));
    InMux I__1532 (
            .O(N__7240),
            .I(N__7225));
    CascadeMux I__1531 (
            .O(N__7239),
            .I(N__7222));
    InMux I__1530 (
            .O(N__7238),
            .I(N__7218));
    InMux I__1529 (
            .O(N__7237),
            .I(N__7215));
    InMux I__1528 (
            .O(N__7236),
            .I(N__7212));
    LocalMux I__1527 (
            .O(N__7231),
            .I(N__7209));
    Span4Mux_v I__1526 (
            .O(N__7228),
            .I(N__7204));
    LocalMux I__1525 (
            .O(N__7225),
            .I(N__7204));
    InMux I__1524 (
            .O(N__7222),
            .I(N__7201));
    InMux I__1523 (
            .O(N__7221),
            .I(N__7198));
    LocalMux I__1522 (
            .O(N__7218),
            .I(\U712_CHIP_RAM.N_274 ));
    LocalMux I__1521 (
            .O(N__7215),
            .I(\U712_CHIP_RAM.N_274 ));
    LocalMux I__1520 (
            .O(N__7212),
            .I(\U712_CHIP_RAM.N_274 ));
    Odrv4 I__1519 (
            .O(N__7209),
            .I(\U712_CHIP_RAM.N_274 ));
    Odrv4 I__1518 (
            .O(N__7204),
            .I(\U712_CHIP_RAM.N_274 ));
    LocalMux I__1517 (
            .O(N__7201),
            .I(\U712_CHIP_RAM.N_274 ));
    LocalMux I__1516 (
            .O(N__7198),
            .I(\U712_CHIP_RAM.N_274 ));
    InMux I__1515 (
            .O(N__7183),
            .I(N__7180));
    LocalMux I__1514 (
            .O(N__7180),
            .I(N__7177));
    Sp12to4 I__1513 (
            .O(N__7177),
            .I(N__7174));
    Span12Mux_v I__1512 (
            .O(N__7174),
            .I(N__7171));
    Span12Mux_h I__1511 (
            .O(N__7171),
            .I(N__7168));
    Odrv12 I__1510 (
            .O(N__7168),
            .I(A_c_17));
    InMux I__1509 (
            .O(N__7165),
            .I(N__7162));
    LocalMux I__1508 (
            .O(N__7162),
            .I(N__7159));
    Odrv4 I__1507 (
            .O(N__7159),
            .I(\U712_CHIP_RAM.CMA_5_i_0_8 ));
    IoInMux I__1506 (
            .O(N__7156),
            .I(N__7153));
    LocalMux I__1505 (
            .O(N__7153),
            .I(N__7150));
    IoSpan4Mux I__1504 (
            .O(N__7150),
            .I(N__7147));
    Span4Mux_s0_h I__1503 (
            .O(N__7147),
            .I(N__7144));
    Sp12to4 I__1502 (
            .O(N__7144),
            .I(N__7141));
    Span12Mux_h I__1501 (
            .O(N__7141),
            .I(N__7138));
    Odrv12 I__1500 (
            .O(N__7138),
            .I(CMA_c_8));
    InMux I__1499 (
            .O(N__7135),
            .I(N__7132));
    LocalMux I__1498 (
            .O(N__7132),
            .I(\U712_CHIP_RAM.N_318 ));
    IoInMux I__1497 (
            .O(N__7129),
            .I(N__7126));
    LocalMux I__1496 (
            .O(N__7126),
            .I(N__7123));
    Span4Mux_s2_h I__1495 (
            .O(N__7123),
            .I(N__7120));
    Span4Mux_v I__1494 (
            .O(N__7120),
            .I(N__7117));
    Sp12to4 I__1493 (
            .O(N__7117),
            .I(N__7114));
    Span12Mux_h I__1492 (
            .O(N__7114),
            .I(N__7111));
    Odrv12 I__1491 (
            .O(N__7111),
            .I(CMA_c_7));
    CascadeMux I__1490 (
            .O(N__7108),
            .I(N__7104));
    InMux I__1489 (
            .O(N__7107),
            .I(N__7096));
    InMux I__1488 (
            .O(N__7104),
            .I(N__7089));
    InMux I__1487 (
            .O(N__7103),
            .I(N__7089));
    InMux I__1486 (
            .O(N__7102),
            .I(N__7084));
    InMux I__1485 (
            .O(N__7101),
            .I(N__7084));
    InMux I__1484 (
            .O(N__7100),
            .I(N__7081));
    InMux I__1483 (
            .O(N__7099),
            .I(N__7078));
    LocalMux I__1482 (
            .O(N__7096),
            .I(N__7070));
    InMux I__1481 (
            .O(N__7095),
            .I(N__7065));
    InMux I__1480 (
            .O(N__7094),
            .I(N__7065));
    LocalMux I__1479 (
            .O(N__7089),
            .I(N__7060));
    LocalMux I__1478 (
            .O(N__7084),
            .I(N__7060));
    LocalMux I__1477 (
            .O(N__7081),
            .I(N__7055));
    LocalMux I__1476 (
            .O(N__7078),
            .I(N__7055));
    InMux I__1475 (
            .O(N__7077),
            .I(N__7052));
    InMux I__1474 (
            .O(N__7076),
            .I(N__7045));
    InMux I__1473 (
            .O(N__7075),
            .I(N__7045));
    InMux I__1472 (
            .O(N__7074),
            .I(N__7045));
    InMux I__1471 (
            .O(N__7073),
            .I(N__7042));
    Span4Mux_v I__1470 (
            .O(N__7070),
            .I(N__7039));
    LocalMux I__1469 (
            .O(N__7065),
            .I(N__7028));
    Span4Mux_h I__1468 (
            .O(N__7060),
            .I(N__7028));
    Span4Mux_v I__1467 (
            .O(N__7055),
            .I(N__7028));
    LocalMux I__1466 (
            .O(N__7052),
            .I(N__7028));
    LocalMux I__1465 (
            .O(N__7045),
            .I(N__7028));
    LocalMux I__1464 (
            .O(N__7042),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1463 (
            .O(N__7039),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1462 (
            .O(N__7028),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    InMux I__1461 (
            .O(N__7021),
            .I(N__7018));
    LocalMux I__1460 (
            .O(N__7018),
            .I(N__7015));
    Odrv4 I__1459 (
            .O(N__7015),
            .I(\U712_CHIP_RAM.N_315 ));
    IoInMux I__1458 (
            .O(N__7012),
            .I(N__7009));
    LocalMux I__1457 (
            .O(N__7009),
            .I(N__7006));
    Span4Mux_s3_h I__1456 (
            .O(N__7006),
            .I(N__7003));
    Sp12to4 I__1455 (
            .O(N__7003),
            .I(N__7000));
    Span12Mux_s10_v I__1454 (
            .O(N__7000),
            .I(N__6997));
    Odrv12 I__1453 (
            .O(N__6997),
            .I(CMA_c_4));
    CEMux I__1452 (
            .O(N__6994),
            .I(N__6990));
    CEMux I__1451 (
            .O(N__6993),
            .I(N__6986));
    LocalMux I__1450 (
            .O(N__6990),
            .I(N__6982));
    CEMux I__1449 (
            .O(N__6989),
            .I(N__6979));
    LocalMux I__1448 (
            .O(N__6986),
            .I(N__6975));
    CEMux I__1447 (
            .O(N__6985),
            .I(N__6972));
    Span4Mux_v I__1446 (
            .O(N__6982),
            .I(N__6968));
    LocalMux I__1445 (
            .O(N__6979),
            .I(N__6965));
    CEMux I__1444 (
            .O(N__6978),
            .I(N__6962));
    Span4Mux_v I__1443 (
            .O(N__6975),
            .I(N__6957));
    LocalMux I__1442 (
            .O(N__6972),
            .I(N__6957));
    CEMux I__1441 (
            .O(N__6971),
            .I(N__6954));
    Span4Mux_h I__1440 (
            .O(N__6968),
            .I(N__6951));
    Span4Mux_v I__1439 (
            .O(N__6965),
            .I(N__6948));
    LocalMux I__1438 (
            .O(N__6962),
            .I(N__6945));
    Span4Mux_v I__1437 (
            .O(N__6957),
            .I(N__6942));
    LocalMux I__1436 (
            .O(N__6954),
            .I(N__6939));
    Odrv4 I__1435 (
            .O(N__6951),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    Odrv4 I__1434 (
            .O(N__6948),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    Odrv4 I__1433 (
            .O(N__6945),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    Odrv4 I__1432 (
            .O(N__6942),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    Odrv4 I__1431 (
            .O(N__6939),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    InMux I__1430 (
            .O(N__6928),
            .I(N__6924));
    InMux I__1429 (
            .O(N__6927),
            .I(N__6921));
    LocalMux I__1428 (
            .O(N__6924),
            .I(N__6918));
    LocalMux I__1427 (
            .O(N__6921),
            .I(N__6915));
    Span4Mux_v I__1426 (
            .O(N__6918),
            .I(N__6912));
    Sp12to4 I__1425 (
            .O(N__6915),
            .I(N__6909));
    Sp12to4 I__1424 (
            .O(N__6912),
            .I(N__6906));
    Span12Mux_v I__1423 (
            .O(N__6909),
            .I(N__6903));
    Span12Mux_h I__1422 (
            .O(N__6906),
            .I(N__6900));
    Span12Mux_h I__1421 (
            .O(N__6903),
            .I(N__6897));
    Span12Mux_v I__1420 (
            .O(N__6900),
            .I(N__6894));
    Odrv12 I__1419 (
            .O(N__6897),
            .I(AWEn_c));
    Odrv12 I__1418 (
            .O(N__6894),
            .I(AWEn_c));
    CascadeMux I__1417 (
            .O(N__6889),
            .I(N__6886));
    InMux I__1416 (
            .O(N__6886),
            .I(N__6883));
    LocalMux I__1415 (
            .O(N__6883),
            .I(N__6880));
    Span4Mux_v I__1414 (
            .O(N__6880),
            .I(N__6875));
    InMux I__1413 (
            .O(N__6879),
            .I(N__6871));
    InMux I__1412 (
            .O(N__6878),
            .I(N__6868));
    Span4Mux_v I__1411 (
            .O(N__6875),
            .I(N__6865));
    InMux I__1410 (
            .O(N__6874),
            .I(N__6862));
    LocalMux I__1409 (
            .O(N__6871),
            .I(N__6859));
    LocalMux I__1408 (
            .O(N__6868),
            .I(N__6856));
    Span4Mux_h I__1407 (
            .O(N__6865),
            .I(N__6853));
    LocalMux I__1406 (
            .O(N__6862),
            .I(N__6850));
    Span4Mux_v I__1405 (
            .O(N__6859),
            .I(N__6847));
    Span4Mux_v I__1404 (
            .O(N__6856),
            .I(N__6844));
    Sp12to4 I__1403 (
            .O(N__6853),
            .I(N__6835));
    Span12Mux_h I__1402 (
            .O(N__6850),
            .I(N__6835));
    Sp12to4 I__1401 (
            .O(N__6847),
            .I(N__6835));
    Sp12to4 I__1400 (
            .O(N__6844),
            .I(N__6835));
    Span12Mux_h I__1399 (
            .O(N__6835),
            .I(N__6832));
    Span12Mux_v I__1398 (
            .O(N__6832),
            .I(N__6829));
    Odrv12 I__1397 (
            .O(N__6829),
            .I(RnW_c));
    InMux I__1396 (
            .O(N__6826),
            .I(N__6817));
    InMux I__1395 (
            .O(N__6825),
            .I(N__6806));
    InMux I__1394 (
            .O(N__6824),
            .I(N__6801));
    InMux I__1393 (
            .O(N__6823),
            .I(N__6801));
    InMux I__1392 (
            .O(N__6822),
            .I(N__6798));
    InMux I__1391 (
            .O(N__6821),
            .I(N__6793));
    InMux I__1390 (
            .O(N__6820),
            .I(N__6793));
    LocalMux I__1389 (
            .O(N__6817),
            .I(N__6787));
    InMux I__1388 (
            .O(N__6816),
            .I(N__6782));
    InMux I__1387 (
            .O(N__6815),
            .I(N__6782));
    CascadeMux I__1386 (
            .O(N__6814),
            .I(N__6777));
    InMux I__1385 (
            .O(N__6813),
            .I(N__6770));
    InMux I__1384 (
            .O(N__6812),
            .I(N__6767));
    InMux I__1383 (
            .O(N__6811),
            .I(N__6764));
    InMux I__1382 (
            .O(N__6810),
            .I(N__6759));
    InMux I__1381 (
            .O(N__6809),
            .I(N__6759));
    LocalMux I__1380 (
            .O(N__6806),
            .I(N__6754));
    LocalMux I__1379 (
            .O(N__6801),
            .I(N__6754));
    LocalMux I__1378 (
            .O(N__6798),
            .I(N__6749));
    LocalMux I__1377 (
            .O(N__6793),
            .I(N__6749));
    InMux I__1376 (
            .O(N__6792),
            .I(N__6744));
    InMux I__1375 (
            .O(N__6791),
            .I(N__6740));
    InMux I__1374 (
            .O(N__6790),
            .I(N__6737));
    Span4Mux_h I__1373 (
            .O(N__6787),
            .I(N__6732));
    LocalMux I__1372 (
            .O(N__6782),
            .I(N__6732));
    InMux I__1371 (
            .O(N__6781),
            .I(N__6723));
    InMux I__1370 (
            .O(N__6780),
            .I(N__6723));
    InMux I__1369 (
            .O(N__6777),
            .I(N__6723));
    InMux I__1368 (
            .O(N__6776),
            .I(N__6723));
    CascadeMux I__1367 (
            .O(N__6775),
            .I(N__6720));
    CascadeMux I__1366 (
            .O(N__6774),
            .I(N__6717));
    CascadeMux I__1365 (
            .O(N__6773),
            .I(N__6714));
    LocalMux I__1364 (
            .O(N__6770),
            .I(N__6711));
    LocalMux I__1363 (
            .O(N__6767),
            .I(N__6706));
    LocalMux I__1362 (
            .O(N__6764),
            .I(N__6706));
    LocalMux I__1361 (
            .O(N__6759),
            .I(N__6701));
    Span4Mux_h I__1360 (
            .O(N__6754),
            .I(N__6701));
    Span4Mux_v I__1359 (
            .O(N__6749),
            .I(N__6698));
    InMux I__1358 (
            .O(N__6748),
            .I(N__6695));
    InMux I__1357 (
            .O(N__6747),
            .I(N__6692));
    LocalMux I__1356 (
            .O(N__6744),
            .I(N__6689));
    InMux I__1355 (
            .O(N__6743),
            .I(N__6686));
    LocalMux I__1354 (
            .O(N__6740),
            .I(N__6683));
    LocalMux I__1353 (
            .O(N__6737),
            .I(N__6676));
    Sp12to4 I__1352 (
            .O(N__6732),
            .I(N__6676));
    LocalMux I__1351 (
            .O(N__6723),
            .I(N__6676));
    InMux I__1350 (
            .O(N__6720),
            .I(N__6669));
    InMux I__1349 (
            .O(N__6717),
            .I(N__6669));
    InMux I__1348 (
            .O(N__6714),
            .I(N__6669));
    Span4Mux_v I__1347 (
            .O(N__6711),
            .I(N__6662));
    Span4Mux_v I__1346 (
            .O(N__6706),
            .I(N__6662));
    Span4Mux_v I__1345 (
            .O(N__6701),
            .I(N__6662));
    Odrv4 I__1344 (
            .O(N__6698),
            .I(CPU_CYCLEm));
    LocalMux I__1343 (
            .O(N__6695),
            .I(CPU_CYCLEm));
    LocalMux I__1342 (
            .O(N__6692),
            .I(CPU_CYCLEm));
    Odrv4 I__1341 (
            .O(N__6689),
            .I(CPU_CYCLEm));
    LocalMux I__1340 (
            .O(N__6686),
            .I(CPU_CYCLEm));
    Odrv4 I__1339 (
            .O(N__6683),
            .I(CPU_CYCLEm));
    Odrv12 I__1338 (
            .O(N__6676),
            .I(CPU_CYCLEm));
    LocalMux I__1337 (
            .O(N__6669),
            .I(CPU_CYCLEm));
    Odrv4 I__1336 (
            .O(N__6662),
            .I(CPU_CYCLEm));
    CEMux I__1335 (
            .O(N__6643),
            .I(N__6640));
    LocalMux I__1334 (
            .O(N__6640),
            .I(N__6637));
    Odrv4 I__1333 (
            .O(N__6637),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_0 ));
    InMux I__1332 (
            .O(N__6634),
            .I(N__6631));
    LocalMux I__1331 (
            .O(N__6631),
            .I(N__6626));
    CascadeMux I__1330 (
            .O(N__6630),
            .I(N__6621));
    InMux I__1329 (
            .O(N__6629),
            .I(N__6616));
    Span4Mux_v I__1328 (
            .O(N__6626),
            .I(N__6613));
    InMux I__1327 (
            .O(N__6625),
            .I(N__6608));
    InMux I__1326 (
            .O(N__6624),
            .I(N__6608));
    InMux I__1325 (
            .O(N__6621),
            .I(N__6601));
    InMux I__1324 (
            .O(N__6620),
            .I(N__6601));
    InMux I__1323 (
            .O(N__6619),
            .I(N__6601));
    LocalMux I__1322 (
            .O(N__6616),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1321 (
            .O(N__6613),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1320 (
            .O(N__6608),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1319 (
            .O(N__6601),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    CEMux I__1318 (
            .O(N__6592),
            .I(N__6589));
    LocalMux I__1317 (
            .O(N__6589),
            .I(N__6586));
    Span4Mux_v I__1316 (
            .O(N__6586),
            .I(N__6583));
    Span4Mux_h I__1315 (
            .O(N__6583),
            .I(N__6580));
    Odrv4 I__1314 (
            .O(N__6580),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_0 ));
    CEMux I__1313 (
            .O(N__6577),
            .I(N__6574));
    LocalMux I__1312 (
            .O(N__6574),
            .I(N__6571));
    Span4Mux_v I__1311 (
            .O(N__6571),
            .I(N__6568));
    Span4Mux_h I__1310 (
            .O(N__6568),
            .I(N__6565));
    Odrv4 I__1309 (
            .O(N__6565),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0 ));
    InMux I__1308 (
            .O(N__6562),
            .I(N__6559));
    LocalMux I__1307 (
            .O(N__6559),
            .I(N__6556));
    Odrv4 I__1306 (
            .O(N__6556),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_i_a2_1_0_a2_1_0 ));
    InMux I__1305 (
            .O(N__6553),
            .I(N__6550));
    LocalMux I__1304 (
            .O(N__6550),
            .I(\U712_CHIP_RAM.N_284 ));
    InMux I__1303 (
            .O(N__6547),
            .I(N__6542));
    InMux I__1302 (
            .O(N__6546),
            .I(N__6539));
    InMux I__1301 (
            .O(N__6545),
            .I(N__6536));
    LocalMux I__1300 (
            .O(N__6542),
            .I(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ));
    LocalMux I__1299 (
            .O(N__6539),
            .I(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ));
    LocalMux I__1298 (
            .O(N__6536),
            .I(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ));
    InMux I__1297 (
            .O(N__6529),
            .I(N__6525));
    InMux I__1296 (
            .O(N__6528),
            .I(N__6522));
    LocalMux I__1295 (
            .O(N__6525),
            .I(\U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ));
    LocalMux I__1294 (
            .O(N__6522),
            .I(\U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ));
    CascadeMux I__1293 (
            .O(N__6517),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER46_cascade_ ));
    CascadeMux I__1292 (
            .O(N__6514),
            .I(N__6511));
    InMux I__1291 (
            .O(N__6511),
            .I(N__6507));
    InMux I__1290 (
            .O(N__6510),
            .I(N__6504));
    LocalMux I__1289 (
            .O(N__6507),
            .I(N__6501));
    LocalMux I__1288 (
            .O(N__6504),
            .I(\U712_CHIP_RAM.N_420 ));
    Odrv4 I__1287 (
            .O(N__6501),
            .I(\U712_CHIP_RAM.N_420 ));
    InMux I__1286 (
            .O(N__6496),
            .I(N__6488));
    InMux I__1285 (
            .O(N__6495),
            .I(N__6479));
    InMux I__1284 (
            .O(N__6494),
            .I(N__6479));
    InMux I__1283 (
            .O(N__6493),
            .I(N__6479));
    InMux I__1282 (
            .O(N__6492),
            .I(N__6475));
    InMux I__1281 (
            .O(N__6491),
            .I(N__6472));
    LocalMux I__1280 (
            .O(N__6488),
            .I(N__6469));
    InMux I__1279 (
            .O(N__6487),
            .I(N__6464));
    InMux I__1278 (
            .O(N__6486),
            .I(N__6464));
    LocalMux I__1277 (
            .O(N__6479),
            .I(N__6461));
    InMux I__1276 (
            .O(N__6478),
            .I(N__6458));
    LocalMux I__1275 (
            .O(N__6475),
            .I(\U712_CHIP_RAM.N_282 ));
    LocalMux I__1274 (
            .O(N__6472),
            .I(\U712_CHIP_RAM.N_282 ));
    Odrv12 I__1273 (
            .O(N__6469),
            .I(\U712_CHIP_RAM.N_282 ));
    LocalMux I__1272 (
            .O(N__6464),
            .I(\U712_CHIP_RAM.N_282 ));
    Odrv4 I__1271 (
            .O(N__6461),
            .I(\U712_CHIP_RAM.N_282 ));
    LocalMux I__1270 (
            .O(N__6458),
            .I(\U712_CHIP_RAM.N_282 ));
    CascadeMux I__1269 (
            .O(N__6445),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_a5_i_0_cascade_ ));
    InMux I__1268 (
            .O(N__6442),
            .I(N__6439));
    LocalMux I__1267 (
            .O(N__6439),
            .I(\U712_CHIP_RAM.N_49 ));
    IoInMux I__1266 (
            .O(N__6436),
            .I(N__6433));
    LocalMux I__1265 (
            .O(N__6433),
            .I(N__6430));
    IoSpan4Mux I__1264 (
            .O(N__6430),
            .I(N__6427));
    IoSpan4Mux I__1263 (
            .O(N__6427),
            .I(N__6423));
    InMux I__1262 (
            .O(N__6426),
            .I(N__6420));
    Sp12to4 I__1261 (
            .O(N__6423),
            .I(N__6417));
    LocalMux I__1260 (
            .O(N__6420),
            .I(N__6414));
    Span12Mux_s9_v I__1259 (
            .O(N__6417),
            .I(N__6410));
    Span4Mux_v I__1258 (
            .O(N__6414),
            .I(N__6407));
    InMux I__1257 (
            .O(N__6413),
            .I(N__6404));
    Odrv12 I__1256 (
            .O(N__6410),
            .I(DBDIR_c));
    Odrv4 I__1255 (
            .O(N__6407),
            .I(DBDIR_c));
    LocalMux I__1254 (
            .O(N__6404),
            .I(DBDIR_c));
    IoInMux I__1253 (
            .O(N__6397),
            .I(N__6394));
    LocalMux I__1252 (
            .O(N__6394),
            .I(N__6391));
    Span12Mux_s8_h I__1251 (
            .O(N__6391),
            .I(N__6388));
    Span12Mux_v I__1250 (
            .O(N__6388),
            .I(N__6385));
    Odrv12 I__1249 (
            .O(N__6385),
            .I(N_218));
    IoInMux I__1248 (
            .O(N__6382),
            .I(N__6379));
    LocalMux I__1247 (
            .O(N__6379),
            .I(N__6376));
    Span4Mux_s0_v I__1246 (
            .O(N__6376),
            .I(N__6373));
    Span4Mux_v I__1245 (
            .O(N__6373),
            .I(N__6370));
    Span4Mux_v I__1244 (
            .O(N__6370),
            .I(N__6367));
    Span4Mux_h I__1243 (
            .O(N__6367),
            .I(N__6364));
    Odrv4 I__1242 (
            .O(N__6364),
            .I(RASn_c));
    InMux I__1241 (
            .O(N__6361),
            .I(N__6358));
    LocalMux I__1240 (
            .O(N__6358),
            .I(N__6355));
    Span4Mux_v I__1239 (
            .O(N__6355),
            .I(N__6352));
    Span4Mux_v I__1238 (
            .O(N__6352),
            .I(N__6349));
    Sp12to4 I__1237 (
            .O(N__6349),
            .I(N__6346));
    Span12Mux_h I__1236 (
            .O(N__6346),
            .I(N__6343));
    Odrv12 I__1235 (
            .O(N__6343),
            .I(A_c_18));
    CascadeMux I__1234 (
            .O(N__6340),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_7_cascade_ ));
    InMux I__1233 (
            .O(N__6337),
            .I(N__6334));
    LocalMux I__1232 (
            .O(N__6334),
            .I(N__6331));
    Span4Mux_v I__1231 (
            .O(N__6331),
            .I(N__6328));
    Span4Mux_v I__1230 (
            .O(N__6328),
            .I(N__6325));
    Sp12to4 I__1229 (
            .O(N__6325),
            .I(N__6322));
    Span12Mux_h I__1228 (
            .O(N__6322),
            .I(N__6319));
    Odrv12 I__1227 (
            .O(N__6319),
            .I(A_c_16));
    CascadeMux I__1226 (
            .O(N__6316),
            .I(\U712_CHIP_RAM.N_296_cascade_ ));
    InMux I__1225 (
            .O(N__6313),
            .I(N__6310));
    LocalMux I__1224 (
            .O(N__6310),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_a2_0_0_0 ));
    InMux I__1223 (
            .O(N__6307),
            .I(N__6304));
    LocalMux I__1222 (
            .O(N__6304),
            .I(N__6301));
    Odrv12 I__1221 (
            .O(N__6301),
            .I(\U712_CHIP_RAM.N_403 ));
    InMux I__1220 (
            .O(N__6298),
            .I(N__6289));
    InMux I__1219 (
            .O(N__6297),
            .I(N__6289));
    InMux I__1218 (
            .O(N__6296),
            .I(N__6289));
    LocalMux I__1217 (
            .O(N__6289),
            .I(\U712_CHIP_RAM.N_309 ));
    CascadeMux I__1216 (
            .O(N__6286),
            .I(N__6281));
    InMux I__1215 (
            .O(N__6285),
            .I(N__6278));
    InMux I__1214 (
            .O(N__6284),
            .I(N__6273));
    InMux I__1213 (
            .O(N__6281),
            .I(N__6273));
    LocalMux I__1212 (
            .O(N__6278),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ));
    LocalMux I__1211 (
            .O(N__6273),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ));
    InMux I__1210 (
            .O(N__6268),
            .I(N__6265));
    LocalMux I__1209 (
            .O(N__6265),
            .I(N__6262));
    Span4Mux_v I__1208 (
            .O(N__6262),
            .I(N__6259));
    Odrv4 I__1207 (
            .O(N__6259),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    CascadeMux I__1206 (
            .O(N__6256),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_1_cascade_ ));
    InMux I__1205 (
            .O(N__6253),
            .I(N__6250));
    LocalMux I__1204 (
            .O(N__6250),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0 ));
    InMux I__1203 (
            .O(N__6247),
            .I(N__6242));
    InMux I__1202 (
            .O(N__6246),
            .I(N__6237));
    InMux I__1201 (
            .O(N__6245),
            .I(N__6237));
    LocalMux I__1200 (
            .O(N__6242),
            .I(\U712_CHIP_RAM.N_285 ));
    LocalMux I__1199 (
            .O(N__6237),
            .I(\U712_CHIP_RAM.N_285 ));
    CascadeMux I__1198 (
            .O(N__6232),
            .I(N__6228));
    InMux I__1197 (
            .O(N__6231),
            .I(N__6225));
    InMux I__1196 (
            .O(N__6228),
            .I(N__6222));
    LocalMux I__1195 (
            .O(N__6225),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ));
    LocalMux I__1194 (
            .O(N__6222),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ));
    InMux I__1193 (
            .O(N__6217),
            .I(N__6214));
    LocalMux I__1192 (
            .O(N__6214),
            .I(N__6211));
    Span4Mux_h I__1191 (
            .O(N__6211),
            .I(N__6208));
    Odrv4 I__1190 (
            .O(N__6208),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    CascadeMux I__1189 (
            .O(N__6205),
            .I(\U712_CHIP_RAM.DMA_CYCLE_7_cascade_ ));
    InMux I__1188 (
            .O(N__6202),
            .I(N__6198));
    InMux I__1187 (
            .O(N__6201),
            .I(N__6195));
    LocalMux I__1186 (
            .O(N__6198),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0 ));
    LocalMux I__1185 (
            .O(N__6195),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0 ));
    IoInMux I__1184 (
            .O(N__6190),
            .I(N__6187));
    LocalMux I__1183 (
            .O(N__6187),
            .I(N__6184));
    IoSpan4Mux I__1182 (
            .O(N__6184),
            .I(N__6181));
    Span4Mux_s3_v I__1181 (
            .O(N__6181),
            .I(N__6174));
    InMux I__1180 (
            .O(N__6180),
            .I(N__6171));
    InMux I__1179 (
            .O(N__6179),
            .I(N__6168));
    InMux I__1178 (
            .O(N__6178),
            .I(N__6163));
    InMux I__1177 (
            .O(N__6177),
            .I(N__6163));
    Sp12to4 I__1176 (
            .O(N__6174),
            .I(N__6160));
    LocalMux I__1175 (
            .O(N__6171),
            .I(N__6155));
    LocalMux I__1174 (
            .O(N__6168),
            .I(N__6155));
    LocalMux I__1173 (
            .O(N__6163),
            .I(N__6152));
    Span12Mux_v I__1172 (
            .O(N__6160),
            .I(N__6148));
    Span4Mux_v I__1171 (
            .O(N__6155),
            .I(N__6145));
    Span4Mux_v I__1170 (
            .O(N__6152),
            .I(N__6142));
    InMux I__1169 (
            .O(N__6151),
            .I(N__6139));
    Odrv12 I__1168 (
            .O(N__6148),
            .I(DBENn_c));
    Odrv4 I__1167 (
            .O(N__6145),
            .I(DBENn_c));
    Odrv4 I__1166 (
            .O(N__6142),
            .I(DBENn_c));
    LocalMux I__1165 (
            .O(N__6139),
            .I(DBENn_c));
    InMux I__1164 (
            .O(N__6130),
            .I(N__6127));
    LocalMux I__1163 (
            .O(N__6127),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_0_a2_0_0 ));
    InMux I__1162 (
            .O(N__6124),
            .I(N__6121));
    LocalMux I__1161 (
            .O(N__6121),
            .I(N__6118));
    Odrv4 I__1160 (
            .O(N__6118),
            .I(\U712_CHIP_RAM.N_427 ));
    InMux I__1159 (
            .O(N__6115),
            .I(N__6112));
    LocalMux I__1158 (
            .O(N__6112),
            .I(\U712_CHIP_RAM.N_421 ));
    InMux I__1157 (
            .O(N__6109),
            .I(N__6106));
    LocalMux I__1156 (
            .O(N__6106),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1 ));
    CascadeMux I__1155 (
            .O(N__6103),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_ ));
    InMux I__1154 (
            .O(N__6100),
            .I(N__6096));
    CascadeMux I__1153 (
            .O(N__6099),
            .I(N__6093));
    LocalMux I__1152 (
            .O(N__6096),
            .I(N__6090));
    InMux I__1151 (
            .O(N__6093),
            .I(N__6087));
    Odrv4 I__1150 (
            .O(N__6090),
            .I(\U712_CHIP_RAM.N_296 ));
    LocalMux I__1149 (
            .O(N__6087),
            .I(\U712_CHIP_RAM.N_296 ));
    InMux I__1148 (
            .O(N__6082),
            .I(N__6079));
    LocalMux I__1147 (
            .O(N__6079),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_4 ));
    CascadeMux I__1146 (
            .O(N__6076),
            .I(N__6073));
    InMux I__1145 (
            .O(N__6073),
            .I(N__6070));
    LocalMux I__1144 (
            .O(N__6070),
            .I(N__6067));
    Span4Mux_v I__1143 (
            .O(N__6067),
            .I(N__6064));
    Sp12to4 I__1142 (
            .O(N__6064),
            .I(N__6061));
    Span12Mux_h I__1141 (
            .O(N__6061),
            .I(N__6058));
    Odrv12 I__1140 (
            .O(N__6058),
            .I(A_c_13));
    CascadeMux I__1139 (
            .O(N__6055),
            .I(\U712_CHIP_RAM.N_493_cascade_ ));
    CascadeMux I__1138 (
            .O(N__6052),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_cascade_ ));
    InMux I__1137 (
            .O(N__6049),
            .I(N__6046));
    LocalMux I__1136 (
            .O(N__6046),
            .I(\U712_CHIP_RAM.N_317 ));
    IoInMux I__1135 (
            .O(N__6043),
            .I(N__6040));
    LocalMux I__1134 (
            .O(N__6040),
            .I(N__6037));
    Span12Mux_s2_h I__1133 (
            .O(N__6037),
            .I(N__6034));
    Span12Mux_h I__1132 (
            .O(N__6034),
            .I(N__6031));
    Odrv12 I__1131 (
            .O(N__6031),
            .I(CMA_c_6));
    InMux I__1130 (
            .O(N__6028),
            .I(N__6025));
    LocalMux I__1129 (
            .O(N__6025),
            .I(N__6022));
    Span4Mux_v I__1128 (
            .O(N__6022),
            .I(N__6019));
    Sp12to4 I__1127 (
            .O(N__6019),
            .I(N__6016));
    Span12Mux_h I__1126 (
            .O(N__6016),
            .I(N__6013));
    Span12Mux_v I__1125 (
            .O(N__6013),
            .I(N__6010));
    Odrv12 I__1124 (
            .O(N__6010),
            .I(A_c_19));
    CascadeMux I__1123 (
            .O(N__6007),
            .I(\U712_CHIP_RAM.CMA_5_i_0_8_cascade_ ));
    IoInMux I__1122 (
            .O(N__6004),
            .I(N__6001));
    LocalMux I__1121 (
            .O(N__6001),
            .I(N__5998));
    IoSpan4Mux I__1120 (
            .O(N__5998),
            .I(N__5995));
    Span4Mux_s3_h I__1119 (
            .O(N__5995),
            .I(N__5992));
    Sp12to4 I__1118 (
            .O(N__5992),
            .I(N__5989));
    Span12Mux_h I__1117 (
            .O(N__5989),
            .I(N__5986));
    Odrv12 I__1116 (
            .O(N__5986),
            .I(CMA_c_9));
    SRMux I__1115 (
            .O(N__5983),
            .I(N__5980));
    LocalMux I__1114 (
            .O(N__5980),
            .I(N__5976));
    InMux I__1113 (
            .O(N__5979),
            .I(N__5973));
    Span4Mux_v I__1112 (
            .O(N__5976),
            .I(N__5970));
    LocalMux I__1111 (
            .O(N__5973),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    Odrv4 I__1110 (
            .O(N__5970),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    CascadeMux I__1109 (
            .O(N__5965),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_cascade_ ));
    InMux I__1108 (
            .O(N__5962),
            .I(N__5959));
    LocalMux I__1107 (
            .O(N__5959),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_0 ));
    InMux I__1106 (
            .O(N__5956),
            .I(N__5952));
    InMux I__1105 (
            .O(N__5955),
            .I(N__5949));
    LocalMux I__1104 (
            .O(N__5952),
            .I(CPU_TACKm));
    LocalMux I__1103 (
            .O(N__5949),
            .I(CPU_TACKm));
    InMux I__1102 (
            .O(N__5944),
            .I(N__5941));
    LocalMux I__1101 (
            .O(N__5941),
            .I(N__5936));
    InMux I__1100 (
            .O(N__5940),
            .I(N__5933));
    InMux I__1099 (
            .O(N__5939),
            .I(N__5930));
    Odrv12 I__1098 (
            .O(N__5936),
            .I(\U712_REG_SM.DS_ENZ0 ));
    LocalMux I__1097 (
            .O(N__5933),
            .I(\U712_REG_SM.DS_ENZ0 ));
    LocalMux I__1096 (
            .O(N__5930),
            .I(\U712_REG_SM.DS_ENZ0 ));
    InMux I__1095 (
            .O(N__5923),
            .I(N__5920));
    LocalMux I__1094 (
            .O(N__5920),
            .I(N__5916));
    InMux I__1093 (
            .O(N__5919),
            .I(N__5913));
    Odrv12 I__1092 (
            .O(N__5916),
            .I(\U712_REG_SM.LDS_OUTZ0 ));
    LocalMux I__1091 (
            .O(N__5913),
            .I(\U712_REG_SM.LDS_OUTZ0 ));
    IoInMux I__1090 (
            .O(N__5908),
            .I(N__5905));
    LocalMux I__1089 (
            .O(N__5905),
            .I(N__5902));
    IoSpan4Mux I__1088 (
            .O(N__5902),
            .I(N__5899));
    Span4Mux_s2_v I__1087 (
            .O(N__5899),
            .I(N__5896));
    Sp12to4 I__1086 (
            .O(N__5896),
            .I(N__5893));
    Span12Mux_v I__1085 (
            .O(N__5893),
            .I(N__5890));
    Odrv12 I__1084 (
            .O(N__5890),
            .I(U712_REG_SM_un1_LDSn_i));
    InMux I__1083 (
            .O(N__5887),
            .I(N__5884));
    LocalMux I__1082 (
            .O(N__5884),
            .I(\U712_CHIP_RAM.N_311 ));
    IoInMux I__1081 (
            .O(N__5881),
            .I(N__5878));
    LocalMux I__1080 (
            .O(N__5878),
            .I(N__5875));
    Span4Mux_s1_v I__1079 (
            .O(N__5875),
            .I(N__5872));
    Span4Mux_v I__1078 (
            .O(N__5872),
            .I(N__5869));
    Span4Mux_v I__1077 (
            .O(N__5869),
            .I(N__5866));
    Odrv4 I__1076 (
            .O(N__5866),
            .I(CMA_c_0));
    InMux I__1075 (
            .O(N__5863),
            .I(N__5860));
    LocalMux I__1074 (
            .O(N__5860),
            .I(\U712_CHIP_RAM.N_312 ));
    IoInMux I__1073 (
            .O(N__5857),
            .I(N__5854));
    LocalMux I__1072 (
            .O(N__5854),
            .I(N__5851));
    Span4Mux_s2_v I__1071 (
            .O(N__5851),
            .I(N__5848));
    Span4Mux_v I__1070 (
            .O(N__5848),
            .I(N__5845));
    Span4Mux_v I__1069 (
            .O(N__5845),
            .I(N__5842));
    Odrv4 I__1068 (
            .O(N__5842),
            .I(CMA_c_1));
    InMux I__1067 (
            .O(N__5839),
            .I(N__5836));
    LocalMux I__1066 (
            .O(N__5836),
            .I(\U712_CHIP_RAM.N_316 ));
    IoInMux I__1065 (
            .O(N__5833),
            .I(N__5830));
    LocalMux I__1064 (
            .O(N__5830),
            .I(N__5827));
    Span4Mux_s2_h I__1063 (
            .O(N__5827),
            .I(N__5824));
    Span4Mux_v I__1062 (
            .O(N__5824),
            .I(N__5821));
    Sp12to4 I__1061 (
            .O(N__5821),
            .I(N__5818));
    Span12Mux_h I__1060 (
            .O(N__5818),
            .I(N__5815));
    Odrv12 I__1059 (
            .O(N__5815),
            .I(CMA_c_5));
    CascadeMux I__1058 (
            .O(N__5812),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_cascade_ ));
    InMux I__1057 (
            .O(N__5809),
            .I(N__5806));
    LocalMux I__1056 (
            .O(N__5806),
            .I(N__5803));
    Span12Mux_v I__1055 (
            .O(N__5803),
            .I(N__5800));
    Span12Mux_h I__1054 (
            .O(N__5800),
            .I(N__5797));
    Odrv12 I__1053 (
            .O(N__5797),
            .I(A_c_6));
    InMux I__1052 (
            .O(N__5794),
            .I(N__5790));
    InMux I__1051 (
            .O(N__5793),
            .I(N__5787));
    LocalMux I__1050 (
            .O(N__5790),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__1049 (
            .O(N__5787),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    CascadeMux I__1048 (
            .O(N__5782),
            .I(N__5779));
    InMux I__1047 (
            .O(N__5779),
            .I(N__5776));
    LocalMux I__1046 (
            .O(N__5776),
            .I(N__5772));
    InMux I__1045 (
            .O(N__5775),
            .I(N__5768));
    Span4Mux_v I__1044 (
            .O(N__5772),
            .I(N__5765));
    InMux I__1043 (
            .O(N__5771),
            .I(N__5762));
    LocalMux I__1042 (
            .O(N__5768),
            .I(U712_REG_SM_DBR_SYNC_0));
    Odrv4 I__1041 (
            .O(N__5765),
            .I(U712_REG_SM_DBR_SYNC_0));
    LocalMux I__1040 (
            .O(N__5762),
            .I(U712_REG_SM_DBR_SYNC_0));
    InMux I__1039 (
            .O(N__5755),
            .I(N__5752));
    LocalMux I__1038 (
            .O(N__5752),
            .I(N__5749));
    Span4Mux_h I__1037 (
            .O(N__5749),
            .I(N__5745));
    InMux I__1036 (
            .O(N__5748),
            .I(N__5742));
    Odrv4 I__1035 (
            .O(N__5745),
            .I(U712_REG_SM_DBR_SYNC_1));
    LocalMux I__1034 (
            .O(N__5742),
            .I(U712_REG_SM_DBR_SYNC_1));
    InMux I__1033 (
            .O(N__5737),
            .I(N__5734));
    LocalMux I__1032 (
            .O(N__5734),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_3_1 ));
    CascadeMux I__1031 (
            .O(N__5731),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_2_1_cascade_ ));
    CascadeMux I__1030 (
            .O(N__5728),
            .I(\U712_CHIP_RAM.N_421_cascade_ ));
    CascadeMux I__1029 (
            .O(N__5725),
            .I(\U712_CHIP_RAM.N_293_cascade_ ));
    CascadeMux I__1028 (
            .O(N__5722),
            .I(\U712_CHIP_RAM.N_309_cascade_ ));
    InMux I__1027 (
            .O(N__5719),
            .I(N__5716));
    LocalMux I__1026 (
            .O(N__5716),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_0_a2_0_a2_0 ));
    InMux I__1025 (
            .O(N__5713),
            .I(N__5710));
    LocalMux I__1024 (
            .O(N__5710),
            .I(N__5707));
    Span4Mux_v I__1023 (
            .O(N__5707),
            .I(N__5704));
    Sp12to4 I__1022 (
            .O(N__5704),
            .I(N__5701));
    Span12Mux_v I__1021 (
            .O(N__5701),
            .I(N__5698));
    Span12Mux_h I__1020 (
            .O(N__5698),
            .I(N__5695));
    Odrv12 I__1019 (
            .O(N__5695),
            .I(DBRn_c));
    CascadeMux I__1018 (
            .O(N__5692),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_0_cascade_ ));
    CascadeMux I__1017 (
            .O(N__5689),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_2_cascade_ ));
    InMux I__1016 (
            .O(N__5686),
            .I(N__5680));
    InMux I__1015 (
            .O(N__5685),
            .I(N__5680));
    LocalMux I__1014 (
            .O(N__5680),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__1013 (
            .O(N__5677),
            .I(N__5672));
    InMux I__1012 (
            .O(N__5676),
            .I(N__5667));
    InMux I__1011 (
            .O(N__5675),
            .I(N__5667));
    LocalMux I__1010 (
            .O(N__5672),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    LocalMux I__1009 (
            .O(N__5667),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    CascadeMux I__1008 (
            .O(N__5662),
            .I(\U712_CHIP_RAM.N_314_cascade_ ));
    IoInMux I__1007 (
            .O(N__5659),
            .I(N__5656));
    LocalMux I__1006 (
            .O(N__5656),
            .I(N__5653));
    IoSpan4Mux I__1005 (
            .O(N__5653),
            .I(N__5650));
    Span4Mux_s1_h I__1004 (
            .O(N__5650),
            .I(N__5647));
    Sp12to4 I__1003 (
            .O(N__5647),
            .I(N__5644));
    Span12Mux_h I__1002 (
            .O(N__5644),
            .I(N__5641));
    Odrv12 I__1001 (
            .O(N__5641),
            .I(CMA_c_3));
    InMux I__1000 (
            .O(N__5638),
            .I(N__5635));
    LocalMux I__999 (
            .O(N__5635),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__998 (
            .O(N__5632),
            .I(N__5629));
    LocalMux I__997 (
            .O(N__5629),
            .I(N__5626));
    Odrv4 I__996 (
            .O(N__5626),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_5 ));
    InMux I__995 (
            .O(N__5623),
            .I(N__5619));
    InMux I__994 (
            .O(N__5622),
            .I(N__5616));
    LocalMux I__993 (
            .O(N__5619),
            .I(N__5611));
    LocalMux I__992 (
            .O(N__5616),
            .I(N__5611));
    Span4Mux_v I__991 (
            .O(N__5611),
            .I(N__5608));
    Span4Mux_v I__990 (
            .O(N__5608),
            .I(N__5605));
    Sp12to4 I__989 (
            .O(N__5605),
            .I(N__5602));
    Span12Mux_h I__988 (
            .O(N__5602),
            .I(N__5599));
    Odrv12 I__987 (
            .O(N__5599),
            .I(DRA_c_6));
    InMux I__986 (
            .O(N__5596),
            .I(N__5593));
    LocalMux I__985 (
            .O(N__5593),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__984 (
            .O(N__5590),
            .I(N__5587));
    LocalMux I__983 (
            .O(N__5587),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__982 (
            .O(N__5584),
            .I(N__5581));
    LocalMux I__981 (
            .O(N__5581),
            .I(N__5577));
    InMux I__980 (
            .O(N__5580),
            .I(N__5574));
    Span4Mux_v I__979 (
            .O(N__5577),
            .I(N__5571));
    LocalMux I__978 (
            .O(N__5574),
            .I(N__5568));
    Span4Mux_v I__977 (
            .O(N__5571),
            .I(N__5565));
    Sp12to4 I__976 (
            .O(N__5568),
            .I(N__5562));
    Sp12to4 I__975 (
            .O(N__5565),
            .I(N__5557));
    Span12Mux_v I__974 (
            .O(N__5562),
            .I(N__5557));
    Span12Mux_h I__973 (
            .O(N__5557),
            .I(N__5554));
    Odrv12 I__972 (
            .O(N__5554),
            .I(DRA_c_5));
    InMux I__971 (
            .O(N__5551),
            .I(N__5548));
    LocalMux I__970 (
            .O(N__5548),
            .I(N__5545));
    Odrv4 I__969 (
            .O(N__5545),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__968 (
            .O(N__5542),
            .I(N__5539));
    LocalMux I__967 (
            .O(N__5539),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__966 (
            .O(N__5536),
            .I(N__5533));
    LocalMux I__965 (
            .O(N__5533),
            .I(N__5530));
    Sp12to4 I__964 (
            .O(N__5530),
            .I(N__5527));
    Span12Mux_v I__963 (
            .O(N__5527),
            .I(N__5524));
    Span12Mux_h I__962 (
            .O(N__5524),
            .I(N__5521));
    Odrv12 I__961 (
            .O(N__5521),
            .I(A_c_8));
    CascadeMux I__960 (
            .O(N__5518),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_6_cascade_ ));
    InMux I__959 (
            .O(N__5515),
            .I(N__5512));
    LocalMux I__958 (
            .O(N__5512),
            .I(N__5509));
    Span4Mux_v I__957 (
            .O(N__5509),
            .I(N__5506));
    Span4Mux_v I__956 (
            .O(N__5506),
            .I(N__5503));
    Sp12to4 I__955 (
            .O(N__5503),
            .I(N__5500));
    Span12Mux_h I__954 (
            .O(N__5500),
            .I(N__5497));
    Odrv12 I__953 (
            .O(N__5497),
            .I(A_c_15));
    InMux I__952 (
            .O(N__5494),
            .I(N__5491));
    LocalMux I__951 (
            .O(N__5491),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__950 (
            .O(N__5488),
            .I(N__5485));
    LocalMux I__949 (
            .O(N__5485),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__948 (
            .O(N__5482),
            .I(N__5479));
    LocalMux I__947 (
            .O(N__5479),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__946 (
            .O(N__5476),
            .I(N__5473));
    LocalMux I__945 (
            .O(N__5473),
            .I(N__5470));
    Span4Mux_v I__944 (
            .O(N__5470),
            .I(N__5467));
    Span4Mux_v I__943 (
            .O(N__5467),
            .I(N__5464));
    Sp12to4 I__942 (
            .O(N__5464),
            .I(N__5461));
    Span12Mux_h I__941 (
            .O(N__5461),
            .I(N__5458));
    Odrv12 I__940 (
            .O(N__5458),
            .I(A_c_9));
    InMux I__939 (
            .O(N__5455),
            .I(N__5452));
    LocalMux I__938 (
            .O(N__5452),
            .I(N__5449));
    Span4Mux_h I__937 (
            .O(N__5449),
            .I(N__5446));
    Span4Mux_v I__936 (
            .O(N__5446),
            .I(N__5443));
    Sp12to4 I__935 (
            .O(N__5443),
            .I(N__5440));
    Span12Mux_h I__934 (
            .O(N__5440),
            .I(N__5437));
    Span12Mux_v I__933 (
            .O(N__5437),
            .I(N__5434));
    Odrv12 I__932 (
            .O(N__5434),
            .I(A_c_2));
    CascadeMux I__931 (
            .O(N__5431),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_0_cascade_ ));
    InMux I__930 (
            .O(N__5428),
            .I(N__5425));
    LocalMux I__929 (
            .O(N__5425),
            .I(N__5422));
    Odrv4 I__928 (
            .O(N__5422),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__927 (
            .O(N__5419),
            .I(N__5416));
    LocalMux I__926 (
            .O(N__5416),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__925 (
            .O(N__5413),
            .I(N__5410));
    LocalMux I__924 (
            .O(N__5410),
            .I(N__5407));
    Span4Mux_v I__923 (
            .O(N__5407),
            .I(N__5404));
    Sp12to4 I__922 (
            .O(N__5404),
            .I(N__5401));
    Span12Mux_h I__921 (
            .O(N__5401),
            .I(N__5398));
    Odrv12 I__920 (
            .O(N__5398),
            .I(A_c_10));
    InMux I__919 (
            .O(N__5395),
            .I(N__5392));
    LocalMux I__918 (
            .O(N__5392),
            .I(N__5389));
    Span4Mux_v I__917 (
            .O(N__5389),
            .I(N__5386));
    Sp12to4 I__916 (
            .O(N__5386),
            .I(N__5383));
    Span12Mux_h I__915 (
            .O(N__5383),
            .I(N__5380));
    Span12Mux_v I__914 (
            .O(N__5380),
            .I(N__5377));
    Odrv12 I__913 (
            .O(N__5377),
            .I(A_c_3));
    CascadeMux I__912 (
            .O(N__5374),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_1_cascade_ ));
    IoInMux I__911 (
            .O(N__5371),
            .I(N__5368));
    LocalMux I__910 (
            .O(N__5368),
            .I(N__5365));
    Span4Mux_s2_v I__909 (
            .O(N__5365),
            .I(N__5362));
    Span4Mux_v I__908 (
            .O(N__5362),
            .I(N__5359));
    Span4Mux_v I__907 (
            .O(N__5359),
            .I(N__5356));
    Span4Mux_h I__906 (
            .O(N__5356),
            .I(N__5353));
    Odrv4 I__905 (
            .O(N__5353),
            .I(CMA_c_10));
    InMux I__904 (
            .O(N__5350),
            .I(N__5347));
    LocalMux I__903 (
            .O(N__5347),
            .I(N__5344));
    Odrv4 I__902 (
            .O(N__5344),
            .I(\U712_CHIP_RAM.N_313 ));
    IoInMux I__901 (
            .O(N__5341),
            .I(N__5338));
    LocalMux I__900 (
            .O(N__5338),
            .I(N__5335));
    IoSpan4Mux I__899 (
            .O(N__5335),
            .I(N__5332));
    Span4Mux_s3_v I__898 (
            .O(N__5332),
            .I(N__5329));
    Span4Mux_v I__897 (
            .O(N__5329),
            .I(N__5326));
    Odrv4 I__896 (
            .O(N__5326),
            .I(CMA_c_2));
    InMux I__895 (
            .O(N__5323),
            .I(N__5320));
    LocalMux I__894 (
            .O(N__5320),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__893 (
            .O(N__5317),
            .I(N__5314));
    LocalMux I__892 (
            .O(N__5314),
            .I(N__5311));
    Span4Mux_v I__891 (
            .O(N__5311),
            .I(N__5308));
    Sp12to4 I__890 (
            .O(N__5308),
            .I(N__5305));
    Span12Mux_h I__889 (
            .O(N__5305),
            .I(N__5302));
    Span12Mux_v I__888 (
            .O(N__5302),
            .I(N__5299));
    Odrv12 I__887 (
            .O(N__5299),
            .I(A_c_5));
    CascadeMux I__886 (
            .O(N__5296),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_3_cascade_ ));
    InMux I__885 (
            .O(N__5293),
            .I(N__5290));
    LocalMux I__884 (
            .O(N__5290),
            .I(N__5287));
    Span4Mux_v I__883 (
            .O(N__5287),
            .I(N__5284));
    Sp12to4 I__882 (
            .O(N__5284),
            .I(N__5281));
    Span12Mux_h I__881 (
            .O(N__5281),
            .I(N__5278));
    Odrv12 I__880 (
            .O(N__5278),
            .I(A_c_12));
    CascadeMux I__879 (
            .O(N__5275),
            .I(N__5272));
    InMux I__878 (
            .O(N__5272),
            .I(N__5269));
    LocalMux I__877 (
            .O(N__5269),
            .I(N__5266));
    Span4Mux_v I__876 (
            .O(N__5266),
            .I(N__5263));
    Odrv4 I__875 (
            .O(N__5263),
            .I(\U712_BYTE_ENABLE.N_392 ));
    InMux I__874 (
            .O(N__5260),
            .I(N__5257));
    LocalMux I__873 (
            .O(N__5257),
            .I(N__5254));
    Span4Mux_v I__872 (
            .O(N__5254),
            .I(N__5251));
    Odrv4 I__871 (
            .O(N__5251),
            .I(\U712_BYTE_ENABLE.N_388 ));
    InMux I__870 (
            .O(N__5248),
            .I(N__5243));
    InMux I__869 (
            .O(N__5247),
            .I(N__5240));
    InMux I__868 (
            .O(N__5246),
            .I(N__5237));
    LocalMux I__867 (
            .O(N__5243),
            .I(N__5234));
    LocalMux I__866 (
            .O(N__5240),
            .I(N__5229));
    LocalMux I__865 (
            .O(N__5237),
            .I(N__5229));
    Span4Mux_v I__864 (
            .O(N__5234),
            .I(N__5226));
    Span12Mux_v I__863 (
            .O(N__5229),
            .I(N__5223));
    Sp12to4 I__862 (
            .O(N__5226),
            .I(N__5220));
    Span12Mux_h I__861 (
            .O(N__5223),
            .I(N__5217));
    Span12Mux_h I__860 (
            .O(N__5220),
            .I(N__5214));
    Span12Mux_v I__859 (
            .O(N__5217),
            .I(N__5211));
    Span12Mux_v I__858 (
            .O(N__5214),
            .I(N__5208));
    Odrv12 I__857 (
            .O(N__5211),
            .I(CASLn_c));
    Odrv12 I__856 (
            .O(N__5208),
            .I(CASLn_c));
    CascadeMux I__855 (
            .O(N__5203),
            .I(N__5199));
    InMux I__854 (
            .O(N__5202),
            .I(N__5191));
    InMux I__853 (
            .O(N__5199),
            .I(N__5191));
    InMux I__852 (
            .O(N__5198),
            .I(N__5191));
    LocalMux I__851 (
            .O(N__5191),
            .I(N__5188));
    Span12Mux_v I__850 (
            .O(N__5188),
            .I(N__5185));
    Span12Mux_h I__849 (
            .O(N__5185),
            .I(N__5182));
    Span12Mux_v I__848 (
            .O(N__5182),
            .I(N__5179));
    Odrv12 I__847 (
            .O(N__5179),
            .I(CASUn_c));
    InMux I__846 (
            .O(N__5176),
            .I(N__5173));
    LocalMux I__845 (
            .O(N__5173),
            .I(N__5170));
    Span4Mux_v I__844 (
            .O(N__5170),
            .I(N__5167));
    Sp12to4 I__843 (
            .O(N__5167),
            .I(N__5163));
    IoInMux I__842 (
            .O(N__5166),
            .I(N__5160));
    Span12Mux_h I__841 (
            .O(N__5163),
            .I(N__5157));
    LocalMux I__840 (
            .O(N__5160),
            .I(N__5154));
    Span12Mux_v I__839 (
            .O(N__5157),
            .I(N__5151));
    IoSpan4Mux I__838 (
            .O(N__5154),
            .I(N__5148));
    Odrv12 I__837 (
            .O(N__5151),
            .I(RAMENn_c));
    Odrv4 I__836 (
            .O(N__5148),
            .I(RAMENn_c));
    CascadeMux I__835 (
            .O(N__5143),
            .I(N__5140));
    InMux I__834 (
            .O(N__5140),
            .I(N__5136));
    InMux I__833 (
            .O(N__5139),
            .I(N__5133));
    LocalMux I__832 (
            .O(N__5136),
            .I(N__5130));
    LocalMux I__831 (
            .O(N__5133),
            .I(N__5127));
    Span4Mux_v I__830 (
            .O(N__5130),
            .I(N__5124));
    Span4Mux_v I__829 (
            .O(N__5127),
            .I(N__5121));
    Sp12to4 I__828 (
            .O(N__5124),
            .I(N__5116));
    Sp12to4 I__827 (
            .O(N__5121),
            .I(N__5116));
    Span12Mux_h I__826 (
            .O(N__5116),
            .I(N__5113));
    Span12Mux_v I__825 (
            .O(N__5113),
            .I(N__5110));
    Odrv12 I__824 (
            .O(N__5110),
            .I(TSn_c));
    InMux I__823 (
            .O(N__5107),
            .I(N__5103));
    InMux I__822 (
            .O(N__5106),
            .I(N__5100));
    LocalMux I__821 (
            .O(N__5103),
            .I(REG_TACK));
    LocalMux I__820 (
            .O(N__5100),
            .I(REG_TACK));
    CascadeMux I__819 (
            .O(N__5095),
            .I(N__5091));
    InMux I__818 (
            .O(N__5094),
            .I(N__5088));
    InMux I__817 (
            .O(N__5091),
            .I(N__5084));
    LocalMux I__816 (
            .O(N__5088),
            .I(N__5081));
    InMux I__815 (
            .O(N__5087),
            .I(N__5078));
    LocalMux I__814 (
            .O(N__5084),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    Odrv4 I__813 (
            .O(N__5081),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__812 (
            .O(N__5078),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    InMux I__811 (
            .O(N__5071),
            .I(N__5065));
    InMux I__810 (
            .O(N__5070),
            .I(N__5065));
    LocalMux I__809 (
            .O(N__5065),
            .I(N__5061));
    InMux I__808 (
            .O(N__5064),
            .I(N__5057));
    Span4Mux_v I__807 (
            .O(N__5061),
            .I(N__5054));
    InMux I__806 (
            .O(N__5060),
            .I(N__5051));
    LocalMux I__805 (
            .O(N__5057),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    Odrv4 I__804 (
            .O(N__5054),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    LocalMux I__803 (
            .O(N__5051),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    InMux I__802 (
            .O(N__5044),
            .I(N__5041));
    LocalMux I__801 (
            .O(N__5041),
            .I(N__5038));
    Span4Mux_v I__800 (
            .O(N__5038),
            .I(N__5035));
    Span4Mux_v I__799 (
            .O(N__5035),
            .I(N__5032));
    Odrv4 I__798 (
            .O(N__5032),
            .I(TACK_EN_i_ess));
    CEMux I__797 (
            .O(N__5029),
            .I(N__5026));
    LocalMux I__796 (
            .O(N__5026),
            .I(\U712_CYCLE_TERM.N_305_i_0_en_0 ));
    IoInMux I__795 (
            .O(N__5023),
            .I(N__5020));
    LocalMux I__794 (
            .O(N__5020),
            .I(N__5017));
    Odrv12 I__793 (
            .O(N__5017),
            .I(RESETn_c_i));
    InMux I__792 (
            .O(N__5014),
            .I(N__5011));
    LocalMux I__791 (
            .O(N__5011),
            .I(N__5008));
    Span4Mux_v I__790 (
            .O(N__5008),
            .I(N__5005));
    Sp12to4 I__789 (
            .O(N__5005),
            .I(N__5002));
    Span12Mux_h I__788 (
            .O(N__5002),
            .I(N__4999));
    Span12Mux_v I__787 (
            .O(N__4999),
            .I(N__4996));
    Odrv12 I__786 (
            .O(N__4996),
            .I(A_c_7));
    CascadeMux I__785 (
            .O(N__4993),
            .I(N__4990));
    InMux I__784 (
            .O(N__4990),
            .I(N__4987));
    LocalMux I__783 (
            .O(N__4987),
            .I(N__4984));
    Span4Mux_v I__782 (
            .O(N__4984),
            .I(N__4981));
    Sp12to4 I__781 (
            .O(N__4981),
            .I(N__4978));
    Span12Mux_h I__780 (
            .O(N__4978),
            .I(N__4975));
    Odrv12 I__779 (
            .O(N__4975),
            .I(A_c_14));
    InMux I__778 (
            .O(N__4972),
            .I(N__4968));
    InMux I__777 (
            .O(N__4971),
            .I(N__4965));
    LocalMux I__776 (
            .O(N__4968),
            .I(N__4962));
    LocalMux I__775 (
            .O(N__4965),
            .I(N__4959));
    Span4Mux_v I__774 (
            .O(N__4962),
            .I(N__4954));
    Span4Mux_v I__773 (
            .O(N__4959),
            .I(N__4954));
    Sp12to4 I__772 (
            .O(N__4954),
            .I(N__4951));
    Span12Mux_h I__771 (
            .O(N__4951),
            .I(N__4948));
    Span12Mux_v I__770 (
            .O(N__4948),
            .I(N__4945));
    Odrv12 I__769 (
            .O(N__4945),
            .I(DRA_c_2));
    InMux I__768 (
            .O(N__4942),
            .I(N__4939));
    LocalMux I__767 (
            .O(N__4939),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__766 (
            .O(N__4936),
            .I(N__4932));
    InMux I__765 (
            .O(N__4935),
            .I(N__4929));
    LocalMux I__764 (
            .O(N__4932),
            .I(N__4924));
    LocalMux I__763 (
            .O(N__4929),
            .I(N__4924));
    Span12Mux_v I__762 (
            .O(N__4924),
            .I(N__4921));
    Span12Mux_h I__761 (
            .O(N__4921),
            .I(N__4918));
    Odrv12 I__760 (
            .O(N__4918),
            .I(DRA_c_4));
    CascadeMux I__759 (
            .O(N__4915),
            .I(\U712_CHIP_RAM.N_341_cascade_ ));
    CascadeMux I__758 (
            .O(N__4912),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_1_1_cascade_ ));
    InMux I__757 (
            .O(N__4909),
            .I(N__4905));
    InMux I__756 (
            .O(N__4908),
            .I(N__4902));
    LocalMux I__755 (
            .O(N__4905),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    LocalMux I__754 (
            .O(N__4902),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    InMux I__753 (
            .O(N__4897),
            .I(N__4893));
    InMux I__752 (
            .O(N__4896),
            .I(N__4890));
    LocalMux I__751 (
            .O(N__4893),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__750 (
            .O(N__4890),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    CascadeMux I__749 (
            .O(N__4885),
            .I(N__4881));
    InMux I__748 (
            .O(N__4884),
            .I(N__4878));
    InMux I__747 (
            .O(N__4881),
            .I(N__4875));
    LocalMux I__746 (
            .O(N__4878),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__745 (
            .O(N__4875),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__744 (
            .O(N__4870),
            .I(N__4866));
    InMux I__743 (
            .O(N__4869),
            .I(N__4863));
    LocalMux I__742 (
            .O(N__4866),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ));
    LocalMux I__741 (
            .O(N__4863),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ));
    InMux I__740 (
            .O(N__4858),
            .I(N__4854));
    InMux I__739 (
            .O(N__4857),
            .I(N__4851));
    LocalMux I__738 (
            .O(N__4854),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__737 (
            .O(N__4851),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__736 (
            .O(N__4846),
            .I(N__4842));
    InMux I__735 (
            .O(N__4845),
            .I(N__4839));
    LocalMux I__734 (
            .O(N__4842),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__733 (
            .O(N__4839),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    CascadeMux I__732 (
            .O(N__4834),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0_cascade_ ));
    InMux I__731 (
            .O(N__4831),
            .I(N__4828));
    LocalMux I__730 (
            .O(N__4828),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ));
    CascadeMux I__729 (
            .O(N__4825),
            .I(N__4821));
    CascadeMux I__728 (
            .O(N__4824),
            .I(N__4818));
    InMux I__727 (
            .O(N__4821),
            .I(N__4815));
    InMux I__726 (
            .O(N__4818),
            .I(N__4812));
    LocalMux I__725 (
            .O(N__4815),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    LocalMux I__724 (
            .O(N__4812),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    CascadeMux I__723 (
            .O(N__4807),
            .I(\U712_CYCLE_TERM.N_305_i_0_en_cascade_ ));
    InMux I__722 (
            .O(N__4804),
            .I(N__4800));
    InMux I__721 (
            .O(N__4803),
            .I(N__4797));
    LocalMux I__720 (
            .O(N__4800),
            .I(N__4792));
    LocalMux I__719 (
            .O(N__4797),
            .I(N__4792));
    Span12Mux_v I__718 (
            .O(N__4792),
            .I(N__4789));
    Span12Mux_v I__717 (
            .O(N__4789),
            .I(N__4786));
    Span12Mux_h I__716 (
            .O(N__4786),
            .I(N__4783));
    Odrv12 I__715 (
            .O(N__4783),
            .I(DRA_c_0));
    InMux I__714 (
            .O(N__4780),
            .I(N__4777));
    LocalMux I__713 (
            .O(N__4777),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__712 (
            .O(N__4774),
            .I(N__4771));
    LocalMux I__711 (
            .O(N__4771),
            .I(N__4767));
    InMux I__710 (
            .O(N__4770),
            .I(N__4764));
    Span4Mux_v I__709 (
            .O(N__4767),
            .I(N__4761));
    LocalMux I__708 (
            .O(N__4764),
            .I(N__4758));
    Span4Mux_h I__707 (
            .O(N__4761),
            .I(N__4753));
    Span4Mux_v I__706 (
            .O(N__4758),
            .I(N__4753));
    Sp12to4 I__705 (
            .O(N__4753),
            .I(N__4750));
    Span12Mux_h I__704 (
            .O(N__4750),
            .I(N__4747));
    Span12Mux_v I__703 (
            .O(N__4747),
            .I(N__4744));
    Odrv12 I__702 (
            .O(N__4744),
            .I(DRA_c_1));
    InMux I__701 (
            .O(N__4741),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__700 (
            .O(N__4738),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__699 (
            .O(N__4735),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__698 (
            .O(N__4732),
            .I(N__4728));
    InMux I__697 (
            .O(N__4731),
            .I(N__4725));
    LocalMux I__696 (
            .O(N__4728),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__695 (
            .O(N__4725),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__694 (
            .O(N__4720),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__693 (
            .O(N__4717),
            .I(N__4713));
    InMux I__692 (
            .O(N__4716),
            .I(N__4710));
    LocalMux I__691 (
            .O(N__4713),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__690 (
            .O(N__4710),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__689 (
            .O(N__4705),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__688 (
            .O(N__4702),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    ClkMux I__687 (
            .O(N__4699),
            .I(N__4696));
    GlobalMux I__686 (
            .O(N__4696),
            .I(N__4693));
    gio2CtrlBuf I__685 (
            .O(N__4693),
            .I(C1_c_g));
    InMux I__684 (
            .O(N__4690),
            .I(N__4686));
    InMux I__683 (
            .O(N__4689),
            .I(N__4683));
    LocalMux I__682 (
            .O(N__4686),
            .I(\U712_REG_SM.N_306 ));
    LocalMux I__681 (
            .O(N__4683),
            .I(\U712_REG_SM.N_306 ));
    CascadeMux I__680 (
            .O(N__4678),
            .I(N__4675));
    InMux I__679 (
            .O(N__4675),
            .I(N__4669));
    InMux I__678 (
            .O(N__4674),
            .I(N__4666));
    InMux I__677 (
            .O(N__4673),
            .I(N__4661));
    InMux I__676 (
            .O(N__4672),
            .I(N__4661));
    LocalMux I__675 (
            .O(N__4669),
            .I(N__4658));
    LocalMux I__674 (
            .O(N__4666),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    LocalMux I__673 (
            .O(N__4661),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    Odrv4 I__672 (
            .O(N__4658),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    InMux I__671 (
            .O(N__4651),
            .I(N__4646));
    InMux I__670 (
            .O(N__4650),
            .I(N__4641));
    InMux I__669 (
            .O(N__4649),
            .I(N__4641));
    LocalMux I__668 (
            .O(N__4646),
            .I(\U712_REG_SM.N_298 ));
    LocalMux I__667 (
            .O(N__4641),
            .I(\U712_REG_SM.N_298 ));
    CascadeMux I__666 (
            .O(N__4636),
            .I(N__4633));
    InMux I__665 (
            .O(N__4633),
            .I(N__4629));
    InMux I__664 (
            .O(N__4632),
            .I(N__4625));
    LocalMux I__663 (
            .O(N__4629),
            .I(N__4622));
    InMux I__662 (
            .O(N__4628),
            .I(N__4619));
    LocalMux I__661 (
            .O(N__4625),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    Odrv4 I__660 (
            .O(N__4622),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__659 (
            .O(N__4619),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    InMux I__658 (
            .O(N__4612),
            .I(N__4608));
    CascadeMux I__657 (
            .O(N__4611),
            .I(N__4605));
    LocalMux I__656 (
            .O(N__4608),
            .I(N__4602));
    InMux I__655 (
            .O(N__4605),
            .I(N__4599));
    Odrv4 I__654 (
            .O(N__4602),
            .I(\U712_REG_SM.UDS_OUTZ0 ));
    LocalMux I__653 (
            .O(N__4599),
            .I(\U712_REG_SM.UDS_OUTZ0 ));
    IoInMux I__652 (
            .O(N__4594),
            .I(N__4591));
    LocalMux I__651 (
            .O(N__4591),
            .I(N__4588));
    Span12Mux_s4_v I__650 (
            .O(N__4588),
            .I(N__4585));
    Span12Mux_h I__649 (
            .O(N__4585),
            .I(N__4582));
    Odrv12 I__648 (
            .O(N__4582),
            .I(U712_REG_SM_un1_UDSn_i));
    InMux I__647 (
            .O(N__4579),
            .I(N__4567));
    InMux I__646 (
            .O(N__4578),
            .I(N__4567));
    InMux I__645 (
            .O(N__4577),
            .I(N__4567));
    InMux I__644 (
            .O(N__4576),
            .I(N__4567));
    LocalMux I__643 (
            .O(N__4567),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    CascadeMux I__642 (
            .O(N__4564),
            .I(N__4560));
    InMux I__641 (
            .O(N__4563),
            .I(N__4554));
    InMux I__640 (
            .O(N__4560),
            .I(N__4554));
    InMux I__639 (
            .O(N__4559),
            .I(N__4551));
    LocalMux I__638 (
            .O(N__4554),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__637 (
            .O(N__4551),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    InMux I__636 (
            .O(N__4546),
            .I(N__4542));
    InMux I__635 (
            .O(N__4545),
            .I(N__4539));
    LocalMux I__634 (
            .O(N__4542),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    LocalMux I__633 (
            .O(N__4539),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    InMux I__632 (
            .O(N__4534),
            .I(N__4531));
    LocalMux I__631 (
            .O(N__4531),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ));
    IoInMux I__630 (
            .O(N__4528),
            .I(N__4525));
    LocalMux I__629 (
            .O(N__4525),
            .I(N__4522));
    IoSpan4Mux I__628 (
            .O(N__4522),
            .I(N__4519));
    Span4Mux_s3_h I__627 (
            .O(N__4519),
            .I(N__4516));
    Span4Mux_h I__626 (
            .O(N__4516),
            .I(N__4513));
    Span4Mux_h I__625 (
            .O(N__4513),
            .I(N__4510));
    Odrv4 I__624 (
            .O(N__4510),
            .I(N_886_i));
    InMux I__623 (
            .O(N__4507),
            .I(N__4504));
    LocalMux I__622 (
            .O(N__4504),
            .I(N__4501));
    Span4Mux_v I__621 (
            .O(N__4501),
            .I(N__4498));
    Sp12to4 I__620 (
            .O(N__4498),
            .I(N__4495));
    Span12Mux_h I__619 (
            .O(N__4495),
            .I(N__4492));
    Span12Mux_v I__618 (
            .O(N__4492),
            .I(N__4489));
    Odrv12 I__617 (
            .O(N__4489),
            .I(A_c_4));
    CascadeMux I__616 (
            .O(N__4486),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_2_cascade_ ));
    InMux I__615 (
            .O(N__4483),
            .I(N__4480));
    LocalMux I__614 (
            .O(N__4480),
            .I(N__4477));
    Span12Mux_h I__613 (
            .O(N__4477),
            .I(N__4474));
    Odrv12 I__612 (
            .O(N__4474),
            .I(A_c_11));
    InMux I__611 (
            .O(N__4471),
            .I(bfn_11_9_0_));
    InMux I__610 (
            .O(N__4468),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__609 (
            .O(N__4465),
            .I(N__4462));
    LocalMux I__608 (
            .O(N__4462),
            .I(N__4456));
    InMux I__607 (
            .O(N__4461),
            .I(N__4453));
    InMux I__606 (
            .O(N__4460),
            .I(N__4448));
    InMux I__605 (
            .O(N__4459),
            .I(N__4448));
    Odrv4 I__604 (
            .O(N__4456),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    LocalMux I__603 (
            .O(N__4453),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    LocalMux I__602 (
            .O(N__4448),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    InMux I__601 (
            .O(N__4441),
            .I(N__4437));
    InMux I__600 (
            .O(N__4440),
            .I(N__4431));
    LocalMux I__599 (
            .O(N__4437),
            .I(N__4428));
    InMux I__598 (
            .O(N__4436),
            .I(N__4425));
    InMux I__597 (
            .O(N__4435),
            .I(N__4420));
    InMux I__596 (
            .O(N__4434),
            .I(N__4420));
    LocalMux I__595 (
            .O(N__4431),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__594 (
            .O(N__4428),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__593 (
            .O(N__4425),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__592 (
            .O(N__4420),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    CascadeMux I__591 (
            .O(N__4411),
            .I(N__4407));
    CascadeMux I__590 (
            .O(N__4410),
            .I(N__4404));
    InMux I__589 (
            .O(N__4407),
            .I(N__4399));
    InMux I__588 (
            .O(N__4404),
            .I(N__4399));
    LocalMux I__587 (
            .O(N__4399),
            .I(\U712_REG_SM.N_289 ));
    InMux I__586 (
            .O(N__4396),
            .I(N__4392));
    InMux I__585 (
            .O(N__4395),
            .I(N__4389));
    LocalMux I__584 (
            .O(N__4392),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    LocalMux I__583 (
            .O(N__4389),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    InMux I__582 (
            .O(N__4384),
            .I(N__4375));
    InMux I__581 (
            .O(N__4383),
            .I(N__4368));
    InMux I__580 (
            .O(N__4382),
            .I(N__4368));
    InMux I__579 (
            .O(N__4381),
            .I(N__4368));
    InMux I__578 (
            .O(N__4380),
            .I(N__4361));
    InMux I__577 (
            .O(N__4379),
            .I(N__4361));
    InMux I__576 (
            .O(N__4378),
            .I(N__4361));
    LocalMux I__575 (
            .O(N__4375),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__574 (
            .O(N__4368),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__573 (
            .O(N__4361),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    CascadeMux I__572 (
            .O(N__4354),
            .I(\U712_REG_SM.N_289_cascade_ ));
    InMux I__571 (
            .O(N__4351),
            .I(N__4341));
    InMux I__570 (
            .O(N__4350),
            .I(N__4341));
    InMux I__569 (
            .O(N__4349),
            .I(N__4336));
    InMux I__568 (
            .O(N__4348),
            .I(N__4331));
    InMux I__567 (
            .O(N__4347),
            .I(N__4331));
    InMux I__566 (
            .O(N__4346),
            .I(N__4328));
    LocalMux I__565 (
            .O(N__4341),
            .I(N__4325));
    InMux I__564 (
            .O(N__4340),
            .I(N__4320));
    InMux I__563 (
            .O(N__4339),
            .I(N__4320));
    LocalMux I__562 (
            .O(N__4336),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__561 (
            .O(N__4331),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__560 (
            .O(N__4328),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    Odrv4 I__559 (
            .O(N__4325),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__558 (
            .O(N__4320),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    InMux I__557 (
            .O(N__4309),
            .I(N__4303));
    InMux I__556 (
            .O(N__4308),
            .I(N__4303));
    LocalMux I__555 (
            .O(N__4303),
            .I(\U712_REG_SM.N_494 ));
    CascadeMux I__554 (
            .O(N__4300),
            .I(N__4296));
    InMux I__553 (
            .O(N__4299),
            .I(N__4288));
    InMux I__552 (
            .O(N__4296),
            .I(N__4288));
    InMux I__551 (
            .O(N__4295),
            .I(N__4281));
    InMux I__550 (
            .O(N__4294),
            .I(N__4281));
    InMux I__549 (
            .O(N__4293),
            .I(N__4281));
    LocalMux I__548 (
            .O(N__4288),
            .I(\U712_REG_SM.N_288 ));
    LocalMux I__547 (
            .O(N__4281),
            .I(\U712_REG_SM.N_288 ));
    CascadeMux I__546 (
            .O(N__4276),
            .I(\U712_REG_SM.N_494_cascade_ ));
    InMux I__545 (
            .O(N__4273),
            .I(N__4269));
    InMux I__544 (
            .O(N__4272),
            .I(N__4266));
    LocalMux I__543 (
            .O(N__4269),
            .I(\U712_REG_SM.N_424 ));
    LocalMux I__542 (
            .O(N__4266),
            .I(\U712_REG_SM.N_424 ));
    InMux I__541 (
            .O(N__4261),
            .I(N__4258));
    LocalMux I__540 (
            .O(N__4258),
            .I(\U712_REG_SM.N_369 ));
    CascadeMux I__539 (
            .O(N__4255),
            .I(\U712_REG_SM.DS_EN_RNOZ0Z_2_cascade_ ));
    InMux I__538 (
            .O(N__4252),
            .I(N__4249));
    LocalMux I__537 (
            .O(N__4249),
            .I(\U712_REG_SM.N_123 ));
    IoInMux I__536 (
            .O(N__4246),
            .I(N__4243));
    LocalMux I__535 (
            .O(N__4243),
            .I(N__4240));
    Span12Mux_s1_h I__534 (
            .O(N__4240),
            .I(N__4237));
    Span12Mux_h I__533 (
            .O(N__4237),
            .I(N__4233));
    InMux I__532 (
            .O(N__4236),
            .I(N__4230));
    Odrv12 I__531 (
            .O(N__4233),
            .I(TACK_OUTn));
    LocalMux I__530 (
            .O(N__4230),
            .I(TACK_OUTn));
    InMux I__529 (
            .O(N__4225),
            .I(N__4222));
    LocalMux I__528 (
            .O(N__4222),
            .I(N__4216));
    InMux I__527 (
            .O(N__4221),
            .I(N__4209));
    InMux I__526 (
            .O(N__4220),
            .I(N__4209));
    InMux I__525 (
            .O(N__4219),
            .I(N__4209));
    Span4Mux_v I__524 (
            .O(N__4216),
            .I(N__4204));
    LocalMux I__523 (
            .O(N__4209),
            .I(N__4204));
    Span4Mux_h I__522 (
            .O(N__4204),
            .I(N__4201));
    Sp12to4 I__521 (
            .O(N__4201),
            .I(N__4198));
    Span12Mux_v I__520 (
            .O(N__4198),
            .I(N__4195));
    Odrv12 I__519 (
            .O(N__4195),
            .I(CLK40_OUT_i));
    InMux I__518 (
            .O(N__4192),
            .I(N__4189));
    LocalMux I__517 (
            .O(N__4189),
            .I(\U712_BYTE_ENABLE.N_395 ));
    IoInMux I__516 (
            .O(N__4186),
            .I(N__4183));
    LocalMux I__515 (
            .O(N__4183),
            .I(N__4180));
    IoSpan4Mux I__514 (
            .O(N__4180),
            .I(N__4177));
    Span4Mux_s3_h I__513 (
            .O(N__4177),
            .I(N__4174));
    Sp12to4 I__512 (
            .O(N__4174),
            .I(N__4171));
    Span12Mux_s8_h I__511 (
            .O(N__4171),
            .I(N__4168));
    Span12Mux_v I__510 (
            .O(N__4168),
            .I(N__4165));
    Odrv12 I__509 (
            .O(N__4165),
            .I(N_74_i));
    InMux I__508 (
            .O(N__4162),
            .I(N__4153));
    InMux I__507 (
            .O(N__4161),
            .I(N__4153));
    InMux I__506 (
            .O(N__4160),
            .I(N__4153));
    LocalMux I__505 (
            .O(N__4153),
            .I(\U712_BYTE_ENABLE.N_387 ));
    InMux I__504 (
            .O(N__4150),
            .I(N__4140));
    InMux I__503 (
            .O(N__4149),
            .I(N__4140));
    InMux I__502 (
            .O(N__4148),
            .I(N__4140));
    InMux I__501 (
            .O(N__4147),
            .I(N__4137));
    LocalMux I__500 (
            .O(N__4140),
            .I(N__4132));
    LocalMux I__499 (
            .O(N__4137),
            .I(N__4132));
    Span4Mux_h I__498 (
            .O(N__4132),
            .I(N__4129));
    Sp12to4 I__497 (
            .O(N__4129),
            .I(N__4126));
    Span12Mux_v I__496 (
            .O(N__4126),
            .I(N__4123));
    Odrv12 I__495 (
            .O(N__4123),
            .I(A_c_1));
    CascadeMux I__494 (
            .O(N__4120),
            .I(N__4117));
    InMux I__493 (
            .O(N__4117),
            .I(N__4111));
    InMux I__492 (
            .O(N__4116),
            .I(N__4111));
    LocalMux I__491 (
            .O(N__4111),
            .I(\U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_0_0 ));
    IoInMux I__490 (
            .O(N__4108),
            .I(N__4105));
    LocalMux I__489 (
            .O(N__4105),
            .I(N__4102));
    Span12Mux_s6_h I__488 (
            .O(N__4102),
            .I(N__4099));
    Span12Mux_h I__487 (
            .O(N__4099),
            .I(N__4096));
    Odrv12 I__486 (
            .O(N__4096),
            .I(N_76_i));
    CascadeMux I__485 (
            .O(N__4093),
            .I(N__4090));
    InMux I__484 (
            .O(N__4090),
            .I(N__4087));
    LocalMux I__483 (
            .O(N__4087),
            .I(\U712_BYTE_ENABLE.N_391 ));
    InMux I__482 (
            .O(N__4084),
            .I(N__4080));
    InMux I__481 (
            .O(N__4083),
            .I(N__4077));
    LocalMux I__480 (
            .O(N__4080),
            .I(\U712_REG_SM.N_304 ));
    LocalMux I__479 (
            .O(N__4077),
            .I(\U712_REG_SM.N_304 ));
    CascadeMux I__478 (
            .O(N__4072),
            .I(N__4068));
    InMux I__477 (
            .O(N__4071),
            .I(N__4060));
    InMux I__476 (
            .O(N__4068),
            .I(N__4060));
    InMux I__475 (
            .O(N__4067),
            .I(N__4060));
    LocalMux I__474 (
            .O(N__4060),
            .I(\U712_REG_SM.N_299 ));
    InMux I__473 (
            .O(N__4057),
            .I(N__4048));
    InMux I__472 (
            .O(N__4056),
            .I(N__4048));
    InMux I__471 (
            .O(N__4055),
            .I(N__4048));
    LocalMux I__470 (
            .O(N__4048),
            .I(\U712_REG_SM.N_281 ));
    InMux I__469 (
            .O(N__4045),
            .I(N__4040));
    InMux I__468 (
            .O(N__4044),
            .I(N__4037));
    InMux I__467 (
            .O(N__4043),
            .I(N__4034));
    LocalMux I__466 (
            .O(N__4040),
            .I(\U712_REG_SM.N_280 ));
    LocalMux I__465 (
            .O(N__4037),
            .I(\U712_REG_SM.N_280 ));
    LocalMux I__464 (
            .O(N__4034),
            .I(\U712_REG_SM.N_280 ));
    CascadeMux I__463 (
            .O(N__4027),
            .I(\U712_REG_SM.N_373_cascade_ ));
    CascadeMux I__462 (
            .O(N__4024),
            .I(\U712_REG_SM.N_288_cascade_ ));
    InMux I__461 (
            .O(N__4021),
            .I(N__4014));
    InMux I__460 (
            .O(N__4020),
            .I(N__4014));
    InMux I__459 (
            .O(N__4019),
            .I(N__4011));
    LocalMux I__458 (
            .O(N__4014),
            .I(\U712_REG_SM.N_307 ));
    LocalMux I__457 (
            .O(N__4011),
            .I(\U712_REG_SM.N_307 ));
    CascadeMux I__456 (
            .O(N__4006),
            .I(N__4003));
    InMux I__455 (
            .O(N__4003),
            .I(N__3999));
    InMux I__454 (
            .O(N__4002),
            .I(N__3996));
    LocalMux I__453 (
            .O(N__3999),
            .I(\U712_REG_SM.C1_SYNCZ0Z_2 ));
    LocalMux I__452 (
            .O(N__3996),
            .I(\U712_REG_SM.C1_SYNCZ0Z_2 ));
    InMux I__451 (
            .O(N__3991),
            .I(N__3988));
    LocalMux I__450 (
            .O(N__3988),
            .I(N__3985));
    Span4Mux_v I__449 (
            .O(N__3985),
            .I(N__3982));
    Sp12to4 I__448 (
            .O(N__3982),
            .I(N__3979));
    Span12Mux_h I__447 (
            .O(N__3979),
            .I(N__3976));
    Odrv12 I__446 (
            .O(N__3976),
            .I(C3_c));
    IoInMux I__445 (
            .O(N__3973),
            .I(N__3969));
    InMux I__444 (
            .O(N__3972),
            .I(N__3966));
    LocalMux I__443 (
            .O(N__3969),
            .I(N__3963));
    LocalMux I__442 (
            .O(N__3966),
            .I(N__3960));
    Span4Mux_s3_h I__441 (
            .O(N__3963),
            .I(N__3957));
    Span12Mux_h I__440 (
            .O(N__3960),
            .I(N__3952));
    Sp12to4 I__439 (
            .O(N__3957),
            .I(N__3952));
    Span12Mux_v I__438 (
            .O(N__3952),
            .I(N__3949));
    Odrv12 I__437 (
            .O(N__3949),
            .I(C1_c));
    InMux I__436 (
            .O(N__3946),
            .I(N__3940));
    InMux I__435 (
            .O(N__3945),
            .I(N__3933));
    InMux I__434 (
            .O(N__3944),
            .I(N__3933));
    InMux I__433 (
            .O(N__3943),
            .I(N__3933));
    LocalMux I__432 (
            .O(N__3940),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__431 (
            .O(N__3933),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    InMux I__430 (
            .O(N__3928),
            .I(N__3924));
    InMux I__429 (
            .O(N__3927),
            .I(N__3921));
    LocalMux I__428 (
            .O(N__3924),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2Z0Z_0 ));
    LocalMux I__427 (
            .O(N__3921),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2Z0Z_0 ));
    IoInMux I__426 (
            .O(N__3916),
            .I(N__3913));
    LocalMux I__425 (
            .O(N__3913),
            .I(N__3910));
    Span4Mux_s2_h I__424 (
            .O(N__3910),
            .I(N__3907));
    Span4Mux_h I__423 (
            .O(N__3907),
            .I(N__3904));
    Sp12to4 I__422 (
            .O(N__3904),
            .I(N__3901));
    Span12Mux_s11_v I__421 (
            .O(N__3901),
            .I(N__3898));
    Span12Mux_h I__420 (
            .O(N__3898),
            .I(N__3895));
    Odrv12 I__419 (
            .O(N__3895),
            .I(N_75_i));
    InMux I__418 (
            .O(N__3892),
            .I(N__3886));
    InMux I__417 (
            .O(N__3891),
            .I(N__3886));
    LocalMux I__416 (
            .O(N__3886),
            .I(\U712_REG_SM.N_301 ));
    InMux I__415 (
            .O(N__3883),
            .I(N__3877));
    InMux I__414 (
            .O(N__3882),
            .I(N__3877));
    LocalMux I__413 (
            .O(N__3877),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    IoInMux I__412 (
            .O(N__3874),
            .I(N__3870));
    IoInMux I__411 (
            .O(N__3873),
            .I(N__3867));
    LocalMux I__410 (
            .O(N__3870),
            .I(N__3864));
    LocalMux I__409 (
            .O(N__3867),
            .I(N__3861));
    IoSpan4Mux I__408 (
            .O(N__3864),
            .I(N__3858));
    IoSpan4Mux I__407 (
            .O(N__3861),
            .I(N__3855));
    Span4Mux_s3_v I__406 (
            .O(N__3858),
            .I(N__3852));
    Span4Mux_s3_v I__405 (
            .O(N__3855),
            .I(N__3849));
    Sp12to4 I__404 (
            .O(N__3852),
            .I(N__3846));
    Sp12to4 I__403 (
            .O(N__3849),
            .I(N__3843));
    Span12Mux_s9_h I__402 (
            .O(N__3846),
            .I(N__3839));
    Span12Mux_s10_h I__401 (
            .O(N__3843),
            .I(N__3836));
    CascadeMux I__400 (
            .O(N__3842),
            .I(N__3833));
    Span12Mux_v I__399 (
            .O(N__3839),
            .I(N__3828));
    Span12Mux_v I__398 (
            .O(N__3836),
            .I(N__3828));
    InMux I__397 (
            .O(N__3833),
            .I(N__3825));
    Odrv12 I__396 (
            .O(N__3828),
            .I(ASn_c));
    LocalMux I__395 (
            .O(N__3825),
            .I(ASn_c));
    InMux I__394 (
            .O(N__3820),
            .I(N__3815));
    InMux I__393 (
            .O(N__3819),
            .I(N__3810));
    InMux I__392 (
            .O(N__3818),
            .I(N__3810));
    LocalMux I__391 (
            .O(N__3815),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__390 (
            .O(N__3810),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    CascadeMux I__389 (
            .O(N__3805),
            .I(N__3802));
    InMux I__388 (
            .O(N__3802),
            .I(N__3795));
    InMux I__387 (
            .O(N__3801),
            .I(N__3795));
    InMux I__386 (
            .O(N__3800),
            .I(N__3792));
    LocalMux I__385 (
            .O(N__3795),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__384 (
            .O(N__3792),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    CascadeMux I__383 (
            .O(N__3787),
            .I(\U712_REG_SM.N_281_cascade_ ));
    CascadeMux I__382 (
            .O(N__3784),
            .I(\U712_REG_SM.N_280_cascade_ ));
    CascadeMux I__381 (
            .O(N__3781),
            .I(N__3777));
    CascadeMux I__380 (
            .O(N__3780),
            .I(N__3774));
    InMux I__379 (
            .O(N__3777),
            .I(N__3769));
    InMux I__378 (
            .O(N__3774),
            .I(N__3766));
    InMux I__377 (
            .O(N__3773),
            .I(N__3761));
    InMux I__376 (
            .O(N__3772),
            .I(N__3761));
    LocalMux I__375 (
            .O(N__3769),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__374 (
            .O(N__3766),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__373 (
            .O(N__3761),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    InMux I__372 (
            .O(N__3754),
            .I(N__3748));
    InMux I__371 (
            .O(N__3753),
            .I(N__3748));
    LocalMux I__370 (
            .O(N__3748),
            .I(\U712_REG_SM.N_308 ));
    InMux I__369 (
            .O(N__3745),
            .I(N__3742));
    LocalMux I__368 (
            .O(N__3742),
            .I(N__3739));
    Span4Mux_v I__367 (
            .O(N__3739),
            .I(N__3735));
    InMux I__366 (
            .O(N__3738),
            .I(N__3732));
    Sp12to4 I__365 (
            .O(N__3735),
            .I(N__3727));
    LocalMux I__364 (
            .O(N__3732),
            .I(N__3727));
    Span12Mux_h I__363 (
            .O(N__3727),
            .I(N__3724));
    Span12Mux_v I__362 (
            .O(N__3724),
            .I(N__3721));
    Odrv12 I__361 (
            .O(N__3721),
            .I(SIZ_c_0));
    CascadeMux I__360 (
            .O(N__3718),
            .I(\U712_BYTE_ENABLE.N_387_cascade_ ));
    IoInMux I__359 (
            .O(N__3715),
            .I(N__3712));
    LocalMux I__358 (
            .O(N__3712),
            .I(N__3709));
    Span4Mux_s2_v I__357 (
            .O(N__3709),
            .I(N__3706));
    Span4Mux_v I__356 (
            .O(N__3706),
            .I(N__3703));
    Span4Mux_v I__355 (
            .O(N__3703),
            .I(N__3700));
    Span4Mux_v I__354 (
            .O(N__3700),
            .I(N__3697));
    Odrv4 I__353 (
            .O(N__3697),
            .I(N_73_i));
    InMux I__352 (
            .O(N__3694),
            .I(N__3690));
    InMux I__351 (
            .O(N__3693),
            .I(N__3687));
    LocalMux I__350 (
            .O(N__3690),
            .I(N__3682));
    LocalMux I__349 (
            .O(N__3687),
            .I(N__3682));
    Span4Mux_v I__348 (
            .O(N__3682),
            .I(N__3677));
    InMux I__347 (
            .O(N__3681),
            .I(N__3672));
    InMux I__346 (
            .O(N__3680),
            .I(N__3672));
    Span4Mux_v I__345 (
            .O(N__3677),
            .I(N__3669));
    LocalMux I__344 (
            .O(N__3672),
            .I(N__3666));
    Sp12to4 I__343 (
            .O(N__3669),
            .I(N__3661));
    Span12Mux_v I__342 (
            .O(N__3666),
            .I(N__3661));
    Odrv12 I__341 (
            .O(N__3661),
            .I(A_c_0));
    InMux I__340 (
            .O(N__3658),
            .I(N__3655));
    LocalMux I__339 (
            .O(N__3655),
            .I(N__3651));
    InMux I__338 (
            .O(N__3654),
            .I(N__3648));
    Span4Mux_v I__337 (
            .O(N__3651),
            .I(N__3643));
    LocalMux I__336 (
            .O(N__3648),
            .I(N__3643));
    Span4Mux_h I__335 (
            .O(N__3643),
            .I(N__3640));
    Sp12to4 I__334 (
            .O(N__3640),
            .I(N__3637));
    Span12Mux_v I__333 (
            .O(N__3637),
            .I(N__3634));
    Odrv12 I__332 (
            .O(N__3634),
            .I(SIZ_c_1));
    InMux I__331 (
            .O(N__3631),
            .I(N__3628));
    LocalMux I__330 (
            .O(N__3628),
            .I(N__3625));
    Span4Mux_v I__329 (
            .O(N__3625),
            .I(N__3622));
    Sp12to4 I__328 (
            .O(N__3622),
            .I(N__3619));
    Span12Mux_h I__327 (
            .O(N__3619),
            .I(N__3616));
    Span12Mux_v I__326 (
            .O(N__3616),
            .I(N__3613));
    Odrv12 I__325 (
            .O(N__3613),
            .I(REGSPACEn_c));
    IoInMux I__324 (
            .O(N__3610),
            .I(N__3607));
    LocalMux I__323 (
            .O(N__3607),
            .I(N__3604));
    Span4Mux_s3_v I__322 (
            .O(N__3604),
            .I(N__3601));
    Span4Mux_h I__321 (
            .O(N__3601),
            .I(N__3598));
    Odrv4 I__320 (
            .O(N__3598),
            .I(CLK80_OUT_i_i));
    IoInMux I__319 (
            .O(N__3595),
            .I(N__3592));
    LocalMux I__318 (
            .O(N__3592),
            .I(N__3589));
    Span12Mux_s6_h I__317 (
            .O(N__3589),
            .I(N__3586));
    Odrv12 I__316 (
            .O(N__3586),
            .I(CLK40_OUT_i_i));
    CascadeMux I__315 (
            .O(N__3583),
            .I(N__3579));
    InMux I__314 (
            .O(N__3582),
            .I(N__3574));
    InMux I__313 (
            .O(N__3579),
            .I(N__3574));
    LocalMux I__312 (
            .O(N__3574),
            .I(\U712_REG_SM.LDS_OUT_2_0_a2Z0Z_0 ));
    IoInMux I__311 (
            .O(N__3571),
            .I(N__3568));
    LocalMux I__310 (
            .O(N__3568),
            .I(N__3565));
    Span4Mux_s1_v I__309 (
            .O(N__3565),
            .I(N__3562));
    Span4Mux_v I__308 (
            .O(N__3562),
            .I(N__3559));
    Span4Mux_v I__307 (
            .O(N__3559),
            .I(N__3556));
    Odrv4 I__306 (
            .O(N__3556),
            .I(VBENn_c));
    IoInMux I__305 (
            .O(N__3553),
            .I(N__3550));
    LocalMux I__304 (
            .O(N__3550),
            .I(N__3547));
    IoSpan4Mux I__303 (
            .O(N__3547),
            .I(N__3544));
    Span4Mux_s2_v I__302 (
            .O(N__3544),
            .I(N__3541));
    Sp12to4 I__301 (
            .O(N__3541),
            .I(N__3538));
    Span12Mux_v I__300 (
            .O(N__3538),
            .I(N__3535));
    Odrv12 I__299 (
            .O(N__3535),
            .I(CLK40_IN_c));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_9_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__5023),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__3973),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_3_1_0.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_3_1_0.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_3_1_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLKRAM_obuf_RNO_LC_3_1_0 (
            .in0(N__9163),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK80_OUT_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDS_OUT_2_0_a2_0_LC_7_12_3 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_2_0_a2_0_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDS_OUT_2_0_a2_0_LC_7_12_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_REG_SM.LDS_OUT_2_0_a2_0_LC_7_12_3  (
            .in0(_gnd_net_),
            .in1(N__6878),
            .in2(_gnd_net_),
            .in3(N__3738),
            .lcout(\U712_REG_SM.LDS_OUT_2_0_a2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLK40C_obuf_RNO_LC_8_10_1.C_ON=1'b0;
    defparam CLK40C_obuf_RNO_LC_8_10_1.SEQ_MODE=4'b0000;
    defparam CLK40C_obuf_RNO_LC_8_10_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLK40C_obuf_RNO_LC_8_10_1 (
            .in0(N__4225),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_OUT_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.UDS_OUT_LC_8_12_4 .C_ON=1'b0;
    defparam \U712_REG_SM.UDS_OUT_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.UDS_OUT_LC_8_12_4 .LUT_INIT=16'b1011000111110101;
    LogicCell40 \U712_REG_SM.UDS_OUT_LC_8_12_4  (
            .in0(N__3754),
            .in1(N__3681),
            .in2(N__4611),
            .in3(N__3582),
            .lcout(\U712_REG_SM.UDS_OUTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9158),
            .ce(),
            .sr(N__8944));
    defparam \U712_REG_SM.LDS_OUT_LC_8_12_7 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_LC_8_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.LDS_OUT_LC_8_12_7 .LUT_INIT=16'b1100110010101111;
    LogicCell40 \U712_REG_SM.LDS_OUT_LC_8_12_7  (
            .in0(N__3680),
            .in1(N__5919),
            .in2(N__3583),
            .in3(N__3753),
            .lcout(\U712_REG_SM.LDS_OUTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9158),
            .ce(),
            .sr(N__8944));
    defparam \U712_BUFFERS.un1_VBENn_0_a2_0_a2_LC_9_4_1 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_0_a2_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_0_a2_LC_9_4_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a2_0_a2_LC_9_4_1  (
            .in0(_gnd_net_),
            .in1(N__6826),
            .in2(_gnd_net_),
            .in3(N__7496),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_1_0_LC_9_9_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_1_0_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_1_0_LC_9_9_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_1_0_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__6820),
            .in2(_gnd_net_),
            .in3(N__3694),
            .lcout(\U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_9_9_2 .LUT_INIT=16'b1000100001000100;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_9_9_2  (
            .in0(N__3658),
            .in1(N__6821),
            .in2(_gnd_net_),
            .in3(N__3745),
            .lcout(\U712_BYTE_ENABLE.N_387 ),
            .ltout(\U712_BYTE_ENABLE.N_387_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_73_i_LC_9_9_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_73_i_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_73_i_LC_9_9_3 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \U712_BYTE_ENABLE.N_73_i_LC_9_9_3  (
            .in0(N__4192),
            .in1(N__4147),
            .in2(N__3718),
            .in3(N__3927),
            .lcout(N_73_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_0_LC_9_10_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_0_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_0_LC_9_10_2 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_0_LC_9_10_2  (
            .in0(N__6822),
            .in1(N__3693),
            .in2(_gnd_net_),
            .in3(N__3654),
            .lcout(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_srsts_0_i_o3_0_LC_9_10_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_srsts_0_i_o3_0_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_srsts_0_i_o3_0_LC_9_10_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_srsts_0_i_o3_0_LC_9_10_7  (
            .in0(N__5139),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3631),
            .lcout(\U712_REG_SM.N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_9_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_9_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_9_11_1 .LUT_INIT=16'b1111010011000100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_9_11_1  (
            .in0(N__3892),
            .in1(N__3882),
            .in2(N__3780),
            .in3(N__4020),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9155),
            .ce(),
            .sr(N__8945));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_9_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_9_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_9_11_2 .LUT_INIT=16'b1101110000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_9_11_2  (
            .in0(N__4021),
            .in1(N__3801),
            .in2(N__3781),
            .in3(N__4084),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9155),
            .ce(),
            .sr(N__8945));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_9_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_9_11_3 .LUT_INIT=16'b1100111000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_9_11_3  (
            .in0(N__3819),
            .in1(N__4632),
            .in2(N__4072),
            .in3(N__4651),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9155),
            .ce(),
            .sr(N__8945));
    defparam \U712_REG_SM.REG_CYCLE_LC_9_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_9_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_9_11_4 .LUT_INIT=16'b1100101011001110;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_9_11_4  (
            .in0(N__7486),
            .in1(N__3818),
            .in2(N__4678),
            .in3(N__4071),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9155),
            .ce(),
            .sr(N__8945));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_9_11_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_9_11_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_9_11_5 .LUT_INIT=16'b1010111000001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_9_11_5  (
            .in0(N__3891),
            .in1(N__4309),
            .in2(N__4300),
            .in3(N__3883),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9155),
            .ce(),
            .sr(N__8945));
    defparam \U712_REG_SM.REGENn_1_LC_9_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_1_LC_9_11_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_1_LC_9_11_6 .LUT_INIT=16'b1111000010111010;
    LogicCell40 \U712_REG_SM.REGENn_1_LC_9_11_6  (
            .in0(N__4308),
            .in1(N__4273),
            .in2(N__3842),
            .in3(N__4299),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9155),
            .ce(),
            .sr(N__8945));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_9_11_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_9_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_9_11_7 .LUT_INIT=16'b0010101000100000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_9_11_7  (
            .in0(N__4067),
            .in1(N__4083),
            .in2(N__3805),
            .in3(N__3820),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9155),
            .ce(),
            .sr(N__8945));
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_9_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_9_12_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_9_12_0  (
            .in0(N__4339),
            .in1(N__3944),
            .in2(N__4006),
            .in3(N__4379),
            .lcout(\U712_REG_SM.N_281 ),
            .ltout(\U712_REG_SM.N_281_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_9_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_9_12_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_1_LC_9_12_1  (
            .in0(N__3800),
            .in1(N__4460),
            .in2(N__3787),
            .in3(N__4435),
            .lcout(\U712_REG_SM.N_369 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_9_12_2 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_9_12_2 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_0_LC_9_12_2  (
            .in0(N__6879),
            .in1(N__3945),
            .in2(_gnd_net_),
            .in3(N__4351),
            .lcout(\U712_REG_SM.N_123 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_0_2_LC_9_12_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_0_2_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_0_2_LC_9_12_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI90BP_0_2_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__4459),
            .in2(_gnd_net_),
            .in3(N__4434),
            .lcout(\U712_REG_SM.N_280 ),
            .ltout(\U712_REG_SM.N_280_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNINB3L1_1_LC_9_12_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNINB3L1_1_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNINB3L1_1_LC_9_12_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNINB3L1_1_LC_9_12_4  (
            .in0(N__3772),
            .in1(N__4350),
            .in2(N__3784),
            .in3(N__4380),
            .lcout(\U712_REG_SM.N_424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_9_12_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_9_12_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(N__3773),
            .in2(_gnd_net_),
            .in3(N__4019),
            .lcout(\U712_REG_SM.N_308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_9_12_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_9_12_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(N__3943),
            .in2(_gnd_net_),
            .in3(N__4002),
            .lcout(\U712_REG_SM.N_288 ),
            .ltout(\U712_REG_SM.N_288_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_9_12_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_9_12_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_9_12_7  (
            .in0(N__4378),
            .in1(N__4340),
            .in2(N__4024),
            .in3(N__4043),
            .lcout(\U712_REG_SM.N_307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_2_LC_9_13_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_2_LC_9_13_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_2_LC_9_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_2_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4384),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9159),
            .ce(),
            .sr(N__8935));
    defparam \U712_REG_SM.C3_SYNC_0_LC_9_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_9_13_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_9_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3991),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9159),
            .ce(),
            .sr(N__8935));
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_13_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_13_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_9_13_2  (
            .in0(N__3972),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9159),
            .ce(),
            .sr(N__8935));
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_13_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4349),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9159),
            .ce(),
            .sr(N__8935));
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_13_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3946),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9159),
            .ce(),
            .sr(N__8935));
    defparam \U712_REG_SM.C3_SYNC_2_LC_9_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_2_LC_9_13_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_2_LC_9_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_2_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4440),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9159),
            .ce(),
            .sr(N__8935));
    defparam \U712_BYTE_ENABLE.N_75_i_LC_10_9_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_75_i_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_75_i_LC_10_9_1 .LUT_INIT=16'b0000010000000101;
    LogicCell40 \U712_BYTE_ENABLE.N_75_i_LC_10_9_1  (
            .in0(N__4161),
            .in1(N__4149),
            .in2(N__4093),
            .in3(N__3928),
            .lcout(N_75_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_10_9_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_10_9_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_10_9_2  (
            .in0(N__7584),
            .in1(N__5247),
            .in2(_gnd_net_),
            .in3(N__6179),
            .lcout(\U712_BYTE_ENABLE.N_395 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_74_i_LC_10_9_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_74_i_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_74_i_LC_10_9_6 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \U712_BYTE_ENABLE.N_74_i_LC_10_9_6  (
            .in0(N__4148),
            .in1(N__4160),
            .in2(N__5275),
            .in3(N__4116),
            .lcout(N_74_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_76_i_LC_10_9_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_76_i_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_76_i_LC_10_9_7 .LUT_INIT=16'b0000000001000101;
    LogicCell40 \U712_BYTE_ENABLE.N_76_i_LC_10_9_7  (
            .in0(N__4162),
            .in1(N__4150),
            .in2(N__4120),
            .in3(N__5260),
            .lcout(N_76_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_LC_10_10_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_LC_10_10_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_LC_10_10_7  (
            .in0(N__5246),
            .in1(N__7585),
            .in2(_gnd_net_),
            .in3(N__6180),
            .lcout(\U712_BYTE_ENABLE.N_391 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_10_11_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_10_11_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_10_11_0  (
            .in0(N__4056),
            .in1(N__4465),
            .in2(_gnd_net_),
            .in3(N__4441),
            .lcout(\U712_REG_SM.N_304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_10_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_10_11_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_10_11_4  (
            .in0(N__4057),
            .in1(N__4045),
            .in2(N__5782),
            .in3(N__5755),
            .lcout(\U712_REG_SM.N_299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNI0ULC2_4_LC_10_11_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI0ULC2_4_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI0ULC2_4_LC_10_11_5 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI0ULC2_4_LC_10_11_5  (
            .in0(N__4628),
            .in1(N__4055),
            .in2(_gnd_net_),
            .in3(N__4044),
            .lcout(\U712_REG_SM.N_298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_10_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_10_12_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_10_12_0  (
            .in0(N__4348),
            .in1(N__4383),
            .in2(N__4411),
            .in3(N__4295),
            .lcout(),
            .ltout(\U712_REG_SM.N_373_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_6_LC_10_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_10_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_10_12_1 .LUT_INIT=16'b0000101000001110;
    LogicCell40 \U712_REG_SM.STATE_COUNT_6_LC_10_12_1  (
            .in0(N__4396),
            .in1(N__4674),
            .in2(N__4027),
            .in3(N__4689),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9156),
            .ce(),
            .sr(N__8936));
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_0_1_LC_10_12_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_0_1_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_0_1_LC_10_12_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNIIDN62_0_1_LC_10_12_2  (
            .in0(N__4347),
            .in1(N__4382),
            .in2(N__4410),
            .in3(N__4293),
            .lcout(\U712_REG_SM.N_306 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_10_12_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_10_12_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(N__4461),
            .in2(_gnd_net_),
            .in3(N__4436),
            .lcout(\U712_REG_SM.N_289 ),
            .ltout(\U712_REG_SM.N_289_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_10_12_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_10_12_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_10_12_4  (
            .in0(N__4395),
            .in1(N__4381),
            .in2(N__4354),
            .in3(N__4346),
            .lcout(\U712_REG_SM.N_494 ),
            .ltout(\U712_REG_SM.N_494_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_10_12_5 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_10_12_5 .LUT_INIT=16'b0101010101010000;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_2_LC_10_12_5  (
            .in0(N__4294),
            .in1(_gnd_net_),
            .in2(N__4276),
            .in3(N__4272),
            .lcout(),
            .ltout(\U712_REG_SM.DS_EN_RNOZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_LC_10_12_6 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_LC_10_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DS_EN_LC_10_12_6 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \U712_REG_SM.DS_EN_LC_10_12_6  (
            .in0(N__5939),
            .in1(N__4261),
            .in2(N__4255),
            .in3(N__4252),
            .lcout(\U712_REG_SM.DS_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9156),
            .ce(),
            .sr(N__8936));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_10_13_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_10_13_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_10_13_0 .LUT_INIT=16'b1111110011110100;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_10_13_0  (
            .in0(N__4578),
            .in1(N__4236),
            .in2(N__4564),
            .in3(N__4219),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9157),
            .ce(),
            .sr(N__8933));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_10_13_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_10_13_1 .LUT_INIT=16'b1100100011111000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_10_13_1  (
            .in0(N__4220),
            .in1(N__4579),
            .in2(N__5095),
            .in3(N__5071),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9157),
            .ce(),
            .sr(N__8933));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_10_13_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_10_13_2 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_10_13_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_10_13_2  (
            .in0(N__4577),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4221),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9157),
            .ce(),
            .sr(N__8933));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_10_13_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_10_13_4 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_10_13_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_10_13_4  (
            .in0(N__4563),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9157),
            .ce(),
            .sr(N__8933));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_10_13_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_10_13_5 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_10_13_5 .LUT_INIT=16'b0011001000110000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_10_13_5  (
            .in0(N__4534),
            .in1(N__4576),
            .in2(N__4825),
            .in3(N__5070),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9157),
            .ce(),
            .sr(N__8933));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_10_13_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_10_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_10_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4546),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9157),
            .ce(),
            .sr(N__8933));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_14_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_14_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(N__4559),
            .in2(_gnd_net_),
            .in3(N__4545),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TACKn_obuft_RNO_LC_10_18_4.C_ON=1'b0;
    defparam TACKn_obuft_RNO_LC_10_18_4.SEQ_MODE=4'b0000;
    defparam TACKn_obuft_RNO_LC_10_18_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 TACKn_obuft_RNO_LC_10_18_4 (
            .in0(N__5044),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_886_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_6_5 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_6_5  (
            .in0(N__4780),
            .in1(N__6809),
            .in2(N__8587),
            .in3(N__4942),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_6_6 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_6_6  (
            .in0(N__6810),
            .in1(N__4507),
            .in2(N__4486),
            .in3(N__4483),
            .lcout(\U712_CHIP_RAM.N_313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(N__4716),
            .in2(_gnd_net_),
            .in3(N__4731),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_9_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_9_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__4870),
            .in2(_gnd_net_),
            .in3(N__4471),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__4699),
            .ce(),
            .sr(N__5983));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_9_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_9_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__4897),
            .in2(_gnd_net_),
            .in3(N__4468),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__4699),
            .ce(),
            .sr(N__5983));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_9_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_9_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__4909),
            .in2(_gnd_net_),
            .in3(N__4741),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__4699),
            .ce(),
            .sr(N__5983));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_9_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_9_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__4846),
            .in2(_gnd_net_),
            .in3(N__4738),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__4699),
            .ce(),
            .sr(N__5983));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_9_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_9_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__4884),
            .in2(_gnd_net_),
            .in3(N__4735),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__4699),
            .ce(),
            .sr(N__5983));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_9_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_9_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__4732),
            .in2(_gnd_net_),
            .in3(N__4720),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__4699),
            .ce(),
            .sr(N__5983));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_9_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_9_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__4717),
            .in2(_gnd_net_),
            .in3(N__4705),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__4699),
            .ce(),
            .sr(N__5983));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_9_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_9_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__4858),
            .in2(_gnd_net_),
            .in3(N__4702),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4699),
            .ce(),
            .sr(N__5983));
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_11_1 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_5_LC_11_11_1  (
            .in0(N__4650),
            .in1(N__4673),
            .in2(_gnd_net_),
            .in3(N__4690),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9148),
            .ce(),
            .sr(N__8937));
    defparam \U712_REG_SM.REG_TACK_LC_11_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_11_11_4 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_11_11_4  (
            .in0(N__4672),
            .in1(N__4649),
            .in2(N__4636),
            .in3(N__5107),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9148),
            .ce(),
            .sr(N__8937));
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_11_12_2 .C_ON=1'b0;
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_11_12_2 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_REG_SM.UDS_OUT_RNIUP9B_LC_11_12_2  (
            .in0(N__5940),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4612),
            .lcout(U712_REG_SM_un1_UDSn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_11_13_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_11_13_1 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_11_13_1  (
            .in0(N__8235),
            .in1(N__5087),
            .in2(N__4824),
            .in3(N__5060),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_305_i_0_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_13_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_13_2 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_13_2  (
            .in0(N__9018),
            .in1(_gnd_net_),
            .in2(N__4807),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.N_305_i_0_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_12_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_12_5_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_12_5_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_12_5_1  (
            .in0(N__4804),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9117),
            .ce(N__8636),
            .sr(N__8965));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_12_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_12_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_12_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4803),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9118),
            .ce(N__8727),
            .sr(N__8956));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_12_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_12_6_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_12_6_1  (
            .in0(N__4774),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9118),
            .ce(N__8727),
            .sr(N__8956));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_12_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_12_6_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_12_6_2  (
            .in0(N__4972),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9118),
            .ce(N__8727),
            .sr(N__8956));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_6_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_6_3  (
            .in0(N__8692),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9118),
            .ce(N__8727),
            .sr(N__8956));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_12_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_12_6_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_12_6_4  (
            .in0(N__4936),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9118),
            .ce(N__8727),
            .sr(N__8956));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_7_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_7_0  (
            .in0(N__4770),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9122),
            .ce(N__8635),
            .sr(N__8951));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_7_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_7_1  (
            .in0(N__5584),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9122),
            .ce(N__8635),
            .sr(N__8951));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4971),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9122),
            .ce(N__8635),
            .sr(N__8951));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_12_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_12_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_12_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_12_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5623),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9122),
            .ce(N__8635),
            .sr(N__8951));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4935),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9126),
            .ce(N__8641),
            .sr(N__8943));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_12_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_12_9_1 .LUT_INIT=16'b1111000111101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_12_9_1  (
            .in0(N__8112),
            .in1(N__7991),
            .in2(N__7848),
            .in3(N__7731),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_341_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_12_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_12_9_2 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_12_9_2  (
            .in0(N__7846),
            .in1(N__7765),
            .in2(N__4915),
            .in3(N__7382),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_12_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_12_9_3 .LUT_INIT=16'b1111100011111001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_12_9_3  (
            .in0(N__7383),
            .in1(N__7733),
            .in2(N__4912),
            .in3(N__7847),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_12_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_12_9_4 .LUT_INIT=16'b0001111101011111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_12_9_4  (
            .in0(N__4908),
            .in1(N__4896),
            .in2(N__4885),
            .in3(N__4869),
            .lcout(),
            .ltout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_12_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_12_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_12_9_5 .LUT_INIT=16'b1010111011111111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_12_9_5  (
            .in0(N__4857),
            .in1(N__4845),
            .in2(N__4834),
            .in3(N__4831),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9130),
            .ce(),
            .sr(N__8939));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_12_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_12_9_7 .LUT_INIT=16'b0101000010100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_12_9_7  (
            .in0(N__7381),
            .in1(_gnd_net_),
            .in2(N__7849),
            .in3(N__7732),
            .lcout(\U712_CHIP_RAM.N_403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_12_10_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_12_10_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_12_10_0  (
            .in0(N__7582),
            .in1(N__5198),
            .in2(_gnd_net_),
            .in3(N__6177),
            .lcout(\U712_BYTE_ENABLE.N_392 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_0_LC_12_10_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_0_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_0_LC_12_10_1 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_0_LC_12_10_1  (
            .in0(N__6178),
            .in1(_gnd_net_),
            .in2(N__5203),
            .in3(N__7583),
            .lcout(\U712_BYTE_ENABLE.N_388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_12_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_12_10_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_12_10_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_12_10_2  (
            .in0(N__5248),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5202),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9135),
            .ce(),
            .sr(N__8934));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_12_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_12_10_3 .LUT_INIT=16'b0101011100000011;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_12_10_3  (
            .in0(N__6813),
            .in1(N__5176),
            .in2(N__5143),
            .in3(N__5794),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9135),
            .ce(),
            .sr(N__8934));
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_12_12_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_12_12_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN6_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(N__5106),
            .in2(_gnd_net_),
            .in3(N__5955),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_12_13_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_12_13_1 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_12_13_1 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_LC_12_13_1  (
            .in0(N__8231),
            .in1(N__5094),
            .in2(_gnd_net_),
            .in3(N__5064),
            .lcout(TACK_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9152),
            .ce(N__5029),
            .sr(N__8929));
    defparam RESETn_ibuf_RNIM9SF_LC_12_17_2.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_17_2.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_17_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8236),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_4_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_4_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_4_1 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_4_1  (
            .in0(N__5014),
            .in1(N__5632),
            .in2(N__4993),
            .in3(N__6825),
            .lcout(\U712_CHIP_RAM.N_316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_5_1 .LUT_INIT=16'b0000101101011011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_5_1  (
            .in0(N__6776),
            .in1(N__5488),
            .in2(N__8588),
            .in3(N__5482),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_5_2 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_5_2  (
            .in0(N__5476),
            .in1(N__5455),
            .in2(N__5431),
            .in3(N__6780),
            .lcout(\U712_CHIP_RAM.N_311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_5_3 .LUT_INIT=16'b0000010111110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_5_3  (
            .in0(N__5428),
            .in1(N__5419),
            .in2(N__6814),
            .in3(N__8575),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_5_4 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_5_4  (
            .in0(N__5413),
            .in1(N__5395),
            .in2(N__5374),
            .in3(N__6781),
            .lcout(\U712_CHIP_RAM.N_312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_13_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_13_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_13_5_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_13_5_6  (
            .in0(N__8576),
            .in1(N__7099),
            .in2(N__8442),
            .in3(N__8328),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9119),
            .ce(N__6989),
            .sr(N__8968));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_13_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_13_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_13_6_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_13_6_2  (
            .in0(N__7094),
            .in1(N__5350),
            .in2(_gnd_net_),
            .in3(N__8431),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9123),
            .ce(N__6971),
            .sr(N__8966));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_13_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_13_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_13_6_3 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_13_6_3  (
            .in0(N__5323),
            .in1(N__6815),
            .in2(N__8586),
            .in3(N__8653),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_13_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_13_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_13_6_4 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_13_6_4  (
            .in0(N__6816),
            .in1(N__5317),
            .in2(N__5296),
            .in3(N__5293),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_314_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_6_5 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_13_6_5  (
            .in0(N__8430),
            .in1(_gnd_net_),
            .in2(N__5662),
            .in3(N__7095),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9123),
            .ce(N__6971),
            .sr(N__8966));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_13_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_13_7_1 .LUT_INIT=16'b0011000100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_13_7_1  (
            .in0(N__5596),
            .in1(N__8537),
            .in2(N__6773),
            .in3(N__5638),
            .lcout(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_13_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_13_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_13_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_13_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5622),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9127),
            .ce(N__8726),
            .sr(N__8957));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_13_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_13_7_3 .LUT_INIT=16'b0011000100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_13_7_3  (
            .in0(N__5551),
            .in1(N__8538),
            .in2(N__6774),
            .in3(N__5590),
            .lcout(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_13_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_13_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_13_7_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_13_7_4  (
            .in0(N__5580),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9127),
            .ce(N__8726),
            .sr(N__8957));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_7_5 .LUT_INIT=16'b0011000100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_7_5  (
            .in0(N__5494),
            .in1(N__8539),
            .in2(N__6775),
            .in3(N__5542),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_7_6 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_7_6  (
            .in0(N__6743),
            .in1(N__5536),
            .in2(N__5518),
            .in3(N__5515),
            .lcout(\U712_CHIP_RAM.N_317 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_13_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_13_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_13_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8800),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9127),
            .ce(N__8726),
            .sr(N__8957));
    defparam \U712_CHIP_RAM.DBDIR_LC_13_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_13_8_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_13_8_0 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_13_8_0  (
            .in0(N__6928),
            .in1(N__6413),
            .in2(_gnd_net_),
            .in3(N__6231),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9131),
            .ce(),
            .sr(N__8952));
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_13_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_13_8_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_13_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DBR_SYNC_0_LC_13_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5713),
            .lcout(U712_REG_SM_DBR_SYNC_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9131),
            .ce(),
            .sr(N__8952));
    defparam \U712_REG_SM.DBR_SYNC_1_LC_13_8_2 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_13_8_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_13_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.DBR_SYNC_1_LC_13_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5775),
            .lcout(U712_REG_SM_DBR_SYNC_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9131),
            .ce(),
            .sr(N__8952));
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_13_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_13_8_7 .LUT_INIT=16'b0101011100000010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_LC_13_8_7  (
            .in0(N__6202),
            .in1(N__6629),
            .in2(N__7740),
            .in3(N__6747),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9131),
            .ce(),
            .sr(N__8952));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI32IV_LC_13_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI32IV_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI32IV_LC_13_9_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNI32IV_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(N__8230),
            .in2(_gnd_net_),
            .in3(N__6619),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIT6BC2_2_LC_13_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIT6BC2_2_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIT6BC2_2_LC_13_9_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIT6BC2_2_LC_13_9_1  (
            .in0(N__7370),
            .in1(N__7696),
            .in2(N__5692),
            .in3(N__8088),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFP3R8_2_LC_13_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFP3R8_2_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFP3R8_2_LC_13_9_2 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIFP3R8_2_LC_13_9_2  (
            .in0(N__6245),
            .in1(N__6486),
            .in2(N__5689),
            .in3(N__6253),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_13_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_13_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_13_9_3 .LUT_INIT=16'b0011000010111010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_13_9_3  (
            .in0(N__5686),
            .in1(N__7572),
            .in2(N__6630),
            .in3(N__5677),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9139),
            .ce(),
            .sr(N__8946));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_13_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_13_9_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_13_9_4  (
            .in0(N__6246),
            .in1(N__6620),
            .in2(_gnd_net_),
            .in3(N__6487),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_13_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_13_9_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_13_9_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_13_9_5  (
            .in0(N__5676),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9139),
            .ce(),
            .sr(N__8946));
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_13_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_13_9_6 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_13_9_6  (
            .in0(N__9020),
            .in1(N__5685),
            .in2(_gnd_net_),
            .in3(N__5675),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIKEL61_LC_13_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIKEL61_LC_13_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIKEL61_LC_13_9_7 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIKEL61_LC_13_9_7  (
            .in0(N__5793),
            .in1(N__5771),
            .in2(_gnd_net_),
            .in3(N__5748),
            .lcout(\U712_CHIP_RAM.N_285 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_13_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_13_10_0 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_13_10_0  (
            .in0(N__8148),
            .in1(N__7373),
            .in2(_gnd_net_),
            .in3(N__6492),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_13_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_13_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_13_10_1 .LUT_INIT=16'b1111111000110010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_13_10_1  (
            .in0(N__5737),
            .in1(N__6285),
            .in2(N__5731),
            .in3(N__8524),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9144),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_2_LC_13_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_2_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_2_LC_13_10_2 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_2_LC_13_10_2  (
            .in0(N__7976),
            .in1(N__8089),
            .in2(N__7827),
            .in3(N__7371),
            .lcout(\U712_CHIP_RAM.N_421 ),
            .ltout(\U712_CHIP_RAM.N_421_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMMGI5_2_LC_13_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMMGI5_2_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMMGI5_2_LC_13_10_3 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIMMGI5_2_LC_13_10_3  (
            .in0(N__6124),
            .in1(_gnd_net_),
            .in2(N__5728),
            .in3(N__6510),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_293_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJ42D8_0_LC_13_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJ42D8_0_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJ42D8_0_LC_13_10_4 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIJ42D8_0_LC_13_10_4  (
            .in0(N__7720),
            .in1(N__9019),
            .in2(N__5725),
            .in3(N__7245),
            .lcout(\U712_CHIP_RAM.N_309 ),
            .ltout(\U712_CHIP_RAM.N_309_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_13_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_13_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_13_10_5 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_13_10_5  (
            .in0(N__7374),
            .in1(_gnd_net_),
            .in2(N__5722),
            .in3(N__7721),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9144),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_13_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_13_10_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_13_10_6  (
            .in0(N__5719),
            .in1(N__8037),
            .in2(_gnd_net_),
            .in3(N__7244),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_1_LC_13_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_1_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_1_LC_13_10_7 .LUT_INIT=16'b0010000100000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_RNO_1_LC_13_10_7  (
            .in0(N__7372),
            .in1(N__7757),
            .in2(N__7735),
            .in3(N__7813),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_0_a2_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_LC_13_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_LC_13_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_LC_13_11_6 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_LC_13_11_6  (
            .in0(N__6100),
            .in1(N__5962),
            .in2(_gnd_net_),
            .in3(N__6547),
            .lcout(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9149),
            .ce(),
            .sr(N__8938));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_13_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_13_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_13_11_7 .LUT_INIT=16'b1000101110001000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_13_11_7  (
            .in0(N__5956),
            .in1(N__6442),
            .in2(N__7407),
            .in3(N__6790),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9149),
            .ce(),
            .sr(N__8938));
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_13_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_13_12_0 .LUT_INIT=16'b0111011101110111;
    LogicCell40 \U712_REG_SM.LDS_OUT_RNIL31J_LC_13_12_0  (
            .in0(N__5944),
            .in1(N__5923),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(U712_REG_SM_un1_LDSn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_14_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_14_4_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_14_4_5 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_14_4_5  (
            .in0(N__5887),
            .in1(N__7100),
            .in2(_gnd_net_),
            .in3(N__8435),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9120),
            .ce(N__6978),
            .sr(N__8980));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_14_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_14_5_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_14_5_0 .LUT_INIT=16'b1010101010100011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_14_5_0  (
            .in0(N__5863),
            .in1(N__8584),
            .in2(N__7108),
            .in3(N__8419),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9124),
            .ce(N__6985),
            .sr(N__8976));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_14_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_14_5_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_14_5_1 .LUT_INIT=16'b1111110100000001;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_14_5_1  (
            .in0(N__8583),
            .in1(N__7103),
            .in2(N__8436),
            .in3(N__5839),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9124),
            .ce(N__6985),
            .sr(N__8976));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI9T531_3_LC_14_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI9T531_3_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI9T531_3_LC_14_6_0 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI9T531_3_LC_14_6_0  (
            .in0(N__7077),
            .in1(N__8321),
            .in2(N__8585),
            .in3(N__5979),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_CMA31_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIV62J1_3_LC_14_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIV62J1_3_LC_14_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIV62J1_3_LC_14_6_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIV62J1_3_LC_14_6_1  (
            .in0(N__9029),
            .in1(_gnd_net_),
            .in2(N__5812),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_CMA31_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_6_3 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_6_3  (
            .in0(N__5809),
            .in1(N__6082),
            .in2(N__6076),
            .in3(N__6791),
            .lcout(\U712_CHIP_RAM.N_315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_2_LC_14_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_2_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_2_LC_14_6_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_2_LC_14_6_5  (
            .in0(N__6496),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7408),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_493_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_1_LC_14_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_1_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_1_LC_14_6_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_1_LC_14_6_6  (
            .in0(N__7246),
            .in1(N__7734),
            .in2(N__6055),
            .in3(N__8038),
            .lcout(),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_14_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_14_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_14_6_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_14_6_7  (
            .in0(N__9030),
            .in1(_gnd_net_),
            .in2(N__6052),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_7_3 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_14_7_3  (
            .in0(N__6049),
            .in1(_gnd_net_),
            .in2(N__8426),
            .in3(N__7076),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9132),
            .ce(N__6993),
            .sr(N__8967));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_14_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_14_7_5 .LUT_INIT=16'b0000111101011111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_14_7_5  (
            .in0(N__8398),
            .in1(_gnd_net_),
            .in2(N__8562),
            .in3(N__7075),
            .lcout(\U712_CHIP_RAM.CMA_5_i_0_8 ),
            .ltout(\U712_CHIP_RAM.CMA_5_i_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_7_6 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_14_7_6  (
            .in0(N__8278),
            .in1(N__6028),
            .in2(N__6007),
            .in3(N__6748),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9132),
            .ce(N__6993),
            .sr(N__8967));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNITDMK_3_LC_14_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNITDMK_3_LC_14_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNITDMK_3_LC_14_7_7 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_RNITDMK_3_LC_14_7_7  (
            .in0(N__8397),
            .in1(N__8311),
            .in2(N__8561),
            .in3(N__7074),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_3_LC_14_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_3_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_3_LC_14_8_0 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_3_LC_14_8_0  (
            .in0(N__6130),
            .in1(N__7240),
            .in2(N__6232),
            .in3(N__7978),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_14_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_14_8_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_14_8_1  (
            .in0(N__9023),
            .in1(_gnd_net_),
            .in2(N__5965),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI7Q5U5_LC_14_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI7Q5U5_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI7Q5U5_LC_14_8_2 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNI7Q5U5_LC_14_8_2  (
            .in0(N__6493),
            .in1(N__6247),
            .in2(N__6099),
            .in3(N__6624),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIAEJU_LC_14_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIAEJU_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIAEJU_LC_14_8_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIAEJU_LC_14_8_3  (
            .in0(N__6625),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7722),
            .lcout(),
            .ltout(\U712_CHIP_RAM.DMA_CYCLE_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_LC_14_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_14_8_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_14_8_4 .LUT_INIT=16'b0101111111001100;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_14_8_4  (
            .in0(N__6217),
            .in1(N__6151),
            .in2(N__6205),
            .in3(N__6201),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9140),
            .ce(),
            .sr(N__8958));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISB5T1_2_LC_14_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISB5T1_2_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISB5T1_2_LC_14_8_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNISB5T1_2_LC_14_8_5  (
            .in0(N__7699),
            .in1(N__7388),
            .in2(N__8115),
            .in3(N__6494),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_2_LC_14_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_2_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_2_LC_14_8_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_2_LC_14_8_7  (
            .in0(N__7977),
            .in1(N__7389),
            .in2(N__8116),
            .in3(N__6495),
            .lcout(\U712_CHIP_RAM.N_427 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3F0BF_0_LC_14_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3F0BF_0_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3F0BF_0_LC_14_9_0 .LUT_INIT=16'b1111111111001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI3F0BF_0_LC_14_9_0  (
            .in0(N__6115),
            .in1(N__8122),
            .in2(N__6514),
            .in3(N__6109),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_sbtinv_3_LC_14_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_sbtinv_3_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_sbtinv_3_LC_14_9_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_sbtinv_3_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6103),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_14_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_14_9_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_14_9_2  (
            .in0(N__7359),
            .in1(N__8016),
            .in2(N__7239),
            .in3(N__7694),
            .lcout(\U712_CHIP_RAM.N_296 ),
            .ltout(\U712_CHIP_RAM.N_296_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_14_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_14_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_14_9_3 .LUT_INIT=16'b0001001000010011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_14_9_3  (
            .in0(N__7695),
            .in1(N__6298),
            .in2(N__6316),
            .in3(N__6313),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9145),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_14_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_14_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_14_9_4 .LUT_INIT=16'b1111111000001110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_14_9_4  (
            .in0(N__6307),
            .in1(N__7441),
            .in2(N__6286),
            .in3(N__7073),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9145),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_14_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_14_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_14_9_5 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_14_9_5  (
            .in0(N__7384),
            .in1(N__7726),
            .in2(N__8114),
            .in3(N__6296),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9145),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_14_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_14_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_14_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_14_9_6  (
            .in0(N__6297),
            .in1(N__7899),
            .in2(_gnd_net_),
            .in3(N__7990),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9145),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_14_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_14_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_14_9_7 .LUT_INIT=16'b1111001111100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_14_9_7  (
            .in0(N__7599),
            .in1(N__6284),
            .in2(N__8425),
            .in3(N__7423),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9145),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_14_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_14_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_14_10_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_14_10_3  (
            .in0(N__6268),
            .in1(N__7579),
            .in2(_gnd_net_),
            .in3(N__6792),
            .lcout(\U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9150),
            .ce(),
            .sr(N__8947));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_14_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_14_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_14_10_4 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_14_10_4  (
            .in0(N__7808),
            .in1(N__7238),
            .in2(_gnd_net_),
            .in3(N__6562),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9150),
            .ce(),
            .sr(N__8947));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83_2_LC_14_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83_2_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83_2_LC_14_10_5 .LUT_INIT=16'b0000000000110111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83_2_LC_14_10_5  (
            .in0(N__7358),
            .in1(N__8087),
            .in2(N__7730),
            .in3(N__7221),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISSMN4_3_LC_14_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISSMN4_3_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISSMN4_3_LC_14_10_6 .LUT_INIT=16'b0000000010001010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNISSMN4_3_LC_14_10_6  (
            .in0(N__8225),
            .in1(N__7975),
            .in2(N__6256),
            .in3(N__6478),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_14_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_14_10_7 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_14_10_7  (
            .in0(N__6545),
            .in1(N__6528),
            .in2(_gnd_net_),
            .in3(N__7807),
            .lcout(\U712_CHIP_RAM.N_282 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI7MV4_LC_14_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI7MV4_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI7MV4_LC_14_11_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI7MV4_LC_14_11_2  (
            .in0(_gnd_net_),
            .in1(N__6546),
            .in2(_gnd_net_),
            .in3(N__6529),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER46 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER46_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVE5T1_LC_14_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVE5T1_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVE5T1_LC_14_11_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVE5T1_LC_14_11_3  (
            .in0(N__8017),
            .in1(N__7360),
            .in2(N__6517),
            .in3(N__7809),
            .lcout(\U712_CHIP_RAM.N_420 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_14_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_14_11_6 .LUT_INIT=16'b1111111110110111;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_14_11_6  (
            .in0(N__7361),
            .in1(N__8113),
            .in2(N__7741),
            .in3(N__6491),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_a5_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_14_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_14_11_7 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_14_11_7  (
            .in0(_gnd_net_),
            .in1(N__7992),
            .in2(N__6445),
            .in3(N__7236),
            .lcout(\U712_CHIP_RAM.N_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DRDDIR_i_LC_14_13_2 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_i_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_i_LC_14_13_2 .LUT_INIT=16'b0011000010111010;
    LogicCell40 \U712_BUFFERS.DRDDIR_i_LC_14_13_2  (
            .in0(N__7581),
            .in1(N__6874),
            .in2(N__7513),
            .in3(N__6426),
            .lcout(N_218),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RASn_LC_15_3_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_15_3_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_15_3_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_15_3_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7107),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9121),
            .ce(),
            .sr(N__8984));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_15_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_15_4_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_15_4_2 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_15_4_2  (
            .in0(N__8737),
            .in1(N__6823),
            .in2(N__8595),
            .in3(N__8767),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_15_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_15_4_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_15_4_3 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_15_4_3  (
            .in0(N__6824),
            .in1(N__6361),
            .in2(N__6340),
            .in3(N__6337),
            .lcout(\U712_CHIP_RAM.N_318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_15_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_15_5_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_15_5_0 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_15_5_0  (
            .in0(N__7183),
            .in1(N__7165),
            .in2(N__7453),
            .in3(N__6812),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9128),
            .ce(N__6994),
            .sr(N__8981));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_15_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_15_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_15_5_2 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_15_5_2  (
            .in0(N__7135),
            .in1(_gnd_net_),
            .in2(N__8443),
            .in3(N__7102),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9128),
            .ce(N__6994),
            .sr(N__8981));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_15_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_15_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_15_5_6 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_15_5_6  (
            .in0(N__8437),
            .in1(N__7101),
            .in2(_gnd_net_),
            .in3(N__7021),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9128),
            .ce(N__6994),
            .sr(N__8981));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_15_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_15_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_15_6_0 .LUT_INIT=16'b0100111101000100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_15_6_0  (
            .in0(N__6927),
            .in1(N__7545),
            .in2(N__6889),
            .in3(N__6811),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9133),
            .ce(N__6643),
            .sr(N__8977));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_15_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_15_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_15_7_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_15_7_0  (
            .in0(_gnd_net_),
            .in1(N__6634),
            .in2(_gnd_net_),
            .in3(N__7739),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9141),
            .ce(N__6592),
            .sr(N__8969));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_3_LC_15_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_3_LC_15_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_3_LC_15_8_1 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_3_LC_15_8_1  (
            .in0(N__7600),
            .in1(N__7411),
            .in2(N__8152),
            .in3(N__7288),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9146),
            .ce(N__6577),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_15_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_15_8_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_15_8_4  (
            .in0(N__7410),
            .in1(N__8099),
            .in2(N__7993),
            .in3(N__6553),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_0_i_a2_1_0_a2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_15_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_15_8_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_15_8_6  (
            .in0(N__7409),
            .in1(N__7716),
            .in2(_gnd_net_),
            .in3(N__8098),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIO6AQ_LC_15_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIO6AQ_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIO6AQ_LC_15_9_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIO6AQ_LC_15_9_0  (
            .in0(_gnd_net_),
            .in1(N__7700),
            .in2(_gnd_net_),
            .in3(N__7819),
            .lcout(\U712_CHIP_RAM.N_284 ),
            .ltout(\U712_CHIP_RAM.N_284_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_15_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_15_9_1 .LUT_INIT=16'b1111111010101111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_15_9_1  (
            .in0(N__8141),
            .in1(N__7413),
            .in2(N__7444),
            .in3(N__8036),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_15_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_15_9_2 .LUT_INIT=16'b0101000001110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_15_9_2  (
            .in0(N__7412),
            .in1(N__7701),
            .in2(N__7839),
            .in3(N__7435),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_15_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_15_9_3 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_15_9_3  (
            .in0(N__8226),
            .in1(N__8035),
            .in2(N__7426),
            .in3(N__7237),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_15_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_15_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_15_9_4 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_15_9_4  (
            .in0(N__7898),
            .in1(N__7920),
            .in2(N__9031),
            .in3(N__7989),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9151),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_15_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_15_9_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_15_9_5  (
            .in0(N__7988),
            .in1(N__7869),
            .in2(N__7921),
            .in3(N__7897),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c6 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_15_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_15_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_15_9_6 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_15_9_6  (
            .in0(N__9027),
            .in1(_gnd_net_),
            .in2(N__7417),
            .in3(N__7273),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9151),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_3_LC_15_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_3_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_3_LC_15_9_7 .LUT_INIT=16'b1111010100101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_3_LC_15_9_7  (
            .in0(N__7702),
            .in1(N__7414),
            .in2(N__7838),
            .in3(N__8034),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_15_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_15_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_15_10_0 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_15_10_0  (
            .in0(N__9022),
            .in1(N__7272),
            .in2(N__7282),
            .in3(N__7257),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9153),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_15_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_15_10_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_15_10_1  (
            .in0(N__7271),
            .in1(N__7862),
            .in2(N__7258),
            .in3(N__7915),
            .lcout(\U712_CHIP_RAM.N_274 ),
            .ltout(\U712_CHIP_RAM.N_274_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_15_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_15_10_2 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_15_10_2  (
            .in0(N__8224),
            .in1(_gnd_net_),
            .in2(N__8155),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_337 ),
            .ltout(\U712_CHIP_RAM.N_337_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITDHQ2_0_LC_15_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITDHQ2_0_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITDHQ2_0_LC_15_10_3 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITDHQ2_0_LC_15_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8125),
            .in3(N__7697),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_15_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_15_10_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_15_10_4  (
            .in0(_gnd_net_),
            .in1(N__7973),
            .in2(_gnd_net_),
            .in3(N__8086),
            .lcout(\U712_CHIP_RAM.N_271 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_5_LC_15_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_5_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_5_LC_15_10_5 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_5_LC_15_10_5  (
            .in0(N__7974),
            .in1(N__7916),
            .in2(N__7873),
            .in3(N__7900),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_15_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_15_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_15_10_6 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_15_10_6  (
            .in0(N__9021),
            .in1(_gnd_net_),
            .in2(N__7876),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9153),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVS9V_LC_15_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVS9V_LC_15_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVS9V_LC_15_10_7 .LUT_INIT=16'b0101010100100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVS9V_LC_15_10_7  (
            .in0(N__7823),
            .in1(N__7761),
            .in2(_gnd_net_),
            .in3(N__7698),
            .lcout(\U712_CHIP_RAM.N_303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_0_a2_LC_15_13_1 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_0_a2_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_0_a2_LC_15_13_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_0_a2_0_a2_LC_15_13_1  (
            .in0(N__7580),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7512),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_5_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8761),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9134),
            .ce(N__8640),
            .sr(N__8983));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8796),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9134),
            .ce(N__8640),
            .sr(N__8983));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_16_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_16_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_16_6_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_16_6_4  (
            .in0(N__8757),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9142),
            .ce(N__8728),
            .sr(N__8982));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_16_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_16_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_16_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_16_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8688),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9147),
            .ce(N__8622),
            .sr(N__8978));
    defparam \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_16_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_16_8_2 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_16_8_2  (
            .in0(N__9028),
            .in1(N__9169),
            .in2(_gnd_net_),
            .in3(N__9180),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CASn_LC_17_2_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_17_2_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_17_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_17_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8596),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9125),
            .ce(),
            .sr(N__8987));
    defparam \U712_CHIP_RAM.WEn_LC_17_3_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_17_3_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_17_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_17_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8441),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9129),
            .ce(),
            .sr(N__8986));
    defparam \U712_CHIP_RAM.CRCSn_LC_17_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_17_5_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_17_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_17_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8329),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9143),
            .ce(),
            .sr(N__8985));
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_17_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_17_8_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_17_8_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_0_LC_17_8_3  (
            .in0(_gnd_net_),
            .in1(N__8277),
            .in2(_gnd_net_),
            .in3(N__8248),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9154),
            .ce(),
            .sr(N__8979));
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_17_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_17_8_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_17_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_1_LC_17_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9181),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9154),
            .ce(),
            .sr(N__8979));
    defparam CONSTANT_ONE_LUT4_LC_22_4_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_22_4_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_22_4_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_22_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U712_TOP

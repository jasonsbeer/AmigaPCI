// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 7 2025 10:58:53

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U409_TOP" view "INTERFACE"

module U409_TOP (
    TT,
    TM,
    A,
    D,
    RESETn,
    OVL,
    CONFIGENn,
    PIO_S0,
    PORTSIZE,
    TICK60,
    CIACS0n,
    CPUCONFn,
    CLK6,
    CLK_CIA,
    BUFENn,
    AUTOBOOT,
    RnW,
    PIO_P2,
    CIACS1n,
    BRIDGE_ENn,
    PIO_S1,
    ATA_MODE_S,
    PIO_P0,
    TICK50,
    TCIn,
    TBIn,
    RAMSPACEn,
    CLK40_IN,
    CLK28_IN,
    REGSPACEn,
    TSn,
    RTC_ENn,
    PIO_S2,
    ATA_ENn,
    TACKn,
    ATA_MODE_P,
    ROMENn,
    PIO_P1);

    input [1:0] TT;
    input [1:0] TM;
    input [31:1] A;
    inout [7:4] D;
    input RESETn;
    input OVL;
    output CONFIGENn;
    output PIO_S0;
    output PORTSIZE;
    output TICK60;
    output CIACS0n;
    input CPUCONFn;
    input CLK6;
    output CLK_CIA;
    output BUFENn;
    input AUTOBOOT;
    input RnW;
    output PIO_P2;
    output CIACS1n;
    output BRIDGE_ENn;
    output PIO_S1;
    input ATA_MODE_S;
    output PIO_P0;
    output TICK50;
    output TCIn;
    output TBIn;
    output RAMSPACEn;
    input CLK40_IN;
    input CLK28_IN;
    output REGSPACEn;
    input TSn;
    output RTC_ENn;
    output PIO_S2;
    output ATA_ENn;
    inout TACKn;
    input ATA_MODE_P;
    output ROMENn;
    output PIO_P1;

    wire N__11402;
    wire N__11401;
    wire N__11400;
    wire N__11392;
    wire N__11391;
    wire N__11390;
    wire N__11382;
    wire N__11381;
    wire N__11380;
    wire N__11371;
    wire N__11370;
    wire N__11369;
    wire N__11362;
    wire N__11361;
    wire N__11360;
    wire N__11353;
    wire N__11352;
    wire N__11351;
    wire N__11344;
    wire N__11343;
    wire N__11342;
    wire N__11335;
    wire N__11334;
    wire N__11333;
    wire N__11326;
    wire N__11325;
    wire N__11324;
    wire N__11317;
    wire N__11316;
    wire N__11315;
    wire N__11308;
    wire N__11307;
    wire N__11306;
    wire N__11299;
    wire N__11298;
    wire N__11297;
    wire N__11290;
    wire N__11289;
    wire N__11288;
    wire N__11281;
    wire N__11280;
    wire N__11279;
    wire N__11272;
    wire N__11271;
    wire N__11270;
    wire N__11263;
    wire N__11262;
    wire N__11261;
    wire N__11254;
    wire N__11253;
    wire N__11252;
    wire N__11245;
    wire N__11244;
    wire N__11243;
    wire N__11236;
    wire N__11235;
    wire N__11234;
    wire N__11227;
    wire N__11226;
    wire N__11225;
    wire N__11218;
    wire N__11217;
    wire N__11216;
    wire N__11209;
    wire N__11208;
    wire N__11207;
    wire N__11200;
    wire N__11199;
    wire N__11198;
    wire N__11191;
    wire N__11190;
    wire N__11189;
    wire N__11182;
    wire N__11181;
    wire N__11180;
    wire N__11173;
    wire N__11172;
    wire N__11171;
    wire N__11164;
    wire N__11163;
    wire N__11162;
    wire N__11155;
    wire N__11154;
    wire N__11153;
    wire N__11146;
    wire N__11145;
    wire N__11144;
    wire N__11137;
    wire N__11136;
    wire N__11135;
    wire N__11128;
    wire N__11127;
    wire N__11126;
    wire N__11119;
    wire N__11118;
    wire N__11117;
    wire N__11110;
    wire N__11109;
    wire N__11108;
    wire N__11101;
    wire N__11100;
    wire N__11099;
    wire N__11092;
    wire N__11091;
    wire N__11090;
    wire N__11083;
    wire N__11082;
    wire N__11081;
    wire N__11074;
    wire N__11073;
    wire N__11072;
    wire N__11065;
    wire N__11064;
    wire N__11063;
    wire N__11056;
    wire N__11055;
    wire N__11054;
    wire N__11047;
    wire N__11046;
    wire N__11045;
    wire N__11038;
    wire N__11037;
    wire N__11036;
    wire N__11029;
    wire N__11028;
    wire N__11027;
    wire N__11020;
    wire N__11019;
    wire N__11018;
    wire N__11011;
    wire N__11010;
    wire N__11009;
    wire N__11002;
    wire N__11001;
    wire N__11000;
    wire N__10993;
    wire N__10992;
    wire N__10991;
    wire N__10984;
    wire N__10983;
    wire N__10982;
    wire N__10975;
    wire N__10974;
    wire N__10973;
    wire N__10966;
    wire N__10965;
    wire N__10964;
    wire N__10957;
    wire N__10956;
    wire N__10955;
    wire N__10948;
    wire N__10947;
    wire N__10946;
    wire N__10939;
    wire N__10938;
    wire N__10937;
    wire N__10930;
    wire N__10929;
    wire N__10928;
    wire N__10921;
    wire N__10920;
    wire N__10919;
    wire N__10912;
    wire N__10911;
    wire N__10910;
    wire N__10903;
    wire N__10902;
    wire N__10901;
    wire N__10894;
    wire N__10893;
    wire N__10892;
    wire N__10885;
    wire N__10884;
    wire N__10883;
    wire N__10876;
    wire N__10875;
    wire N__10874;
    wire N__10867;
    wire N__10866;
    wire N__10865;
    wire N__10858;
    wire N__10857;
    wire N__10856;
    wire N__10849;
    wire N__10848;
    wire N__10847;
    wire N__10840;
    wire N__10839;
    wire N__10838;
    wire N__10831;
    wire N__10830;
    wire N__10829;
    wire N__10822;
    wire N__10821;
    wire N__10820;
    wire N__10813;
    wire N__10812;
    wire N__10811;
    wire N__10804;
    wire N__10803;
    wire N__10802;
    wire N__10785;
    wire N__10782;
    wire N__10779;
    wire N__10778;
    wire N__10777;
    wire N__10776;
    wire N__10775;
    wire N__10774;
    wire N__10773;
    wire N__10772;
    wire N__10761;
    wire N__10754;
    wire N__10749;
    wire N__10748;
    wire N__10747;
    wire N__10746;
    wire N__10745;
    wire N__10742;
    wire N__10741;
    wire N__10740;
    wire N__10739;
    wire N__10730;
    wire N__10721;
    wire N__10716;
    wire N__10715;
    wire N__10714;
    wire N__10713;
    wire N__10712;
    wire N__10709;
    wire N__10706;
    wire N__10705;
    wire N__10702;
    wire N__10701;
    wire N__10700;
    wire N__10697;
    wire N__10688;
    wire N__10683;
    wire N__10678;
    wire N__10671;
    wire N__10668;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10656;
    wire N__10655;
    wire N__10654;
    wire N__10653;
    wire N__10652;
    wire N__10651;
    wire N__10650;
    wire N__10649;
    wire N__10648;
    wire N__10629;
    wire N__10626;
    wire N__10623;
    wire N__10620;
    wire N__10619;
    wire N__10618;
    wire N__10615;
    wire N__10612;
    wire N__10609;
    wire N__10606;
    wire N__10605;
    wire N__10602;
    wire N__10599;
    wire N__10598;
    wire N__10595;
    wire N__10592;
    wire N__10589;
    wire N__10586;
    wire N__10583;
    wire N__10578;
    wire N__10575;
    wire N__10570;
    wire N__10567;
    wire N__10564;
    wire N__10561;
    wire N__10554;
    wire N__10551;
    wire N__10550;
    wire N__10547;
    wire N__10544;
    wire N__10539;
    wire N__10538;
    wire N__10535;
    wire N__10532;
    wire N__10527;
    wire N__10526;
    wire N__10525;
    wire N__10524;
    wire N__10521;
    wire N__10518;
    wire N__10515;
    wire N__10512;
    wire N__10509;
    wire N__10500;
    wire N__10499;
    wire N__10496;
    wire N__10493;
    wire N__10488;
    wire N__10485;
    wire N__10482;
    wire N__10479;
    wire N__10476;
    wire N__10475;
    wire N__10472;
    wire N__10469;
    wire N__10464;
    wire N__10461;
    wire N__10458;
    wire N__10455;
    wire N__10454;
    wire N__10451;
    wire N__10448;
    wire N__10443;
    wire N__10440;
    wire N__10437;
    wire N__10434;
    wire N__10431;
    wire N__10430;
    wire N__10427;
    wire N__10424;
    wire N__10419;
    wire N__10418;
    wire N__10415;
    wire N__10412;
    wire N__10407;
    wire N__10406;
    wire N__10403;
    wire N__10400;
    wire N__10395;
    wire N__10392;
    wire N__10389;
    wire N__10386;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10374;
    wire N__10371;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10359;
    wire N__10356;
    wire N__10353;
    wire N__10352;
    wire N__10351;
    wire N__10350;
    wire N__10349;
    wire N__10348;
    wire N__10345;
    wire N__10344;
    wire N__10337;
    wire N__10334;
    wire N__10327;
    wire N__10320;
    wire N__10319;
    wire N__10318;
    wire N__10317;
    wire N__10316;
    wire N__10313;
    wire N__10312;
    wire N__10311;
    wire N__10308;
    wire N__10301;
    wire N__10298;
    wire N__10293;
    wire N__10284;
    wire N__10283;
    wire N__10282;
    wire N__10275;
    wire N__10272;
    wire N__10269;
    wire N__10268;
    wire N__10267;
    wire N__10266;
    wire N__10263;
    wire N__10260;
    wire N__10255;
    wire N__10248;
    wire N__10247;
    wire N__10246;
    wire N__10245;
    wire N__10244;
    wire N__10241;
    wire N__10236;
    wire N__10231;
    wire N__10224;
    wire N__10223;
    wire N__10222;
    wire N__10221;
    wire N__10218;
    wire N__10215;
    wire N__10210;
    wire N__10203;
    wire N__10200;
    wire N__10197;
    wire N__10194;
    wire N__10191;
    wire N__10188;
    wire N__10185;
    wire N__10182;
    wire N__10179;
    wire N__10176;
    wire N__10173;
    wire N__10172;
    wire N__10169;
    wire N__10166;
    wire N__10161;
    wire N__10158;
    wire N__10155;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10143;
    wire N__10142;
    wire N__10139;
    wire N__10136;
    wire N__10131;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10123;
    wire N__10118;
    wire N__10115;
    wire N__10110;
    wire N__10109;
    wire N__10106;
    wire N__10103;
    wire N__10098;
    wire N__10097;
    wire N__10094;
    wire N__10091;
    wire N__10086;
    wire N__10083;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10071;
    wire N__10068;
    wire N__10065;
    wire N__10062;
    wire N__10059;
    wire N__10056;
    wire N__10055;
    wire N__10050;
    wire N__10047;
    wire N__10044;
    wire N__10043;
    wire N__10038;
    wire N__10035;
    wire N__10032;
    wire N__10031;
    wire N__10030;
    wire N__10027;
    wire N__10022;
    wire N__10017;
    wire N__10016;
    wire N__10013;
    wire N__10012;
    wire N__10009;
    wire N__10004;
    wire N__9999;
    wire N__9998;
    wire N__9997;
    wire N__9994;
    wire N__9989;
    wire N__9984;
    wire N__9981;
    wire N__9978;
    wire N__9977;
    wire N__9974;
    wire N__9973;
    wire N__9972;
    wire N__9969;
    wire N__9966;
    wire N__9961;
    wire N__9958;
    wire N__9951;
    wire N__9948;
    wire N__9945;
    wire N__9944;
    wire N__9941;
    wire N__9938;
    wire N__9933;
    wire N__9932;
    wire N__9929;
    wire N__9926;
    wire N__9921;
    wire N__9918;
    wire N__9915;
    wire N__9914;
    wire N__9911;
    wire N__9908;
    wire N__9903;
    wire N__9900;
    wire N__9897;
    wire N__9894;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9882;
    wire N__9881;
    wire N__9880;
    wire N__9879;
    wire N__9878;
    wire N__9877;
    wire N__9874;
    wire N__9873;
    wire N__9866;
    wire N__9861;
    wire N__9856;
    wire N__9849;
    wire N__9848;
    wire N__9847;
    wire N__9846;
    wire N__9845;
    wire N__9844;
    wire N__9843;
    wire N__9838;
    wire N__9835;
    wire N__9826;
    wire N__9823;
    wire N__9816;
    wire N__9815;
    wire N__9814;
    wire N__9813;
    wire N__9810;
    wire N__9807;
    wire N__9804;
    wire N__9803;
    wire N__9802;
    wire N__9801;
    wire N__9790;
    wire N__9787;
    wire N__9784;
    wire N__9781;
    wire N__9774;
    wire N__9771;
    wire N__9768;
    wire N__9767;
    wire N__9764;
    wire N__9761;
    wire N__9756;
    wire N__9753;
    wire N__9750;
    wire N__9747;
    wire N__9744;
    wire N__9741;
    wire N__9738;
    wire N__9735;
    wire N__9732;
    wire N__9729;
    wire N__9728;
    wire N__9725;
    wire N__9722;
    wire N__9717;
    wire N__9714;
    wire N__9711;
    wire N__9708;
    wire N__9705;
    wire N__9702;
    wire N__9699;
    wire N__9696;
    wire N__9693;
    wire N__9690;
    wire N__9689;
    wire N__9688;
    wire N__9685;
    wire N__9682;
    wire N__9679;
    wire N__9672;
    wire N__9669;
    wire N__9666;
    wire N__9663;
    wire N__9660;
    wire N__9657;
    wire N__9654;
    wire N__9651;
    wire N__9648;
    wire N__9647;
    wire N__9644;
    wire N__9641;
    wire N__9636;
    wire N__9635;
    wire N__9632;
    wire N__9629;
    wire N__9624;
    wire N__9621;
    wire N__9618;
    wire N__9617;
    wire N__9614;
    wire N__9611;
    wire N__9606;
    wire N__9603;
    wire N__9600;
    wire N__9597;
    wire N__9594;
    wire N__9591;
    wire N__9588;
    wire N__9585;
    wire N__9582;
    wire N__9581;
    wire N__9578;
    wire N__9575;
    wire N__9570;
    wire N__9567;
    wire N__9564;
    wire N__9561;
    wire N__9558;
    wire N__9555;
    wire N__9552;
    wire N__9549;
    wire N__9548;
    wire N__9547;
    wire N__9544;
    wire N__9541;
    wire N__9538;
    wire N__9531;
    wire N__9528;
    wire N__9525;
    wire N__9524;
    wire N__9521;
    wire N__9518;
    wire N__9513;
    wire N__9510;
    wire N__9507;
    wire N__9504;
    wire N__9503;
    wire N__9500;
    wire N__9497;
    wire N__9492;
    wire N__9489;
    wire N__9486;
    wire N__9485;
    wire N__9482;
    wire N__9479;
    wire N__9474;
    wire N__9471;
    wire N__9470;
    wire N__9467;
    wire N__9464;
    wire N__9459;
    wire N__9456;
    wire N__9453;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9438;
    wire N__9435;
    wire N__9432;
    wire N__9429;
    wire N__9426;
    wire N__9425;
    wire N__9424;
    wire N__9421;
    wire N__9420;
    wire N__9419;
    wire N__9418;
    wire N__9417;
    wire N__9416;
    wire N__9415;
    wire N__9414;
    wire N__9413;
    wire N__9412;
    wire N__9387;
    wire N__9384;
    wire N__9381;
    wire N__9380;
    wire N__9377;
    wire N__9374;
    wire N__9369;
    wire N__9366;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9347;
    wire N__9342;
    wire N__9339;
    wire N__9336;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9328;
    wire N__9325;
    wire N__9322;
    wire N__9319;
    wire N__9312;
    wire N__9309;
    wire N__9308;
    wire N__9305;
    wire N__9304;
    wire N__9303;
    wire N__9302;
    wire N__9301;
    wire N__9298;
    wire N__9295;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9272;
    wire N__9271;
    wire N__9270;
    wire N__9267;
    wire N__9264;
    wire N__9261;
    wire N__9258;
    wire N__9249;
    wire N__9248;
    wire N__9247;
    wire N__9246;
    wire N__9243;
    wire N__9240;
    wire N__9237;
    wire N__9236;
    wire N__9231;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9208;
    wire N__9205;
    wire N__9202;
    wire N__9199;
    wire N__9192;
    wire N__9189;
    wire N__9186;
    wire N__9183;
    wire N__9180;
    wire N__9179;
    wire N__9178;
    wire N__9177;
    wire N__9174;
    wire N__9171;
    wire N__9170;
    wire N__9169;
    wire N__9168;
    wire N__9167;
    wire N__9164;
    wire N__9163;
    wire N__9160;
    wire N__9159;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9137;
    wire N__9136;
    wire N__9135;
    wire N__9132;
    wire N__9127;
    wire N__9122;
    wire N__9119;
    wire N__9114;
    wire N__9111;
    wire N__9108;
    wire N__9107;
    wire N__9106;
    wire N__9105;
    wire N__9100;
    wire N__9099;
    wire N__9090;
    wire N__9087;
    wire N__9084;
    wire N__9079;
    wire N__9076;
    wire N__9073;
    wire N__9072;
    wire N__9071;
    wire N__9070;
    wire N__9067;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9053;
    wire N__9050;
    wire N__9045;
    wire N__9044;
    wire N__9037;
    wire N__9028;
    wire N__9025;
    wire N__9018;
    wire N__9015;
    wire N__9012;
    wire N__9009;
    wire N__9006;
    wire N__9003;
    wire N__9000;
    wire N__8999;
    wire N__8996;
    wire N__8991;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8979;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8967;
    wire N__8964;
    wire N__8961;
    wire N__8958;
    wire N__8955;
    wire N__8952;
    wire N__8949;
    wire N__8946;
    wire N__8943;
    wire N__8940;
    wire N__8937;
    wire N__8934;
    wire N__8931;
    wire N__8928;
    wire N__8925;
    wire N__8922;
    wire N__8919;
    wire N__8916;
    wire N__8913;
    wire N__8912;
    wire N__8911;
    wire N__8910;
    wire N__8909;
    wire N__8908;
    wire N__8905;
    wire N__8900;
    wire N__8897;
    wire N__8892;
    wire N__8883;
    wire N__8880;
    wire N__8877;
    wire N__8876;
    wire N__8875;
    wire N__8874;
    wire N__8873;
    wire N__8870;
    wire N__8863;
    wire N__8860;
    wire N__8853;
    wire N__8850;
    wire N__8847;
    wire N__8846;
    wire N__8845;
    wire N__8844;
    wire N__8841;
    wire N__8834;
    wire N__8829;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8821;
    wire N__8814;
    wire N__8811;
    wire N__8808;
    wire N__8807;
    wire N__8806;
    wire N__8805;
    wire N__8802;
    wire N__8797;
    wire N__8794;
    wire N__8787;
    wire N__8786;
    wire N__8785;
    wire N__8780;
    wire N__8777;
    wire N__8772;
    wire N__8769;
    wire N__8766;
    wire N__8763;
    wire N__8760;
    wire N__8757;
    wire N__8754;
    wire N__8751;
    wire N__8748;
    wire N__8745;
    wire N__8742;
    wire N__8739;
    wire N__8736;
    wire N__8733;
    wire N__8730;
    wire N__8727;
    wire N__8724;
    wire N__8721;
    wire N__8718;
    wire N__8715;
    wire N__8712;
    wire N__8709;
    wire N__8706;
    wire N__8703;
    wire N__8702;
    wire N__8699;
    wire N__8698;
    wire N__8695;
    wire N__8692;
    wire N__8689;
    wire N__8686;
    wire N__8681;
    wire N__8676;
    wire N__8673;
    wire N__8670;
    wire N__8667;
    wire N__8664;
    wire N__8661;
    wire N__8658;
    wire N__8655;
    wire N__8652;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8634;
    wire N__8633;
    wire N__8632;
    wire N__8631;
    wire N__8630;
    wire N__8627;
    wire N__8626;
    wire N__8625;
    wire N__8620;
    wire N__8617;
    wire N__8614;
    wire N__8611;
    wire N__8608;
    wire N__8605;
    wire N__8592;
    wire N__8591;
    wire N__8590;
    wire N__8587;
    wire N__8586;
    wire N__8585;
    wire N__8582;
    wire N__8581;
    wire N__8578;
    wire N__8575;
    wire N__8572;
    wire N__8569;
    wire N__8564;
    wire N__8553;
    wire N__8552;
    wire N__8551;
    wire N__8548;
    wire N__8547;
    wire N__8546;
    wire N__8545;
    wire N__8540;
    wire N__8535;
    wire N__8532;
    wire N__8529;
    wire N__8520;
    wire N__8519;
    wire N__8518;
    wire N__8517;
    wire N__8516;
    wire N__8515;
    wire N__8512;
    wire N__8507;
    wire N__8504;
    wire N__8499;
    wire N__8490;
    wire N__8487;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8469;
    wire N__8466;
    wire N__8465;
    wire N__8464;
    wire N__8461;
    wire N__8458;
    wire N__8455;
    wire N__8450;
    wire N__8447;
    wire N__8442;
    wire N__8439;
    wire N__8438;
    wire N__8435;
    wire N__8432;
    wire N__8429;
    wire N__8426;
    wire N__8421;
    wire N__8418;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8406;
    wire N__8403;
    wire N__8400;
    wire N__8397;
    wire N__8394;
    wire N__8391;
    wire N__8388;
    wire N__8385;
    wire N__8384;
    wire N__8383;
    wire N__8382;
    wire N__8381;
    wire N__8380;
    wire N__8377;
    wire N__8374;
    wire N__8373;
    wire N__8370;
    wire N__8365;
    wire N__8362;
    wire N__8359;
    wire N__8354;
    wire N__8351;
    wire N__8350;
    wire N__8349;
    wire N__8348;
    wire N__8347;
    wire N__8346;
    wire N__8345;
    wire N__8344;
    wire N__8343;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8330;
    wire N__8329;
    wire N__8298;
    wire N__8295;
    wire N__8292;
    wire N__8289;
    wire N__8286;
    wire N__8283;
    wire N__8280;
    wire N__8277;
    wire N__8274;
    wire N__8271;
    wire N__8268;
    wire N__8265;
    wire N__8262;
    wire N__8259;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8247;
    wire N__8246;
    wire N__8243;
    wire N__8240;
    wire N__8237;
    wire N__8234;
    wire N__8229;
    wire N__8226;
    wire N__8223;
    wire N__8222;
    wire N__8221;
    wire N__8218;
    wire N__8213;
    wire N__8208;
    wire N__8207;
    wire N__8206;
    wire N__8205;
    wire N__8202;
    wire N__8199;
    wire N__8196;
    wire N__8193;
    wire N__8186;
    wire N__8181;
    wire N__8180;
    wire N__8179;
    wire N__8178;
    wire N__8175;
    wire N__8168;
    wire N__8163;
    wire N__8162;
    wire N__8161;
    wire N__8158;
    wire N__8153;
    wire N__8148;
    wire N__8145;
    wire N__8144;
    wire N__8141;
    wire N__8138;
    wire N__8133;
    wire N__8130;
    wire N__8129;
    wire N__8126;
    wire N__8123;
    wire N__8120;
    wire N__8117;
    wire N__8112;
    wire N__8109;
    wire N__8106;
    wire N__8105;
    wire N__8102;
    wire N__8099;
    wire N__8094;
    wire N__8091;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8079;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8067;
    wire N__8066;
    wire N__8061;
    wire N__8058;
    wire N__8055;
    wire N__8052;
    wire N__8049;
    wire N__8046;
    wire N__8043;
    wire N__8040;
    wire N__8039;
    wire N__8036;
    wire N__8033;
    wire N__8030;
    wire N__8027;
    wire N__8022;
    wire N__8019;
    wire N__8016;
    wire N__8013;
    wire N__8010;
    wire N__8007;
    wire N__8004;
    wire N__8001;
    wire N__7998;
    wire N__7995;
    wire N__7992;
    wire N__7989;
    wire N__7986;
    wire N__7983;
    wire N__7980;
    wire N__7977;
    wire N__7974;
    wire N__7971;
    wire N__7968;
    wire N__7965;
    wire N__7964;
    wire N__7963;
    wire N__7962;
    wire N__7959;
    wire N__7956;
    wire N__7953;
    wire N__7952;
    wire N__7949;
    wire N__7944;
    wire N__7941;
    wire N__7938;
    wire N__7937;
    wire N__7936;
    wire N__7933;
    wire N__7926;
    wire N__7923;
    wire N__7920;
    wire N__7917;
    wire N__7912;
    wire N__7909;
    wire N__7906;
    wire N__7903;
    wire N__7900;
    wire N__7897;
    wire N__7894;
    wire N__7891;
    wire N__7886;
    wire N__7881;
    wire N__7878;
    wire N__7875;
    wire N__7874;
    wire N__7871;
    wire N__7870;
    wire N__7867;
    wire N__7864;
    wire N__7861;
    wire N__7858;
    wire N__7857;
    wire N__7850;
    wire N__7847;
    wire N__7842;
    wire N__7839;
    wire N__7836;
    wire N__7835;
    wire N__7832;
    wire N__7829;
    wire N__7828;
    wire N__7823;
    wire N__7820;
    wire N__7815;
    wire N__7812;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7804;
    wire N__7803;
    wire N__7802;
    wire N__7797;
    wire N__7794;
    wire N__7791;
    wire N__7788;
    wire N__7787;
    wire N__7784;
    wire N__7781;
    wire N__7778;
    wire N__7775;
    wire N__7772;
    wire N__7767;
    wire N__7764;
    wire N__7759;
    wire N__7756;
    wire N__7751;
    wire N__7746;
    wire N__7743;
    wire N__7740;
    wire N__7737;
    wire N__7736;
    wire N__7733;
    wire N__7730;
    wire N__7725;
    wire N__7722;
    wire N__7719;
    wire N__7718;
    wire N__7715;
    wire N__7712;
    wire N__7711;
    wire N__7708;
    wire N__7705;
    wire N__7702;
    wire N__7701;
    wire N__7700;
    wire N__7699;
    wire N__7696;
    wire N__7691;
    wire N__7688;
    wire N__7685;
    wire N__7682;
    wire N__7679;
    wire N__7676;
    wire N__7673;
    wire N__7668;
    wire N__7659;
    wire N__7656;
    wire N__7655;
    wire N__7650;
    wire N__7647;
    wire N__7646;
    wire N__7645;
    wire N__7644;
    wire N__7643;
    wire N__7640;
    wire N__7639;
    wire N__7638;
    wire N__7629;
    wire N__7626;
    wire N__7625;
    wire N__7624;
    wire N__7623;
    wire N__7620;
    wire N__7619;
    wire N__7618;
    wire N__7615;
    wire N__7612;
    wire N__7609;
    wire N__7594;
    wire N__7591;
    wire N__7588;
    wire N__7585;
    wire N__7578;
    wire N__7577;
    wire N__7574;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire N__7562;
    wire N__7559;
    wire N__7558;
    wire N__7555;
    wire N__7552;
    wire N__7549;
    wire N__7546;
    wire N__7543;
    wire N__7540;
    wire N__7535;
    wire N__7532;
    wire N__7527;
    wire N__7524;
    wire N__7523;
    wire N__7518;
    wire N__7515;
    wire N__7512;
    wire N__7509;
    wire N__7506;
    wire N__7505;
    wire N__7502;
    wire N__7499;
    wire N__7494;
    wire N__7493;
    wire N__7492;
    wire N__7491;
    wire N__7482;
    wire N__7479;
    wire N__7476;
    wire N__7475;
    wire N__7472;
    wire N__7471;
    wire N__7470;
    wire N__7469;
    wire N__7468;
    wire N__7465;
    wire N__7464;
    wire N__7461;
    wire N__7458;
    wire N__7455;
    wire N__7452;
    wire N__7451;
    wire N__7450;
    wire N__7447;
    wire N__7444;
    wire N__7443;
    wire N__7440;
    wire N__7435;
    wire N__7432;
    wire N__7429;
    wire N__7424;
    wire N__7421;
    wire N__7418;
    wire N__7413;
    wire N__7398;
    wire N__7395;
    wire N__7394;
    wire N__7393;
    wire N__7392;
    wire N__7391;
    wire N__7388;
    wire N__7383;
    wire N__7378;
    wire N__7371;
    wire N__7370;
    wire N__7369;
    wire N__7368;
    wire N__7367;
    wire N__7366;
    wire N__7365;
    wire N__7364;
    wire N__7363;
    wire N__7362;
    wire N__7357;
    wire N__7350;
    wire N__7347;
    wire N__7346;
    wire N__7343;
    wire N__7340;
    wire N__7337;
    wire N__7334;
    wire N__7333;
    wire N__7332;
    wire N__7331;
    wire N__7330;
    wire N__7329;
    wire N__7328;
    wire N__7327;
    wire N__7326;
    wire N__7325;
    wire N__7320;
    wire N__7317;
    wire N__7312;
    wire N__7305;
    wire N__7294;
    wire N__7291;
    wire N__7286;
    wire N__7285;
    wire N__7284;
    wire N__7281;
    wire N__7280;
    wire N__7275;
    wire N__7272;
    wire N__7263;
    wire N__7258;
    wire N__7255;
    wire N__7252;
    wire N__7249;
    wire N__7246;
    wire N__7243;
    wire N__7236;
    wire N__7229;
    wire N__7226;
    wire N__7223;
    wire N__7220;
    wire N__7217;
    wire N__7212;
    wire N__7209;
    wire N__7206;
    wire N__7203;
    wire N__7202;
    wire N__7201;
    wire N__7198;
    wire N__7195;
    wire N__7192;
    wire N__7189;
    wire N__7188;
    wire N__7183;
    wire N__7182;
    wire N__7179;
    wire N__7176;
    wire N__7173;
    wire N__7170;
    wire N__7161;
    wire N__7160;
    wire N__7157;
    wire N__7154;
    wire N__7149;
    wire N__7146;
    wire N__7143;
    wire N__7140;
    wire N__7139;
    wire N__7136;
    wire N__7135;
    wire N__7134;
    wire N__7131;
    wire N__7128;
    wire N__7125;
    wire N__7122;
    wire N__7121;
    wire N__7118;
    wire N__7113;
    wire N__7110;
    wire N__7107;
    wire N__7104;
    wire N__7101;
    wire N__7094;
    wire N__7091;
    wire N__7088;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7074;
    wire N__7071;
    wire N__7068;
    wire N__7067;
    wire N__7064;
    wire N__7061;
    wire N__7060;
    wire N__7059;
    wire N__7056;
    wire N__7053;
    wire N__7048;
    wire N__7041;
    wire N__7040;
    wire N__7039;
    wire N__7038;
    wire N__7037;
    wire N__7036;
    wire N__7035;
    wire N__7032;
    wire N__7027;
    wire N__7024;
    wire N__7017;
    wire N__7008;
    wire N__7007;
    wire N__7006;
    wire N__7005;
    wire N__7002;
    wire N__6999;
    wire N__6994;
    wire N__6987;
    wire N__6986;
    wire N__6985;
    wire N__6984;
    wire N__6983;
    wire N__6980;
    wire N__6977;
    wire N__6974;
    wire N__6971;
    wire N__6968;
    wire N__6957;
    wire N__6956;
    wire N__6953;
    wire N__6952;
    wire N__6949;
    wire N__6944;
    wire N__6939;
    wire N__6936;
    wire N__6933;
    wire N__6932;
    wire N__6931;
    wire N__6928;
    wire N__6925;
    wire N__6922;
    wire N__6921;
    wire N__6920;
    wire N__6915;
    wire N__6912;
    wire N__6911;
    wire N__6906;
    wire N__6901;
    wire N__6900;
    wire N__6897;
    wire N__6894;
    wire N__6893;
    wire N__6890;
    wire N__6887;
    wire N__6884;
    wire N__6881;
    wire N__6878;
    wire N__6867;
    wire N__6864;
    wire N__6861;
    wire N__6858;
    wire N__6855;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6843;
    wire N__6842;
    wire N__6839;
    wire N__6836;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6822;
    wire N__6819;
    wire N__6816;
    wire N__6813;
    wire N__6810;
    wire N__6809;
    wire N__6808;
    wire N__6805;
    wire N__6802;
    wire N__6799;
    wire N__6792;
    wire N__6789;
    wire N__6786;
    wire N__6783;
    wire N__6782;
    wire N__6779;
    wire N__6776;
    wire N__6775;
    wire N__6774;
    wire N__6771;
    wire N__6768;
    wire N__6765;
    wire N__6764;
    wire N__6763;
    wire N__6760;
    wire N__6753;
    wire N__6750;
    wire N__6747;
    wire N__6738;
    wire N__6737;
    wire N__6736;
    wire N__6735;
    wire N__6732;
    wire N__6727;
    wire N__6724;
    wire N__6723;
    wire N__6722;
    wire N__6717;
    wire N__6714;
    wire N__6709;
    wire N__6702;
    wire N__6699;
    wire N__6698;
    wire N__6697;
    wire N__6696;
    wire N__6695;
    wire N__6694;
    wire N__6689;
    wire N__6686;
    wire N__6683;
    wire N__6680;
    wire N__6677;
    wire N__6674;
    wire N__6671;
    wire N__6666;
    wire N__6663;
    wire N__6662;
    wire N__6661;
    wire N__6654;
    wire N__6651;
    wire N__6646;
    wire N__6639;
    wire N__6636;
    wire N__6633;
    wire N__6630;
    wire N__6627;
    wire N__6624;
    wire N__6621;
    wire N__6618;
    wire N__6615;
    wire N__6614;
    wire N__6613;
    wire N__6612;
    wire N__6609;
    wire N__6608;
    wire N__6607;
    wire N__6606;
    wire N__6603;
    wire N__6600;
    wire N__6597;
    wire N__6594;
    wire N__6591;
    wire N__6590;
    wire N__6587;
    wire N__6586;
    wire N__6583;
    wire N__6578;
    wire N__6573;
    wire N__6570;
    wire N__6567;
    wire N__6564;
    wire N__6561;
    wire N__6558;
    wire N__6551;
    wire N__6548;
    wire N__6541;
    wire N__6538;
    wire N__6533;
    wire N__6528;
    wire N__6525;
    wire N__6522;
    wire N__6519;
    wire N__6516;
    wire N__6515;
    wire N__6512;
    wire N__6509;
    wire N__6504;
    wire N__6501;
    wire N__6498;
    wire N__6495;
    wire N__6494;
    wire N__6491;
    wire N__6488;
    wire N__6485;
    wire N__6480;
    wire N__6477;
    wire N__6476;
    wire N__6471;
    wire N__6468;
    wire N__6465;
    wire N__6462;
    wire N__6459;
    wire N__6456;
    wire N__6455;
    wire N__6452;
    wire N__6449;
    wire N__6448;
    wire N__6443;
    wire N__6440;
    wire N__6437;
    wire N__6434;
    wire N__6431;
    wire N__6428;
    wire N__6425;
    wire N__6422;
    wire N__6417;
    wire N__6414;
    wire N__6411;
    wire N__6410;
    wire N__6407;
    wire N__6404;
    wire N__6401;
    wire N__6398;
    wire N__6393;
    wire N__6390;
    wire N__6389;
    wire N__6386;
    wire N__6383;
    wire N__6378;
    wire N__6377;
    wire N__6376;
    wire N__6373;
    wire N__6370;
    wire N__6367;
    wire N__6364;
    wire N__6363;
    wire N__6362;
    wire N__6359;
    wire N__6354;
    wire N__6351;
    wire N__6348;
    wire N__6339;
    wire N__6336;
    wire N__6333;
    wire N__6330;
    wire N__6327;
    wire N__6324;
    wire N__6321;
    wire N__6320;
    wire N__6319;
    wire N__6318;
    wire N__6313;
    wire N__6310;
    wire N__6307;
    wire N__6306;
    wire N__6303;
    wire N__6300;
    wire N__6297;
    wire N__6294;
    wire N__6291;
    wire N__6284;
    wire N__6281;
    wire N__6278;
    wire N__6275;
    wire N__6272;
    wire N__6267;
    wire N__6264;
    wire N__6263;
    wire N__6262;
    wire N__6261;
    wire N__6260;
    wire N__6257;
    wire N__6256;
    wire N__6253;
    wire N__6248;
    wire N__6241;
    wire N__6234;
    wire N__6233;
    wire N__6230;
    wire N__6227;
    wire N__6222;
    wire N__6221;
    wire N__6218;
    wire N__6215;
    wire N__6210;
    wire N__6209;
    wire N__6206;
    wire N__6203;
    wire N__6200;
    wire N__6197;
    wire N__6192;
    wire N__6191;
    wire N__6188;
    wire N__6185;
    wire N__6182;
    wire N__6179;
    wire N__6176;
    wire N__6173;
    wire N__6168;
    wire N__6165;
    wire N__6164;
    wire N__6161;
    wire N__6158;
    wire N__6153;
    wire N__6150;
    wire N__6149;
    wire N__6146;
    wire N__6143;
    wire N__6138;
    wire N__6137;
    wire N__6134;
    wire N__6131;
    wire N__6126;
    wire N__6123;
    wire N__6120;
    wire N__6117;
    wire N__6116;
    wire N__6113;
    wire N__6112;
    wire N__6111;
    wire N__6108;
    wire N__6105;
    wire N__6102;
    wire N__6099;
    wire N__6092;
    wire N__6089;
    wire N__6088;
    wire N__6085;
    wire N__6082;
    wire N__6079;
    wire N__6072;
    wire N__6069;
    wire N__6066;
    wire N__6063;
    wire N__6062;
    wire N__6059;
    wire N__6056;
    wire N__6051;
    wire N__6048;
    wire N__6045;
    wire N__6042;
    wire N__6039;
    wire N__6038;
    wire N__6033;
    wire N__6030;
    wire N__6029;
    wire N__6024;
    wire N__6021;
    wire N__6018;
    wire N__6015;
    wire N__6012;
    wire N__6011;
    wire N__6008;
    wire N__6007;
    wire N__6006;
    wire N__6003;
    wire N__6002;
    wire N__6001;
    wire N__5996;
    wire N__5993;
    wire N__5990;
    wire N__5985;
    wire N__5976;
    wire N__5975;
    wire N__5974;
    wire N__5971;
    wire N__5970;
    wire N__5969;
    wire N__5966;
    wire N__5963;
    wire N__5960;
    wire N__5955;
    wire N__5946;
    wire N__5943;
    wire N__5942;
    wire N__5939;
    wire N__5936;
    wire N__5933;
    wire N__5930;
    wire N__5925;
    wire N__5922;
    wire N__5919;
    wire N__5918;
    wire N__5915;
    wire N__5912;
    wire N__5907;
    wire N__5904;
    wire N__5901;
    wire N__5898;
    wire N__5895;
    wire N__5892;
    wire N__5889;
    wire N__5888;
    wire N__5883;
    wire N__5880;
    wire N__5879;
    wire N__5874;
    wire N__5871;
    wire N__5870;
    wire N__5869;
    wire N__5866;
    wire N__5861;
    wire N__5858;
    wire N__5855;
    wire N__5852;
    wire N__5849;
    wire N__5846;
    wire N__5841;
    wire N__5838;
    wire N__5835;
    wire N__5832;
    wire N__5831;
    wire N__5826;
    wire N__5823;
    wire N__5822;
    wire N__5819;
    wire N__5816;
    wire N__5813;
    wire N__5810;
    wire N__5807;
    wire N__5804;
    wire N__5799;
    wire N__5796;
    wire N__5793;
    wire N__5790;
    wire N__5789;
    wire N__5788;
    wire N__5787;
    wire N__5782;
    wire N__5777;
    wire N__5772;
    wire N__5771;
    wire N__5768;
    wire N__5767;
    wire N__5764;
    wire N__5759;
    wire N__5754;
    wire N__5751;
    wire N__5748;
    wire N__5745;
    wire N__5742;
    wire N__5741;
    wire N__5736;
    wire N__5733;
    wire N__5732;
    wire N__5729;
    wire N__5724;
    wire N__5721;
    wire N__5718;
    wire N__5715;
    wire N__5714;
    wire N__5713;
    wire N__5710;
    wire N__5707;
    wire N__5706;
    wire N__5703;
    wire N__5696;
    wire N__5691;
    wire N__5688;
    wire N__5685;
    wire N__5684;
    wire N__5683;
    wire N__5680;
    wire N__5677;
    wire N__5674;
    wire N__5669;
    wire N__5666;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5652;
    wire N__5651;
    wire N__5648;
    wire N__5645;
    wire N__5640;
    wire N__5637;
    wire N__5636;
    wire N__5633;
    wire N__5630;
    wire N__5625;
    wire N__5624;
    wire N__5621;
    wire N__5618;
    wire N__5615;
    wire N__5614;
    wire N__5611;
    wire N__5608;
    wire N__5605;
    wire N__5602;
    wire N__5597;
    wire N__5594;
    wire N__5591;
    wire N__5588;
    wire N__5585;
    wire N__5580;
    wire N__5577;
    wire N__5574;
    wire N__5573;
    wire N__5572;
    wire N__5571;
    wire N__5562;
    wire N__5559;
    wire N__5558;
    wire N__5557;
    wire N__5556;
    wire N__5553;
    wire N__5548;
    wire N__5545;
    wire N__5538;
    wire N__5537;
    wire N__5536;
    wire N__5529;
    wire N__5526;
    wire N__5525;
    wire N__5522;
    wire N__5519;
    wire N__5516;
    wire N__5513;
    wire N__5508;
    wire N__5505;
    wire N__5502;
    wire N__5499;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5487;
    wire N__5484;
    wire N__5481;
    wire N__5478;
    wire N__5475;
    wire N__5472;
    wire N__5469;
    wire N__5466;
    wire N__5463;
    wire N__5460;
    wire N__5457;
    wire N__5454;
    wire N__5451;
    wire N__5448;
    wire N__5447;
    wire N__5446;
    wire N__5443;
    wire N__5440;
    wire N__5437;
    wire N__5432;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5409;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5397;
    wire N__5396;
    wire N__5395;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5351;
    wire N__5346;
    wire N__5345;
    wire N__5342;
    wire N__5339;
    wire N__5334;
    wire N__5331;
    wire N__5328;
    wire N__5325;
    wire N__5324;
    wire N__5323;
    wire N__5320;
    wire N__5317;
    wire N__5314;
    wire N__5307;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5289;
    wire N__5286;
    wire N__5283;
    wire N__5280;
    wire N__5277;
    wire N__5274;
    wire N__5271;
    wire N__5268;
    wire N__5265;
    wire N__5262;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5250;
    wire N__5249;
    wire N__5248;
    wire N__5247;
    wire N__5244;
    wire N__5241;
    wire N__5236;
    wire N__5233;
    wire N__5232;
    wire N__5231;
    wire N__5230;
    wire N__5229;
    wire N__5228;
    wire N__5227;
    wire N__5224;
    wire N__5221;
    wire N__5218;
    wire N__5211;
    wire N__5208;
    wire N__5205;
    wire N__5204;
    wire N__5201;
    wire N__5196;
    wire N__5191;
    wire N__5182;
    wire N__5175;
    wire N__5172;
    wire N__5169;
    wire N__5168;
    wire N__5167;
    wire N__5166;
    wire N__5165;
    wire N__5162;
    wire N__5155;
    wire N__5154;
    wire N__5153;
    wire N__5152;
    wire N__5151;
    wire N__5148;
    wire N__5143;
    wire N__5140;
    wire N__5137;
    wire N__5132;
    wire N__5125;
    wire N__5120;
    wire N__5117;
    wire N__5114;
    wire N__5111;
    wire N__5108;
    wire N__5103;
    wire N__5100;
    wire N__5097;
    wire N__5094;
    wire N__5091;
    wire N__5088;
    wire N__5085;
    wire N__5082;
    wire N__5079;
    wire N__5076;
    wire N__5073;
    wire N__5070;
    wire N__5067;
    wire N__5064;
    wire N__5061;
    wire N__5058;
    wire N__5055;
    wire N__5054;
    wire N__5051;
    wire N__5048;
    wire N__5043;
    wire N__5042;
    wire N__5039;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5027;
    wire N__5024;
    wire N__5019;
    wire N__5018;
    wire N__5015;
    wire N__5012;
    wire N__5011;
    wire N__5006;
    wire N__5003;
    wire N__4998;
    wire N__4995;
    wire N__4992;
    wire N__4989;
    wire N__4986;
    wire N__4983;
    wire N__4980;
    wire N__4977;
    wire N__4974;
    wire N__4973;
    wire N__4972;
    wire N__4969;
    wire N__4966;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4934;
    wire N__4931;
    wire N__4928;
    wire N__4923;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4905;
    wire N__4902;
    wire N__4899;
    wire N__4896;
    wire N__4895;
    wire N__4892;
    wire N__4889;
    wire N__4884;
    wire N__4881;
    wire N__4878;
    wire N__4877;
    wire N__4874;
    wire N__4871;
    wire N__4866;
    wire N__4863;
    wire N__4860;
    wire N__4857;
    wire N__4854;
    wire N__4853;
    wire N__4850;
    wire N__4845;
    wire N__4842;
    wire N__4841;
    wire N__4840;
    wire N__4837;
    wire N__4836;
    wire N__4835;
    wire N__4834;
    wire N__4831;
    wire N__4830;
    wire N__4827;
    wire N__4818;
    wire N__4817;
    wire N__4816;
    wire N__4813;
    wire N__4812;
    wire N__4811;
    wire N__4810;
    wire N__4809;
    wire N__4806;
    wire N__4801;
    wire N__4796;
    wire N__4793;
    wire N__4786;
    wire N__4783;
    wire N__4780;
    wire N__4775;
    wire N__4768;
    wire N__4765;
    wire N__4762;
    wire N__4759;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4743;
    wire N__4742;
    wire N__4741;
    wire N__4740;
    wire N__4739;
    wire N__4738;
    wire N__4737;
    wire N__4736;
    wire N__4733;
    wire N__4732;
    wire N__4729;
    wire N__4726;
    wire N__4725;
    wire N__4722;
    wire N__4721;
    wire N__4718;
    wire N__4711;
    wire N__4704;
    wire N__4699;
    wire N__4696;
    wire N__4693;
    wire N__4692;
    wire N__4687;
    wire N__4684;
    wire N__4677;
    wire N__4676;
    wire N__4673;
    wire N__4672;
    wire N__4669;
    wire N__4664;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4644;
    wire N__4641;
    wire N__4638;
    wire N__4635;
    wire N__4632;
    wire N__4629;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4617;
    wire N__4616;
    wire N__4613;
    wire N__4608;
    wire N__4605;
    wire N__4602;
    wire N__4599;
    wire N__4596;
    wire N__4593;
    wire N__4590;
    wire N__4587;
    wire N__4584;
    wire N__4581;
    wire N__4578;
    wire N__4575;
    wire N__4574;
    wire N__4573;
    wire N__4572;
    wire N__4563;
    wire N__4560;
    wire N__4557;
    wire N__4554;
    wire N__4551;
    wire N__4548;
    wire N__4545;
    wire N__4542;
    wire N__4539;
    wire N__4536;
    wire N__4533;
    wire N__4532;
    wire N__4531;
    wire N__4530;
    wire N__4521;
    wire N__4518;
    wire N__4515;
    wire N__4512;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4504;
    wire N__4501;
    wire N__4498;
    wire N__4495;
    wire N__4494;
    wire N__4493;
    wire N__4492;
    wire N__4489;
    wire N__4484;
    wire N__4477;
    wire N__4470;
    wire N__4467;
    wire N__4466;
    wire N__4465;
    wire N__4464;
    wire N__4463;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4447;
    wire N__4444;
    wire N__4441;
    wire N__4438;
    wire N__4431;
    wire N__4428;
    wire N__4425;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4407;
    wire N__4404;
    wire N__4401;
    wire N__4398;
    wire N__4395;
    wire N__4392;
    wire N__4389;
    wire N__4386;
    wire N__4383;
    wire N__4380;
    wire N__4377;
    wire N__4374;
    wire N__4371;
    wire N__4368;
    wire N__4365;
    wire N__4362;
    wire N__4361;
    wire N__4360;
    wire N__4359;
    wire N__4354;
    wire N__4351;
    wire N__4348;
    wire N__4345;
    wire N__4342;
    wire N__4339;
    wire N__4332;
    wire N__4331;
    wire N__4328;
    wire N__4325;
    wire N__4320;
    wire N__4317;
    wire N__4314;
    wire N__4311;
    wire N__4310;
    wire N__4305;
    wire N__4302;
    wire N__4299;
    wire N__4298;
    wire N__4295;
    wire N__4292;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4280;
    wire N__4277;
    wire N__4274;
    wire N__4269;
    wire N__4266;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4254;
    wire N__4251;
    wire N__4248;
    wire N__4245;
    wire N__4242;
    wire N__4239;
    wire N__4236;
    wire N__4233;
    wire N__4230;
    wire N__4227;
    wire N__4224;
    wire N__4221;
    wire N__4218;
    wire N__4215;
    wire N__4214;
    wire N__4209;
    wire N__4206;
    wire N__4203;
    wire N__4200;
    wire N__4197;
    wire N__4196;
    wire N__4191;
    wire N__4188;
    wire N__4185;
    wire N__4182;
    wire N__4179;
    wire N__4178;
    wire N__4175;
    wire N__4170;
    wire N__4167;
    wire N__4164;
    wire N__4161;
    wire N__4158;
    wire N__4155;
    wire N__4152;
    wire N__4149;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4137;
    wire N__4134;
    wire N__4131;
    wire N__4128;
    wire N__4125;
    wire N__4122;
    wire N__4119;
    wire N__4116;
    wire N__4113;
    wire N__4110;
    wire N__4109;
    wire N__4108;
    wire N__4107;
    wire N__4106;
    wire N__4105;
    wire N__4104;
    wire N__4103;
    wire N__4102;
    wire N__4101;
    wire N__4100;
    wire N__4077;
    wire CLK80_OUT;
    wire PIO_S0_c;
    wire GNDG0;
    wire PIO_P0_c;
    wire VCCG0;
    wire A_c_25;
    wire A_c_27;
    wire A_c_26;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_8_cascade_ ;
    wire A_c_24;
    wire \U409_AUTOCONFIG.N_270 ;
    wire \U409_AUTOCONFIG.N_271 ;
    wire \U409_AUTOCONFIG.N_433_cascade_ ;
    wire \U409_AUTOCONFIG.N_433 ;
    wire \U409_AUTOCONFIG.N_373 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_2_3_0_cascade_ ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_0_0 ;
    wire \U409_AUTOCONFIG.N_269 ;
    wire \U409_AUTOCONFIG.N_370 ;
    wire \U409_AUTOCONFIG.N_195_cascade_ ;
    wire \U409_AUTOCONFIG.N_383 ;
    wire \U409_AUTOCONFIG.N_274 ;
    wire \U409_AUTOCONFIG.N_383_cascade_ ;
    wire TT_c_0;
    wire TT_c_1;
    wire \U409_ADDRESS_DECODE.N_345 ;
    wire \U409_ADDRESS_DECODE.N_344 ;
    wire \U409_AUTOCONFIG.N_288_cascade_ ;
    wire \U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_0_0_a2Z0Z_1 ;
    wire \U409_AUTOCONFIG.N_405_cascade_ ;
    wire \U409_AUTOCONFIG.N_414 ;
    wire \U409_AUTOCONFIG.N_285 ;
    wire \U409_AUTOCONFIG.N_9 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_0_1 ;
    wire \U409_AUTOCONFIG.N_405 ;
    wire \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net ;
    wire \U409_AUTOCONFIG.LIDE_OUTc_0_1 ;
    wire \U409_AUTOCONFIG.LIDE_OUTc_0_0 ;
    wire \U409_AUTOCONFIG.N_286 ;
    wire \U409_AUTOCONFIG.AC_START_RNI3D7VZ0Z2 ;
    wire \INVU409_AUTOCONFIG.LIDE_OUT_0C_net ;
    wire \U409_AUTOCONFIG.N_287 ;
    wire A_c_6;
    wire A_c_7;
    wire \U409_AUTOCONFIG.N_273 ;
    wire \U409_AUTOCONFIG.N_400 ;
    wire A_c_2;
    wire A_c_4;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_10 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_11 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_9_cascade_ ;
    wire N_374;
    wire N_401_cascade_;
    wire N_436;
    wire N_265_i;
    wire U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_o2_4;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_0 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ1Z_0 ;
    wire N_124;
    wire \U409_AUTOCONFIG.un1_STATE_1_0_a2_0Z0Z_2 ;
    wire CPUCONFn_c;
    wire \U409_AUTOCONFIG.AC_STARTZ0 ;
    wire \INVU409_AUTOCONFIG.STATE_0C_net ;
    wire N_354_cascade_;
    wire D_1_i;
    wire AUTOBOOT_c;
    wire \U409_AUTOCONFIG.N_360 ;
    wire A_c_5;
    wire A_c_3;
    wire \U409_AUTOCONFIG.N_276 ;
    wire \U409_ADDRESS_DECODE.PORTSIZE_iZ0Z_1_cascade_ ;
    wire N_139;
    wire \U409_ADDRESS_DECODE.N_343 ;
    wire TM_c_1;
    wire TM_c_0;
    wire U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_o2_5;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ;
    wire N_126;
    wire \INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net ;
    wire N_96;
    wire A_c_29;
    wire BRIDGE_BASE_1;
    wire A_c_28;
    wire BRIDGE_BASE_0;
    wire \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0Z0Z_0 ;
    wire A_c_31;
    wire BRIDGE_BASE_3;
    wire BRIDGE_BASE_2;
    wire A_c_30;
    wire \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0Z0Z_1 ;
    wire \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa ;
    wire \U409_AUTOCONFIG.STATEZ0Z_0 ;
    wire \INVU409_AUTOCONFIG.AC_TACKC_net ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_a2_3_cascade_ ;
    wire \U409_TRANSFER_ACK.N_268_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ;
    wire N_130;
    wire ATA_BASE_4;
    wire ATA_BASE_5;
    wire D_in_4;
    wire D_in_5;
    wire D_in_6;
    wire \INVU409_AUTOCONFIG.ATA_BASE_ness_4C_net ;
    wire ATA_BASE_6;
    wire ATA_BASE_1;
    wire ATA_BASE_0;
    wire \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_7Z0Z_0_cascade_ ;
    wire \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_7_cascade_ ;
    wire \U409_ADDRESS_DECODE.ATA_EN_2_0_o2_3_cascade_ ;
    wire A_c_18;
    wire ATA_BASE_2;
    wire \U409_ADDRESS_DECODE.N_183_i ;
    wire \U409_ADDRESS_DECODE.ATA_EN_2_0_o2_2 ;
    wire \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_2 ;
    wire \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_0 ;
    wire \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_7 ;
    wire \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_o2dupZ0 ;
    wire \U409_ADDRESS_DECODE.un1_ATA_ENn_i_0Z0Z_3_cascade_ ;
    wire \U409_ADDRESS_DECODE.ATA_ENZ0 ;
    wire N_107;
    wire A_c_16;
    wire \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_2 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ;
    wire \U409_AUTOCONFIG.BRIDGE_CONFZ0 ;
    wire N_128;
    wire TSn_c;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ;
    wire \U409_TRANSFER_ACK.N_268 ;
    wire \U409_TRANSFER_ACK.N_237 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ;
    wire RnW_c;
    wire N_356;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ;
    wire A_c_20;
    wire \U409_TRANSFER_ACK.N_346_cascade_ ;
    wire N_434;
    wire N_190_cascade_;
    wire TACKn_in;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ;
    wire A_c_21;
    wire N_351;
    wire N_436_i;
    wire A_c_17;
    wire N_431;
    wire A_c_22;
    wire N_401;
    wire N_431_cascade_;
    wire N_422;
    wire A_c_19;
    wire ATA_BASE_7;
    wire A_c_23;
    wire \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_5 ;
    wire N_361;
    wire D_in_7;
    wire ATA_BASE_3;
    wire \INVU409_AUTOCONFIG.ATA_BASE_ness_3C_net ;
    wire \U409_AUTOCONFIG.un1_STATE_1_0_0 ;
    wire \U409_AUTOCONFIG.N_172 ;
    wire \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ;
    wire \U409_AUTOCONFIG.LIDE_CONFZ0 ;
    wire \U409_AUTOCONFIG.un1_STATE_1_0_a2_0 ;
    wire A_c_1;
    wire CONFIGENn_c;
    wire \INVU409_AUTOCONFIG.CONFIGENnC_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ;
    wire AC_TACK;
    wire \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_ ;
    wire \U409_TRANSFER_ACK.CIA_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net ;
    wire \U409_TRANSFER_ACK.N_159 ;
    wire \U409_TRANSFER_ACK.N_380 ;
    wire \U409_TRANSFER_ACK.N_380_cascade_ ;
    wire N_190;
    wire N_297;
    wire N_94_i;
    wire A_c_13;
    wire U409_ADDRESS_DECODE_un1_CIACS1n_i;
    wire \U409_TRANSFER_ACK.CIA_STATE_d_2_cascade_ ;
    wire \U409_TRANSFER_ACK.N_289 ;
    wire \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ;
    wire TACK_OUTn;
    wire \INVU409_TRANSFER_ACK.TACK_OUTnC_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER6 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.N_379 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0 ;
    wire \U409_TRANSFER_ACK.N_307 ;
    wire \U409_TRANSFER_ACK.N_381 ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0 ;
    wire \U409_TRANSFER_ACK.ROMENn_e_1 ;
    wire ROMENn_c;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ;
    wire TACK_EN;
    wire N_357;
    wire N_339;
    wire TCIn_1_i;
    wire CLK40_IN_c_g;
    wire GB_BUFFER_CLK40_IN_c_g_THRU_CO;
    wire CIA_ENABLE;
    wire CIA_ENABLE_cascade_;
    wire A_c_12;
    wire U409_ADDRESS_DECODE_un1_CIACS0n_i;
    wire \U409_TICK.TICK603_10_cascade_ ;
    wire \U409_TRANSFER_ACK.m12_i_a2_1_0_cascade_ ;
    wire \U409_TRANSFER_ACK.m12_i_0_cascade_ ;
    wire \U409_TRANSFER_ACK.N_293 ;
    wire \U409_TRANSFER_ACK.N_191 ;
    wire \U409_TRANSFER_ACK.N_191_cascade_ ;
    wire \U409_TRANSFER_ACK.N_223 ;
    wire \U409_TRANSFER_ACK.i5_mux_cascade_ ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_0C_net ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ;
    wire \U409_TRANSFER_ACK.N_290 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_0 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ;
    wire RESETn_c_i_g;
    wire OVL_c;
    wire N_429;
    wire N_348;
    wire N_156_i;
    wire N_264_i;
    wire RESETn_c;
    wire RESETn_c_i;
    wire \U409_TICK.COUNTER60Z0Z_1 ;
    wire bfn_13_6_0_;
    wire \U409_TICK.COUNTER60Z0Z_2 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_1 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_2 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_3 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_4 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_6 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_5 ;
    wire \U409_TICK.COUNTER60Z0Z_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_6 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_8 ;
    wire bfn_13_7_0_;
    wire \U409_TICK.COUNTER60Z0Z_10 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_9 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_10 ;
    wire \U409_TICK.COUNTER60Z0Z_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_11 ;
    wire \U409_TICK.COUNTER60Z0Z_13 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_13 ;
    wire \U409_TICK.COUNTER60Z0Z_15 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_15 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_15 ;
    wire \U409_TICK.COUNTER60Z0Z_16 ;
    wire \U409_TICK.COUNTER60Z0Z_11 ;
    wire \U409_TICK.COUNTER60Z0Z_3 ;
    wire \U409_TICK.TICK603_11 ;
    wire \U409_TICK.TICK603_14_cascade_ ;
    wire TICK60_c;
    wire \U409_CIA.CLK_CIA6_0_a2_0_cascade_ ;
    wire \U409_CIA.CLK_CIA6_cascade_ ;
    wire CLK_CIA_c;
    wire \U409_CIA.un1_CIA_CLK_COUNT_3_0_a2_0_cascade_ ;
    wire \U409_CIA.VMA_3_0_a2_2 ;
    wire \U409_CIA.VMA_RNOZ0Z_1_cascade_ ;
    wire \U409_CIA.VMAZ0 ;
    wire bfn_14_5_0_;
    wire \U409_TICK.un2_COUNTER50_1_cry_1 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_3 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_4 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_6 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_8 ;
    wire bfn_14_6_0_;
    wire \U409_TICK.un2_COUNTER50_1_cry_9 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_10 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_11 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_13 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_15 ;
    wire \U409_TICK.COUNTER60Z0Z_5 ;
    wire \U409_TICK.TICK603_8 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_9 ;
    wire \U409_TICK.COUNTER60Z0Z_0 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_4 ;
    wire \U409_TICK.COUNTER60Z0Z_4 ;
    wire \U409_TICK.COUNTER60Z0Z_9 ;
    wire \U409_TICK.COUNTER60Z0Z_6 ;
    wire \U409_TICK.TICK603_9_cascade_ ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_14 ;
    wire \U409_TICK.COUNTER60Z0Z_14 ;
    wire \U409_TICK.TICK603_14 ;
    wire \U409_TICK.TICK603_9 ;
    wire \U409_TICK.TICK603_10 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_8 ;
    wire \U409_TICK.COUNTER60Z0Z_8 ;
    wire bfn_14_9_0_;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_1 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_5 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_6 ;
    wire \U409_CIA.N_427 ;
    wire \U409_CIA.N_427_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNT11 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_6 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_7 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_3 ;
    wire \U409_CIA.un1_CIA_CLK_COUNT_2_0_a2_2_cascade_ ;
    wire \U409_CIA.N_420 ;
    wire \U409_CIA.CLK_CIA_RNOZ0Z_1 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_0 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_1 ;
    wire CLK28_IN_c_g;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_5 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_4 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_2 ;
    wire \U409_CIA.CIA_CLK_COUNT11_0_a2_2 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_5 ;
    wire TICK50_c;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_6 ;
    wire \U409_TICK.COUNTER50Z0Z_8 ;
    wire \U409_TICK.COUNTER50Z0Z_2 ;
    wire \U409_TICK.COUNTER50Z0Z_1 ;
    wire \U409_TICK.COUNTER50Z0Z_16 ;
    wire \U409_TICK.COUNTER50Z0Z_7 ;
    wire \U409_TICK.COUNTER50Z0Z_4 ;
    wire \U409_TICK.TICK503_10_cascade_ ;
    wire \U409_TICK.COUNTER50Z0Z_5 ;
    wire \U409_TICK.COUNTER50Z0Z_3 ;
    wire \U409_TICK.COUNTER50Z0Z_0 ;
    wire \U409_TICK.COUNTER50Z0Z_12 ;
    wire \U409_TICK.TICK503_11 ;
    wire \U409_TICK.TICK503_8_cascade_ ;
    wire \U409_TICK.COUNTER50Z0Z_10 ;
    wire \U409_TICK.TICK503_14_cascade_ ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER50Z0Z_15 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_13 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_14 ;
    wire \U409_TICK.COUNTER50Z0Z_14 ;
    wire \U409_TICK.COUNTER50Z0Z_6 ;
    wire \U409_TICK.COUNTER50Z0Z_13 ;
    wire \U409_TICK.TICK503_9_cascade_ ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_11 ;
    wire \U409_TICK.COUNTER50Z0Z_11 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_9 ;
    wire \U409_TICK.TICK503_10 ;
    wire \U409_TICK.TICK503_14 ;
    wire \U409_TICK.TICK503_9 ;
    wire \U409_TICK.COUNTER50Z0Z_9 ;
    wire CLK6_c_g;
    wire CONSTANT_ONE_NET;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="SIMPLE";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0001111;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE pll (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__8292),
            .RESETB(N__10619),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(CLK80_OUT));
    PRE_IO_GBUF CLK28_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__11400),
            .GLOBALBUFFEROUTPUT(CLK28_IN_c_g));
    IO_PAD CLK28_IN_ibuf_gb_io_iopad (
            .OE(N__11402),
            .DIN(N__11401),
            .DOUT(N__11400),
            .PACKAGEPIN(CLK28_IN));
    defparam CLK28_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK28_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK28_IN_ibuf_gb_io_preio (
            .PADOEN(N__11402),
            .PADOUT(N__11401),
            .PADIN(N__11400),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK6_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__11390),
            .GLOBALBUFFEROUTPUT(CLK6_c_g));
    IO_PAD CLK6_ibuf_gb_io_iopad (
            .OE(N__11392),
            .DIN(N__11391),
            .DOUT(N__11390),
            .PACKAGEPIN(CLK6));
    defparam CLK6_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK6_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK6_ibuf_gb_io_preio (
            .PADOEN(N__11392),
            .PADOUT(N__11391),
            .PADIN(N__11390),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK40_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__11380),
            .GLOBALBUFFEROUTPUT(CLK40_IN_c_g));
    IO_PAD CLK40_IN_ibuf_gb_io_iopad (
            .OE(N__11382),
            .DIN(N__11381),
            .DOUT(N__11380),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_gb_io_preio (
            .PADOEN(N__11382),
            .PADOUT(N__11381),
            .PADIN(N__11380),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__11371),
            .DIN(N__11370),
            .DOUT(N__11369),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__11371),
            .PADOUT(N__11370),
            .PADIN(N__11369),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_0_iopad (
            .OE(N__11362),
            .DIN(N__11361),
            .DOUT(N__11360),
            .PACKAGEPIN(TT[0]));
    defparam TT_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_0_preio (
            .PADOEN(N__11362),
            .PADOUT(N__11361),
            .PADIN(N__11360),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_P1_obuf_iopad (
            .OE(N__11353),
            .DIN(N__11352),
            .DOUT(N__11351),
            .PACKAGEPIN(PIO_P1));
    defparam PIO_P1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_P1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_P1_obuf_preio (
            .PADOEN(N__11353),
            .PADOUT(N__11352),
            .PADIN(N__11351),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10623),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_7_iopad (
            .OE(N__11344),
            .DIN(N__11343),
            .DOUT(N__11342),
            .PACKAGEPIN(D[7]));
    defparam D_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_7_preio (
            .PADOEN(N__11344),
            .PADOUT(N__11343),
            .PADIN(N__11342),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5328),
            .DIN0(D_in_7),
            .DOUT0(N__5907),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__11335),
            .DIN(N__11334),
            .DOUT(N__11333),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__11335),
            .PADOUT(N__11334),
            .PADIN(N__11333),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CPUCONFn_ibuf_iopad (
            .OE(N__11326),
            .DIN(N__11325),
            .DOUT(N__11324),
            .PACKAGEPIN(CPUCONFn));
    defparam CPUCONFn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CPUCONFn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CPUCONFn_ibuf_preio (
            .PADOEN(N__11326),
            .PADOUT(N__11325),
            .PADIN(N__11324),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CPUCONFn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RTC_ENn_obuf_iopad (
            .OE(N__11317),
            .DIN(N__11316),
            .DOUT(N__11315),
            .PACKAGEPIN(RTC_ENn));
    defparam RTC_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RTC_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RTC_ENn_obuf_preio (
            .PADOEN(N__11317),
            .PADOUT(N__11316),
            .PADIN(N__11315),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6639),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_24_iopad (
            .OE(N__11308),
            .DIN(N__11307),
            .DOUT(N__11306),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__11308),
            .PADOUT(N__11307),
            .PADIN(N__11306),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ATA_MODE_P_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ATA_MODE_P_ibuf_iopad (
            .OE(N__11299),
            .DIN(N__11298),
            .DOUT(N__11297),
            .PACKAGEPIN(ATA_MODE_P));
    defparam ATA_MODE_P_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ATA_MODE_P_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ATA_MODE_P_ibuf_preio (
            .PADOEN(N__11299),
            .PADOUT(N__11298),
            .PADIN(N__11297),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(PIO_P0_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_4_iopad (
            .OE(N__11290),
            .DIN(N__11289),
            .DOUT(N__11288),
            .PACKAGEPIN(D[4]));
    defparam D_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_4_preio (
            .PADOEN(N__11290),
            .PADOUT(N__11289),
            .PADIN(N__11288),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5306),
            .DIN0(D_in_4),
            .DOUT0(N__4923),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__11281),
            .DIN(N__11280),
            .DOUT(N__11279),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__11281),
            .PADOUT(N__11280),
            .PADIN(N__11279),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TM_ibuf_1_iopad (
            .OE(N__11272),
            .DIN(N__11271),
            .DOUT(N__11270),
            .PACKAGEPIN(TM[1]));
    defparam TM_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TM_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TM_ibuf_1_preio (
            .PADOEN(N__11272),
            .PADOUT(N__11271),
            .PADIN(N__11270),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TM_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_21_iopad (
            .OE(N__11263),
            .DIN(N__11262),
            .DOUT(N__11261),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__11263),
            .PADOUT(N__11262),
            .PADIN(N__11261),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_obuf_iopad (
            .OE(N__11254),
            .DIN(N__11253),
            .DOUT(N__11252),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMSPACEn_obuf_preio (
            .PADOEN(N__11254),
            .PADOUT(N__11253),
            .PADIN(N__11252),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9192),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__11245),
            .DIN(N__11244),
            .DOUT(N__11243),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__11245),
            .PADOUT(N__11244),
            .PADIN(N__11243),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ROMENn_obuf_iopad (
            .OE(N__11236),
            .DIN(N__11235),
            .DOUT(N__11234),
            .PACKAGEPIN(ROMENn));
    defparam ROMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ROMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ROMENn_obuf_preio (
            .PADOEN(N__11236),
            .PADOUT(N__11235),
            .PADIN(N__11234),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8664),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuft_iopad (
            .OE(N__11227),
            .DIN(N__11226),
            .DOUT(N__11225),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TBIn_obuft_preio (
            .PADOEN(N__11227),
            .PADOUT(N__11226),
            .PADIN(N__11225),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8490),
            .DIN0(),
            .DOUT0(N__8258),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam AUTOBOOT_ibuf_iopad.PULLUP=1'b1;
    IO_PAD AUTOBOOT_ibuf_iopad (
            .OE(N__11218),
            .DIN(N__11217),
            .DOUT(N__11216),
            .PACKAGEPIN(AUTOBOOT));
    defparam AUTOBOOT_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AUTOBOOT_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AUTOBOOT_ibuf_preio (
            .PADOEN(N__11218),
            .PADOUT(N__11217),
            .PADIN(N__11216),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AUTOBOOT_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__11209),
            .DIN(N__11208),
            .DOUT(N__11207),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__11209),
            .PADOUT(N__11208),
            .PADIN(N__11207),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORTSIZE_obuf_iopad (
            .OE(N__11200),
            .DIN(N__11199),
            .DOUT(N__11198),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PORTSIZE_obuf_preio (
            .PADOEN(N__11200),
            .PADOUT(N__11199),
            .PADIN(N__11198),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5085),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_P2_obuf_iopad (
            .OE(N__11191),
            .DIN(N__11190),
            .DOUT(N__11189),
            .PACKAGEPIN(PIO_P2));
    defparam PIO_P2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_P2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_P2_obuf_preio (
            .PADOEN(N__11191),
            .PADOUT(N__11190),
            .PADIN(N__11189),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10605),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__11182),
            .DIN(N__11181),
            .DOUT(N__11180),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__11182),
            .PADOUT(N__11181),
            .PADIN(N__11180),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BRIDGE_ENn_obuf_iopad (
            .OE(N__11173),
            .DIN(N__11172),
            .DOUT(N__11171),
            .PACKAGEPIN(BRIDGE_ENn));
    defparam BRIDGE_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BRIDGE_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BRIDGE_ENn_obuf_preio (
            .PADOEN(N__11173),
            .PADOUT(N__11172),
            .PADIN(N__11171),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5472),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_22_iopad (
            .OE(N__11164),
            .DIN(N__11163),
            .DOUT(N__11162),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__11164),
            .PADOUT(N__11163),
            .PADIN(N__11162),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__11155),
            .DIN(N__11154),
            .DOUT(N__11153),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__11155),
            .PADOUT(N__11154),
            .PADIN(N__11153),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__11146),
            .DIN(N__11145),
            .DOUT(N__11144),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__11146),
            .PADOUT(N__11145),
            .PADIN(N__11144),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_25_iopad (
            .OE(N__11137),
            .DIN(N__11136),
            .DOUT(N__11135),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__11137),
            .PADOUT(N__11136),
            .PADIN(N__11135),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS0n_obuf_iopad (
            .OE(N__11128),
            .DIN(N__11127),
            .DOUT(N__11126),
            .PACKAGEPIN(CIACS0n));
    defparam CIACS0n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS0n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS0n_obuf_preio (
            .PADOEN(N__11128),
            .PADOUT(N__11127),
            .PADIN(N__11126),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8757),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK50_obuf_iopad (
            .OE(N__11119),
            .DIN(N__11118),
            .DOUT(N__11117),
            .PACKAGEPIN(TICK50));
    defparam TICK50_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK50_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK50_obuf_preio (
            .PADOEN(N__11119),
            .PADOUT(N__11118),
            .PADIN(N__11117),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10185),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__11110),
            .DIN(N__11109),
            .DOUT(N__11108),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__11110),
            .PADOUT(N__11109),
            .PADIN(N__11108),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_28_iopad (
            .OE(N__11101),
            .DIN(N__11100),
            .DOUT(N__11099),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__11101),
            .PADOUT(N__11100),
            .PADIN(N__11099),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_30_iopad (
            .OE(N__11092),
            .DIN(N__11091),
            .DOUT(N__11090),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__11092),
            .PADOUT(N__11091),
            .PADIN(N__11090),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD OVL_ibuf_iopad (
            .OE(N__11083),
            .DIN(N__11082),
            .DOUT(N__11081),
            .PACKAGEPIN(OVL));
    defparam OVL_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam OVL_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO OVL_ibuf_preio (
            .PADOEN(N__11083),
            .PADOUT(N__11082),
            .PADIN(N__11081),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(OVL_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuft_iopad (
            .OE(N__11074),
            .DIN(N__11073),
            .DOUT(N__11072),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TCIn_obuft_preio (
            .PADOEN(N__11074),
            .PADOUT(N__11073),
            .PADIN(N__11072),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8406),
            .DIN0(),
            .DOUT0(N__8259),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_5_iopad (
            .OE(N__11065),
            .DIN(N__11064),
            .DOUT(N__11063),
            .PACKAGEPIN(D[5]));
    defparam D_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_5_preio (
            .PADOEN(N__11065),
            .PADOUT(N__11064),
            .PADIN(N__11063),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5323),
            .DIN0(D_in_5),
            .DOUT0(N__5487),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__11056),
            .DIN(N__11055),
            .DOUT(N__11054),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__11056),
            .PADOUT(N__11055),
            .PADIN(N__11054),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__11047),
            .DIN(N__11046),
            .DOUT(N__11045),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__11047),
            .PADOUT(N__11046),
            .PADIN(N__11045),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__11038),
            .DIN(N__11037),
            .DOUT(N__11036),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__11038),
            .PADOUT(N__11037),
            .PADIN(N__11036),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CONFIGENn_obuf_iopad (
            .OE(N__11029),
            .DIN(N__11028),
            .DOUT(N__11027),
            .PACKAGEPIN(CONFIGENn));
    defparam CONFIGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CONFIGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CONFIGENn_obuf_preio (
            .PADOEN(N__11029),
            .PADOUT(N__11028),
            .PADIN(N__11027),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7212),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK60_obuf_iopad (
            .OE(N__11020),
            .DIN(N__11019),
            .DOUT(N__11018),
            .PACKAGEPIN(TICK60));
    defparam TICK60_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK60_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK60_obuf_preio (
            .PADOEN(N__11020),
            .PADOUT(N__11019),
            .PADIN(N__11018),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9597),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_26_iopad (
            .OE(N__11011),
            .DIN(N__11010),
            .DOUT(N__11009),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__11011),
            .PADOUT(N__11010),
            .PADIN(N__11009),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_P0_obuf_iopad (
            .OE(N__11002),
            .DIN(N__11001),
            .DOUT(N__11000),
            .PACKAGEPIN(PIO_P0));
    defparam PIO_P0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_P0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_P0_obuf_preio (
            .PADOEN(N__11002),
            .PADOUT(N__11001),
            .PADIN(N__11000),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4155),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ATA_MODE_S_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ATA_MODE_S_ibuf_iopad (
            .OE(N__10993),
            .DIN(N__10992),
            .DOUT(N__10991),
            .PACKAGEPIN(ATA_MODE_S));
    defparam ATA_MODE_S_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ATA_MODE_S_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ATA_MODE_S_ibuf_preio (
            .PADOEN(N__10993),
            .PADOUT(N__10992),
            .PADIN(N__10991),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(PIO_S0_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_23_iopad (
            .OE(N__10984),
            .DIN(N__10983),
            .DOUT(N__10982),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__10984),
            .PADOUT(N__10983),
            .PADIN(N__10982),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ATA_ENn_obuf_iopad (
            .OE(N__10975),
            .DIN(N__10974),
            .DOUT(N__10973),
            .PACKAGEPIN(ATA_ENn));
    defparam ATA_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ATA_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ATA_ENn_obuf_preio (
            .PADOEN(N__10975),
            .PADOUT(N__10974),
            .PADIN(N__10973),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6468),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_31_iopad (
            .OE(N__10966),
            .DIN(N__10965),
            .DOUT(N__10964),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__10966),
            .PADOUT(N__10965),
            .PADIN(N__10964),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS1n_obuf_iopad (
            .OE(N__10957),
            .DIN(N__10956),
            .DOUT(N__10955),
            .PACKAGEPIN(CIACS1n));
    defparam CIACS1n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS1n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS1n_obuf_preio (
            .PADOEN(N__10957),
            .PADOUT(N__10956),
            .PADIN(N__10955),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7989),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_obuf_iopad (
            .OE(N__10948),
            .DIN(N__10947),
            .DOUT(N__10946),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGSPACEn_obuf_preio (
            .PADOEN(N__10948),
            .PADOUT(N__10947),
            .PADIN(N__10946),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4989),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__10939),
            .DIN(N__10938),
            .DOUT(N__10937),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__10939),
            .PADOUT(N__10938),
            .PADIN(N__10937),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_CIA_obuf_iopad (
            .OE(N__10930),
            .DIN(N__10929),
            .DOUT(N__10928),
            .PACKAGEPIN(CLK_CIA));
    defparam CLK_CIA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_CIA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_CIA_obuf_preio (
            .PADOEN(N__10930),
            .PADOUT(N__10929),
            .PADIN(N__10928),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9564),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__10921),
            .DIN(N__10920),
            .DOUT(N__10919),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__10921),
            .PADOUT(N__10920),
            .PADIN(N__10919),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__10912),
            .DIN(N__10911),
            .DOUT(N__10910),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__10912),
            .PADOUT(N__10911),
            .PADIN(N__10910),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8486),
            .DIN0(TACKn_in),
            .DOUT0(N__8246),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_1_iopad (
            .OE(N__10903),
            .DIN(N__10902),
            .DOUT(N__10901),
            .PACKAGEPIN(TT[1]));
    defparam TT_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_1_preio (
            .PADOEN(N__10903),
            .PADOUT(N__10902),
            .PADIN(N__10901),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__10894),
            .DIN(N__10893),
            .DOUT(N__10892),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__10894),
            .PADOUT(N__10893),
            .PADIN(N__10892),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8022),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_S0_obuf_iopad (
            .OE(N__10885),
            .DIN(N__10884),
            .DOUT(N__10883),
            .PACKAGEPIN(PIO_S0));
    defparam PIO_S0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_S0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_S0_obuf_preio (
            .PADOEN(N__10885),
            .PADOUT(N__10884),
            .PADIN(N__10883),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4134),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_29_iopad (
            .OE(N__10876),
            .DIN(N__10875),
            .DOUT(N__10874),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__10876),
            .PADOUT(N__10875),
            .PADIN(N__10874),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_S2_obuf_iopad (
            .OE(N__10867),
            .DIN(N__10866),
            .DOUT(N__10865),
            .PACKAGEPIN(PIO_S2));
    defparam PIO_S2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_S2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_S2_obuf_preio (
            .PADOEN(N__10867),
            .PADOUT(N__10866),
            .PADIN(N__10865),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10618),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_6_iopad (
            .OE(N__10858),
            .DIN(N__10857),
            .DOUT(N__10856),
            .PACKAGEPIN(D[6]));
    defparam D_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_6_preio (
            .PADOEN(N__10858),
            .PADOUT(N__10857),
            .PADIN(N__10856),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5324),
            .DIN0(D_in_6),
            .DOUT0(N__6339),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__10849),
            .DIN(N__10848),
            .DOUT(N__10847),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__10849),
            .PADOUT(N__10848),
            .PADIN(N__10847),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_27_iopad (
            .OE(N__10840),
            .DIN(N__10839),
            .DOUT(N__10838),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__10840),
            .PADOUT(N__10839),
            .PADIN(N__10838),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_S1_obuf_iopad (
            .OE(N__10831),
            .DIN(N__10830),
            .DOUT(N__10829),
            .PACKAGEPIN(PIO_S1));
    defparam PIO_S1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_S1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_S1_obuf_preio (
            .PADOEN(N__10831),
            .PADOUT(N__10830),
            .PADIN(N__10829),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10598),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TM_ibuf_0_iopad (
            .OE(N__10822),
            .DIN(N__10821),
            .DOUT(N__10820),
            .PACKAGEPIN(TM[0]));
    defparam TM_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TM_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TM_ibuf_0_preio (
            .PADOEN(N__10822),
            .PADOUT(N__10821),
            .PADIN(N__10820),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TM_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__10813),
            .DIN(N__10812),
            .DOUT(N__10811),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__10813),
            .PADOUT(N__10812),
            .PADIN(N__10811),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__10804),
            .DIN(N__10803),
            .DOUT(N__10802),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__10804),
            .PADOUT(N__10803),
            .PADIN(N__10802),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2593 (
            .O(N__10785),
            .I(N__10782));
    LocalMux I__2592 (
            .O(N__10782),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ));
    InMux I__2591 (
            .O(N__10779),
            .I(N__10761));
    InMux I__2590 (
            .O(N__10778),
            .I(N__10761));
    InMux I__2589 (
            .O(N__10777),
            .I(N__10761));
    InMux I__2588 (
            .O(N__10776),
            .I(N__10761));
    InMux I__2587 (
            .O(N__10775),
            .I(N__10761));
    InMux I__2586 (
            .O(N__10774),
            .I(N__10754));
    InMux I__2585 (
            .O(N__10773),
            .I(N__10754));
    InMux I__2584 (
            .O(N__10772),
            .I(N__10754));
    LocalMux I__2583 (
            .O(N__10761),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__2582 (
            .O(N__10754),
            .I(\U409_TICK.TICK503_10 ));
    CascadeMux I__2581 (
            .O(N__10749),
            .I(N__10742));
    InMux I__2580 (
            .O(N__10748),
            .I(N__10730));
    InMux I__2579 (
            .O(N__10747),
            .I(N__10730));
    InMux I__2578 (
            .O(N__10746),
            .I(N__10730));
    InMux I__2577 (
            .O(N__10745),
            .I(N__10730));
    InMux I__2576 (
            .O(N__10742),
            .I(N__10721));
    InMux I__2575 (
            .O(N__10741),
            .I(N__10721));
    InMux I__2574 (
            .O(N__10740),
            .I(N__10721));
    InMux I__2573 (
            .O(N__10739),
            .I(N__10721));
    LocalMux I__2572 (
            .O(N__10730),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__2571 (
            .O(N__10721),
            .I(\U409_TICK.TICK503_14 ));
    CascadeMux I__2570 (
            .O(N__10716),
            .I(N__10709));
    CascadeMux I__2569 (
            .O(N__10715),
            .I(N__10706));
    CascadeMux I__2568 (
            .O(N__10714),
            .I(N__10702));
    CascadeMux I__2567 (
            .O(N__10713),
            .I(N__10697));
    InMux I__2566 (
            .O(N__10712),
            .I(N__10688));
    InMux I__2565 (
            .O(N__10709),
            .I(N__10688));
    InMux I__2564 (
            .O(N__10706),
            .I(N__10688));
    InMux I__2563 (
            .O(N__10705),
            .I(N__10688));
    InMux I__2562 (
            .O(N__10702),
            .I(N__10683));
    InMux I__2561 (
            .O(N__10701),
            .I(N__10683));
    InMux I__2560 (
            .O(N__10700),
            .I(N__10678));
    InMux I__2559 (
            .O(N__10697),
            .I(N__10678));
    LocalMux I__2558 (
            .O(N__10688),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__2557 (
            .O(N__10683),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__2556 (
            .O(N__10678),
            .I(\U409_TICK.TICK503_9 ));
    CascadeMux I__2555 (
            .O(N__10671),
            .I(N__10668));
    InMux I__2554 (
            .O(N__10668),
            .I(N__10664));
    InMux I__2553 (
            .O(N__10667),
            .I(N__10661));
    LocalMux I__2552 (
            .O(N__10664),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    LocalMux I__2551 (
            .O(N__10661),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    ClkMux I__2550 (
            .O(N__10656),
            .I(N__10629));
    ClkMux I__2549 (
            .O(N__10655),
            .I(N__10629));
    ClkMux I__2548 (
            .O(N__10654),
            .I(N__10629));
    ClkMux I__2547 (
            .O(N__10653),
            .I(N__10629));
    ClkMux I__2546 (
            .O(N__10652),
            .I(N__10629));
    ClkMux I__2545 (
            .O(N__10651),
            .I(N__10629));
    ClkMux I__2544 (
            .O(N__10650),
            .I(N__10629));
    ClkMux I__2543 (
            .O(N__10649),
            .I(N__10629));
    ClkMux I__2542 (
            .O(N__10648),
            .I(N__10629));
    GlobalMux I__2541 (
            .O(N__10629),
            .I(N__10626));
    gio2CtrlBuf I__2540 (
            .O(N__10626),
            .I(CLK6_c_g));
    IoInMux I__2539 (
            .O(N__10623),
            .I(N__10620));
    LocalMux I__2538 (
            .O(N__10620),
            .I(N__10615));
    IoInMux I__2537 (
            .O(N__10619),
            .I(N__10612));
    IoInMux I__2536 (
            .O(N__10618),
            .I(N__10609));
    IoSpan4Mux I__2535 (
            .O(N__10615),
            .I(N__10606));
    LocalMux I__2534 (
            .O(N__10612),
            .I(N__10602));
    LocalMux I__2533 (
            .O(N__10609),
            .I(N__10599));
    Span4Mux_s2_h I__2532 (
            .O(N__10606),
            .I(N__10595));
    IoInMux I__2531 (
            .O(N__10605),
            .I(N__10592));
    IoSpan4Mux I__2530 (
            .O(N__10602),
            .I(N__10589));
    IoSpan4Mux I__2529 (
            .O(N__10599),
            .I(N__10586));
    IoInMux I__2528 (
            .O(N__10598),
            .I(N__10583));
    Sp12to4 I__2527 (
            .O(N__10595),
            .I(N__10578));
    LocalMux I__2526 (
            .O(N__10592),
            .I(N__10578));
    Sp12to4 I__2525 (
            .O(N__10589),
            .I(N__10575));
    Sp12to4 I__2524 (
            .O(N__10586),
            .I(N__10570));
    LocalMux I__2523 (
            .O(N__10583),
            .I(N__10570));
    Span12Mux_s9_h I__2522 (
            .O(N__10578),
            .I(N__10567));
    Span12Mux_s9_v I__2521 (
            .O(N__10575),
            .I(N__10564));
    Span12Mux_s1_h I__2520 (
            .O(N__10570),
            .I(N__10561));
    Odrv12 I__2519 (
            .O(N__10567),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__2518 (
            .O(N__10564),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__2517 (
            .O(N__10561),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__2516 (
            .O(N__10554),
            .I(\U409_TICK.TICK503_10_cascade_ ));
    InMux I__2515 (
            .O(N__10551),
            .I(N__10547));
    InMux I__2514 (
            .O(N__10550),
            .I(N__10544));
    LocalMux I__2513 (
            .O(N__10547),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    LocalMux I__2512 (
            .O(N__10544),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    InMux I__2511 (
            .O(N__10539),
            .I(N__10535));
    InMux I__2510 (
            .O(N__10538),
            .I(N__10532));
    LocalMux I__2509 (
            .O(N__10535),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    LocalMux I__2508 (
            .O(N__10532),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    CascadeMux I__2507 (
            .O(N__10527),
            .I(N__10521));
    InMux I__2506 (
            .O(N__10526),
            .I(N__10518));
    InMux I__2505 (
            .O(N__10525),
            .I(N__10515));
    InMux I__2504 (
            .O(N__10524),
            .I(N__10512));
    InMux I__2503 (
            .O(N__10521),
            .I(N__10509));
    LocalMux I__2502 (
            .O(N__10518),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__2501 (
            .O(N__10515),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__2500 (
            .O(N__10512),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__2499 (
            .O(N__10509),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    InMux I__2498 (
            .O(N__10500),
            .I(N__10496));
    InMux I__2497 (
            .O(N__10499),
            .I(N__10493));
    LocalMux I__2496 (
            .O(N__10496),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    LocalMux I__2495 (
            .O(N__10493),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    InMux I__2494 (
            .O(N__10488),
            .I(N__10485));
    LocalMux I__2493 (
            .O(N__10485),
            .I(N__10482));
    Odrv4 I__2492 (
            .O(N__10482),
            .I(\U409_TICK.TICK503_11 ));
    CascadeMux I__2491 (
            .O(N__10479),
            .I(\U409_TICK.TICK503_8_cascade_ ));
    InMux I__2490 (
            .O(N__10476),
            .I(N__10472));
    InMux I__2489 (
            .O(N__10475),
            .I(N__10469));
    LocalMux I__2488 (
            .O(N__10472),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    LocalMux I__2487 (
            .O(N__10469),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    CascadeMux I__2486 (
            .O(N__10464),
            .I(\U409_TICK.TICK503_14_cascade_ ));
    InMux I__2485 (
            .O(N__10461),
            .I(N__10458));
    LocalMux I__2484 (
            .O(N__10458),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ));
    InMux I__2483 (
            .O(N__10455),
            .I(N__10451));
    InMux I__2482 (
            .O(N__10454),
            .I(N__10448));
    LocalMux I__2481 (
            .O(N__10451),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    LocalMux I__2480 (
            .O(N__10448),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    InMux I__2479 (
            .O(N__10443),
            .I(N__10440));
    LocalMux I__2478 (
            .O(N__10440),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ));
    InMux I__2477 (
            .O(N__10437),
            .I(N__10434));
    LocalMux I__2476 (
            .O(N__10434),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ));
    InMux I__2475 (
            .O(N__10431),
            .I(N__10427));
    InMux I__2474 (
            .O(N__10430),
            .I(N__10424));
    LocalMux I__2473 (
            .O(N__10427),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    LocalMux I__2472 (
            .O(N__10424),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    InMux I__2471 (
            .O(N__10419),
            .I(N__10415));
    InMux I__2470 (
            .O(N__10418),
            .I(N__10412));
    LocalMux I__2469 (
            .O(N__10415),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    LocalMux I__2468 (
            .O(N__10412),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    InMux I__2467 (
            .O(N__10407),
            .I(N__10403));
    InMux I__2466 (
            .O(N__10406),
            .I(N__10400));
    LocalMux I__2465 (
            .O(N__10403),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    LocalMux I__2464 (
            .O(N__10400),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    CascadeMux I__2463 (
            .O(N__10395),
            .I(\U409_TICK.TICK503_9_cascade_ ));
    InMux I__2462 (
            .O(N__10392),
            .I(N__10389));
    LocalMux I__2461 (
            .O(N__10389),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ));
    InMux I__2460 (
            .O(N__10386),
            .I(N__10382));
    InMux I__2459 (
            .O(N__10385),
            .I(N__10379));
    LocalMux I__2458 (
            .O(N__10382),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    LocalMux I__2457 (
            .O(N__10379),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    CascadeMux I__2456 (
            .O(N__10374),
            .I(\U409_CIA.un1_CIA_CLK_COUNT_2_0_a2_2_cascade_ ));
    InMux I__2455 (
            .O(N__10371),
            .I(N__10367));
    InMux I__2454 (
            .O(N__10370),
            .I(N__10364));
    LocalMux I__2453 (
            .O(N__10367),
            .I(\U409_CIA.N_420 ));
    LocalMux I__2452 (
            .O(N__10364),
            .I(\U409_CIA.N_420 ));
    InMux I__2451 (
            .O(N__10359),
            .I(N__10356));
    LocalMux I__2450 (
            .O(N__10356),
            .I(\U409_CIA.CLK_CIA_RNOZ0Z_1 ));
    CascadeMux I__2449 (
            .O(N__10353),
            .I(N__10345));
    InMux I__2448 (
            .O(N__10352),
            .I(N__10337));
    InMux I__2447 (
            .O(N__10351),
            .I(N__10337));
    InMux I__2446 (
            .O(N__10350),
            .I(N__10337));
    InMux I__2445 (
            .O(N__10349),
            .I(N__10334));
    InMux I__2444 (
            .O(N__10348),
            .I(N__10327));
    InMux I__2443 (
            .O(N__10345),
            .I(N__10327));
    InMux I__2442 (
            .O(N__10344),
            .I(N__10327));
    LocalMux I__2441 (
            .O(N__10337),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__2440 (
            .O(N__10334),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__2439 (
            .O(N__10327),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    CascadeMux I__2438 (
            .O(N__10320),
            .I(N__10313));
    InMux I__2437 (
            .O(N__10319),
            .I(N__10308));
    InMux I__2436 (
            .O(N__10318),
            .I(N__10301));
    InMux I__2435 (
            .O(N__10317),
            .I(N__10301));
    InMux I__2434 (
            .O(N__10316),
            .I(N__10301));
    InMux I__2433 (
            .O(N__10313),
            .I(N__10298));
    InMux I__2432 (
            .O(N__10312),
            .I(N__10293));
    InMux I__2431 (
            .O(N__10311),
            .I(N__10293));
    LocalMux I__2430 (
            .O(N__10308),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__2429 (
            .O(N__10301),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__2428 (
            .O(N__10298),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__2427 (
            .O(N__10293),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    ClkMux I__2426 (
            .O(N__10284),
            .I(N__10275));
    ClkMux I__2425 (
            .O(N__10283),
            .I(N__10275));
    ClkMux I__2424 (
            .O(N__10282),
            .I(N__10275));
    GlobalMux I__2423 (
            .O(N__10275),
            .I(N__10272));
    gio2CtrlBuf I__2422 (
            .O(N__10272),
            .I(CLK28_IN_c_g));
    InMux I__2421 (
            .O(N__10269),
            .I(N__10263));
    InMux I__2420 (
            .O(N__10268),
            .I(N__10260));
    InMux I__2419 (
            .O(N__10267),
            .I(N__10255));
    InMux I__2418 (
            .O(N__10266),
            .I(N__10255));
    LocalMux I__2417 (
            .O(N__10263),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__2416 (
            .O(N__10260),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__2415 (
            .O(N__10255),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    InMux I__2414 (
            .O(N__10248),
            .I(N__10241));
    InMux I__2413 (
            .O(N__10247),
            .I(N__10236));
    InMux I__2412 (
            .O(N__10246),
            .I(N__10236));
    InMux I__2411 (
            .O(N__10245),
            .I(N__10231));
    InMux I__2410 (
            .O(N__10244),
            .I(N__10231));
    LocalMux I__2409 (
            .O(N__10241),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__2408 (
            .O(N__10236),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__2407 (
            .O(N__10231),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    InMux I__2406 (
            .O(N__10224),
            .I(N__10218));
    InMux I__2405 (
            .O(N__10223),
            .I(N__10215));
    InMux I__2404 (
            .O(N__10222),
            .I(N__10210));
    InMux I__2403 (
            .O(N__10221),
            .I(N__10210));
    LocalMux I__2402 (
            .O(N__10218),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__2401 (
            .O(N__10215),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__2400 (
            .O(N__10210),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    InMux I__2399 (
            .O(N__10203),
            .I(N__10200));
    LocalMux I__2398 (
            .O(N__10200),
            .I(\U409_CIA.CIA_CLK_COUNT11_0_a2_2 ));
    CascadeMux I__2397 (
            .O(N__10197),
            .I(N__10194));
    InMux I__2396 (
            .O(N__10194),
            .I(N__10191));
    LocalMux I__2395 (
            .O(N__10191),
            .I(N__10188));
    Odrv4 I__2394 (
            .O(N__10188),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ));
    IoInMux I__2393 (
            .O(N__10185),
            .I(N__10182));
    LocalMux I__2392 (
            .O(N__10182),
            .I(N__10179));
    Span4Mux_s3_v I__2391 (
            .O(N__10179),
            .I(N__10176));
    Span4Mux_v I__2390 (
            .O(N__10176),
            .I(N__10173));
    Span4Mux_h I__2389 (
            .O(N__10173),
            .I(N__10169));
    InMux I__2388 (
            .O(N__10172),
            .I(N__10166));
    Odrv4 I__2387 (
            .O(N__10169),
            .I(TICK50_c));
    LocalMux I__2386 (
            .O(N__10166),
            .I(TICK50_c));
    InMux I__2385 (
            .O(N__10161),
            .I(N__10158));
    LocalMux I__2384 (
            .O(N__10158),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ));
    InMux I__2383 (
            .O(N__10155),
            .I(N__10151));
    InMux I__2382 (
            .O(N__10154),
            .I(N__10148));
    LocalMux I__2381 (
            .O(N__10151),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    LocalMux I__2380 (
            .O(N__10148),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    InMux I__2379 (
            .O(N__10143),
            .I(N__10139));
    InMux I__2378 (
            .O(N__10142),
            .I(N__10136));
    LocalMux I__2377 (
            .O(N__10139),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    LocalMux I__2376 (
            .O(N__10136),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    CascadeMux I__2375 (
            .O(N__10131),
            .I(N__10127));
    CascadeMux I__2374 (
            .O(N__10130),
            .I(N__10124));
    InMux I__2373 (
            .O(N__10127),
            .I(N__10118));
    InMux I__2372 (
            .O(N__10124),
            .I(N__10118));
    InMux I__2371 (
            .O(N__10123),
            .I(N__10115));
    LocalMux I__2370 (
            .O(N__10118),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__2369 (
            .O(N__10115),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    InMux I__2368 (
            .O(N__10110),
            .I(N__10106));
    InMux I__2367 (
            .O(N__10109),
            .I(N__10103));
    LocalMux I__2366 (
            .O(N__10106),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    LocalMux I__2365 (
            .O(N__10103),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    InMux I__2364 (
            .O(N__10098),
            .I(N__10094));
    InMux I__2363 (
            .O(N__10097),
            .I(N__10091));
    LocalMux I__2362 (
            .O(N__10094),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    LocalMux I__2361 (
            .O(N__10091),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    CascadeMux I__2360 (
            .O(N__10086),
            .I(N__10083));
    InMux I__2359 (
            .O(N__10083),
            .I(N__10079));
    InMux I__2358 (
            .O(N__10082),
            .I(N__10076));
    LocalMux I__2357 (
            .O(N__10079),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    LocalMux I__2356 (
            .O(N__10076),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    InMux I__2355 (
            .O(N__10071),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ));
    InMux I__2354 (
            .O(N__10068),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ));
    InMux I__2353 (
            .O(N__10065),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ));
    InMux I__2352 (
            .O(N__10062),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ));
    InMux I__2351 (
            .O(N__10059),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ));
    InMux I__2350 (
            .O(N__10056),
            .I(N__10050));
    InMux I__2349 (
            .O(N__10055),
            .I(N__10050));
    LocalMux I__2348 (
            .O(N__10050),
            .I(\U409_CIA.N_427 ));
    CascadeMux I__2347 (
            .O(N__10047),
            .I(\U409_CIA.N_427_cascade_ ));
    InMux I__2346 (
            .O(N__10044),
            .I(N__10038));
    InMux I__2345 (
            .O(N__10043),
            .I(N__10038));
    LocalMux I__2344 (
            .O(N__10038),
            .I(N__10035));
    Odrv4 I__2343 (
            .O(N__10035),
            .I(\U409_CIA.CIA_CLK_COUNT11 ));
    InMux I__2342 (
            .O(N__10032),
            .I(N__10027));
    InMux I__2341 (
            .O(N__10031),
            .I(N__10022));
    InMux I__2340 (
            .O(N__10030),
            .I(N__10022));
    LocalMux I__2339 (
            .O(N__10027),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__2338 (
            .O(N__10022),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    CascadeMux I__2337 (
            .O(N__10017),
            .I(N__10013));
    InMux I__2336 (
            .O(N__10016),
            .I(N__10009));
    InMux I__2335 (
            .O(N__10013),
            .I(N__10004));
    InMux I__2334 (
            .O(N__10012),
            .I(N__10004));
    LocalMux I__2333 (
            .O(N__10009),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    LocalMux I__2332 (
            .O(N__10004),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    InMux I__2331 (
            .O(N__9999),
            .I(N__9994));
    InMux I__2330 (
            .O(N__9998),
            .I(N__9989));
    InMux I__2329 (
            .O(N__9997),
            .I(N__9989));
    LocalMux I__2328 (
            .O(N__9994),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__2327 (
            .O(N__9989),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    InMux I__2326 (
            .O(N__9984),
            .I(N__9981));
    LocalMux I__2325 (
            .O(N__9981),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ));
    InMux I__2324 (
            .O(N__9978),
            .I(N__9974));
    CascadeMux I__2323 (
            .O(N__9977),
            .I(N__9969));
    LocalMux I__2322 (
            .O(N__9974),
            .I(N__9966));
    InMux I__2321 (
            .O(N__9973),
            .I(N__9961));
    InMux I__2320 (
            .O(N__9972),
            .I(N__9961));
    InMux I__2319 (
            .O(N__9969),
            .I(N__9958));
    Odrv4 I__2318 (
            .O(N__9966),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__2317 (
            .O(N__9961),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__2316 (
            .O(N__9958),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    InMux I__2315 (
            .O(N__9951),
            .I(N__9948));
    LocalMux I__2314 (
            .O(N__9948),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ));
    InMux I__2313 (
            .O(N__9945),
            .I(N__9941));
    InMux I__2312 (
            .O(N__9944),
            .I(N__9938));
    LocalMux I__2311 (
            .O(N__9941),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    LocalMux I__2310 (
            .O(N__9938),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    InMux I__2309 (
            .O(N__9933),
            .I(N__9929));
    InMux I__2308 (
            .O(N__9932),
            .I(N__9926));
    LocalMux I__2307 (
            .O(N__9929),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    LocalMux I__2306 (
            .O(N__9926),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    CascadeMux I__2305 (
            .O(N__9921),
            .I(N__9918));
    InMux I__2304 (
            .O(N__9918),
            .I(N__9915));
    LocalMux I__2303 (
            .O(N__9915),
            .I(N__9911));
    InMux I__2302 (
            .O(N__9914),
            .I(N__9908));
    Odrv4 I__2301 (
            .O(N__9911),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    LocalMux I__2300 (
            .O(N__9908),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    CascadeMux I__2299 (
            .O(N__9903),
            .I(\U409_TICK.TICK603_9_cascade_ ));
    InMux I__2298 (
            .O(N__9900),
            .I(N__9897));
    LocalMux I__2297 (
            .O(N__9897),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ));
    InMux I__2296 (
            .O(N__9894),
            .I(N__9890));
    InMux I__2295 (
            .O(N__9893),
            .I(N__9887));
    LocalMux I__2294 (
            .O(N__9890),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    LocalMux I__2293 (
            .O(N__9887),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    CascadeMux I__2292 (
            .O(N__9882),
            .I(N__9874));
    InMux I__2291 (
            .O(N__9881),
            .I(N__9866));
    InMux I__2290 (
            .O(N__9880),
            .I(N__9866));
    InMux I__2289 (
            .O(N__9879),
            .I(N__9866));
    InMux I__2288 (
            .O(N__9878),
            .I(N__9861));
    InMux I__2287 (
            .O(N__9877),
            .I(N__9861));
    InMux I__2286 (
            .O(N__9874),
            .I(N__9856));
    InMux I__2285 (
            .O(N__9873),
            .I(N__9856));
    LocalMux I__2284 (
            .O(N__9866),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__2283 (
            .O(N__9861),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__2282 (
            .O(N__9856),
            .I(\U409_TICK.TICK603_14 ));
    InMux I__2281 (
            .O(N__9849),
            .I(N__9838));
    InMux I__2280 (
            .O(N__9848),
            .I(N__9838));
    InMux I__2279 (
            .O(N__9847),
            .I(N__9835));
    InMux I__2278 (
            .O(N__9846),
            .I(N__9826));
    InMux I__2277 (
            .O(N__9845),
            .I(N__9826));
    InMux I__2276 (
            .O(N__9844),
            .I(N__9826));
    InMux I__2275 (
            .O(N__9843),
            .I(N__9826));
    LocalMux I__2274 (
            .O(N__9838),
            .I(N__9823));
    LocalMux I__2273 (
            .O(N__9835),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__2272 (
            .O(N__9826),
            .I(\U409_TICK.TICK603_9 ));
    Odrv4 I__2271 (
            .O(N__9823),
            .I(\U409_TICK.TICK603_9 ));
    CascadeMux I__2270 (
            .O(N__9816),
            .I(N__9810));
    CascadeMux I__2269 (
            .O(N__9815),
            .I(N__9807));
    CascadeMux I__2268 (
            .O(N__9814),
            .I(N__9804));
    InMux I__2267 (
            .O(N__9813),
            .I(N__9790));
    InMux I__2266 (
            .O(N__9810),
            .I(N__9790));
    InMux I__2265 (
            .O(N__9807),
            .I(N__9790));
    InMux I__2264 (
            .O(N__9804),
            .I(N__9790));
    InMux I__2263 (
            .O(N__9803),
            .I(N__9790));
    InMux I__2262 (
            .O(N__9802),
            .I(N__9787));
    InMux I__2261 (
            .O(N__9801),
            .I(N__9784));
    LocalMux I__2260 (
            .O(N__9790),
            .I(N__9781));
    LocalMux I__2259 (
            .O(N__9787),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__2258 (
            .O(N__9784),
            .I(\U409_TICK.TICK603_10 ));
    Odrv12 I__2257 (
            .O(N__9781),
            .I(\U409_TICK.TICK603_10 ));
    InMux I__2256 (
            .O(N__9774),
            .I(N__9771));
    LocalMux I__2255 (
            .O(N__9771),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ));
    InMux I__2254 (
            .O(N__9768),
            .I(N__9764));
    InMux I__2253 (
            .O(N__9767),
            .I(N__9761));
    LocalMux I__2252 (
            .O(N__9764),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    LocalMux I__2251 (
            .O(N__9761),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    InMux I__2250 (
            .O(N__9756),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ));
    InMux I__2249 (
            .O(N__9753),
            .I(bfn_14_6_0_));
    InMux I__2248 (
            .O(N__9750),
            .I(\U409_TICK.un2_COUNTER50_1_cry_9 ));
    InMux I__2247 (
            .O(N__9747),
            .I(\U409_TICK.un2_COUNTER50_1_cry_10 ));
    InMux I__2246 (
            .O(N__9744),
            .I(\U409_TICK.un2_COUNTER50_1_cry_11 ));
    InMux I__2245 (
            .O(N__9741),
            .I(\U409_TICK.un2_COUNTER50_1_cry_12 ));
    InMux I__2244 (
            .O(N__9738),
            .I(\U409_TICK.un2_COUNTER50_1_cry_13 ));
    InMux I__2243 (
            .O(N__9735),
            .I(\U409_TICK.un2_COUNTER50_1_cry_14 ));
    InMux I__2242 (
            .O(N__9732),
            .I(\U409_TICK.un2_COUNTER50_1_cry_15 ));
    InMux I__2241 (
            .O(N__9729),
            .I(N__9725));
    InMux I__2240 (
            .O(N__9728),
            .I(N__9722));
    LocalMux I__2239 (
            .O(N__9725),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    LocalMux I__2238 (
            .O(N__9722),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    InMux I__2237 (
            .O(N__9717),
            .I(N__9714));
    LocalMux I__2236 (
            .O(N__9714),
            .I(\U409_TICK.TICK603_8 ));
    InMux I__2235 (
            .O(N__9711),
            .I(N__9708));
    LocalMux I__2234 (
            .O(N__9708),
            .I(N__9705));
    Span4Mux_h I__2233 (
            .O(N__9705),
            .I(N__9702));
    Odrv4 I__2232 (
            .O(N__9702),
            .I(\U409_CIA.VMA_3_0_a2_2 ));
    CascadeMux I__2231 (
            .O(N__9699),
            .I(\U409_CIA.VMA_RNOZ0Z_1_cascade_ ));
    InMux I__2230 (
            .O(N__9696),
            .I(N__9693));
    LocalMux I__2229 (
            .O(N__9693),
            .I(N__9690));
    Span4Mux_v I__2228 (
            .O(N__9690),
            .I(N__9685));
    InMux I__2227 (
            .O(N__9689),
            .I(N__9682));
    InMux I__2226 (
            .O(N__9688),
            .I(N__9679));
    Odrv4 I__2225 (
            .O(N__9685),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__2224 (
            .O(N__9682),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__2223 (
            .O(N__9679),
            .I(\U409_CIA.VMAZ0 ));
    InMux I__2222 (
            .O(N__9672),
            .I(\U409_TICK.un2_COUNTER50_1_cry_1 ));
    InMux I__2221 (
            .O(N__9669),
            .I(\U409_TICK.un2_COUNTER50_1_cry_2 ));
    InMux I__2220 (
            .O(N__9666),
            .I(\U409_TICK.un2_COUNTER50_1_cry_3 ));
    InMux I__2219 (
            .O(N__9663),
            .I(\U409_TICK.un2_COUNTER50_1_cry_4 ));
    InMux I__2218 (
            .O(N__9660),
            .I(\U409_TICK.un2_COUNTER50_1_cry_5 ));
    InMux I__2217 (
            .O(N__9657),
            .I(\U409_TICK.un2_COUNTER50_1_cry_6 ));
    InMux I__2216 (
            .O(N__9654),
            .I(\U409_TICK.un2_COUNTER50_1_cry_7 ));
    InMux I__2215 (
            .O(N__9651),
            .I(\U409_TICK.un3_COUNTER60_1_cry_15 ));
    InMux I__2214 (
            .O(N__9648),
            .I(N__9644));
    InMux I__2213 (
            .O(N__9647),
            .I(N__9641));
    LocalMux I__2212 (
            .O(N__9644),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    LocalMux I__2211 (
            .O(N__9641),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    InMux I__2210 (
            .O(N__9636),
            .I(N__9632));
    InMux I__2209 (
            .O(N__9635),
            .I(N__9629));
    LocalMux I__2208 (
            .O(N__9632),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    LocalMux I__2207 (
            .O(N__9629),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    CascadeMux I__2206 (
            .O(N__9624),
            .I(N__9621));
    InMux I__2205 (
            .O(N__9621),
            .I(N__9618));
    LocalMux I__2204 (
            .O(N__9618),
            .I(N__9614));
    InMux I__2203 (
            .O(N__9617),
            .I(N__9611));
    Odrv12 I__2202 (
            .O(N__9614),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    LocalMux I__2201 (
            .O(N__9611),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    InMux I__2200 (
            .O(N__9606),
            .I(N__9603));
    LocalMux I__2199 (
            .O(N__9603),
            .I(\U409_TICK.TICK603_11 ));
    CascadeMux I__2198 (
            .O(N__9600),
            .I(\U409_TICK.TICK603_14_cascade_ ));
    IoInMux I__2197 (
            .O(N__9597),
            .I(N__9594));
    LocalMux I__2196 (
            .O(N__9594),
            .I(N__9591));
    Span4Mux_s3_v I__2195 (
            .O(N__9591),
            .I(N__9588));
    Span4Mux_v I__2194 (
            .O(N__9588),
            .I(N__9585));
    Span4Mux_v I__2193 (
            .O(N__9585),
            .I(N__9582));
    Span4Mux_h I__2192 (
            .O(N__9582),
            .I(N__9578));
    InMux I__2191 (
            .O(N__9581),
            .I(N__9575));
    Odrv4 I__2190 (
            .O(N__9578),
            .I(TICK60_c));
    LocalMux I__2189 (
            .O(N__9575),
            .I(TICK60_c));
    CascadeMux I__2188 (
            .O(N__9570),
            .I(\U409_CIA.CLK_CIA6_0_a2_0_cascade_ ));
    CascadeMux I__2187 (
            .O(N__9567),
            .I(\U409_CIA.CLK_CIA6_cascade_ ));
    IoInMux I__2186 (
            .O(N__9564),
            .I(N__9561));
    LocalMux I__2185 (
            .O(N__9561),
            .I(N__9558));
    IoSpan4Mux I__2184 (
            .O(N__9558),
            .I(N__9555));
    Span4Mux_s2_v I__2183 (
            .O(N__9555),
            .I(N__9552));
    Span4Mux_v I__2182 (
            .O(N__9552),
            .I(N__9549));
    Sp12to4 I__2181 (
            .O(N__9549),
            .I(N__9544));
    InMux I__2180 (
            .O(N__9548),
            .I(N__9541));
    InMux I__2179 (
            .O(N__9547),
            .I(N__9538));
    Odrv12 I__2178 (
            .O(N__9544),
            .I(CLK_CIA_c));
    LocalMux I__2177 (
            .O(N__9541),
            .I(CLK_CIA_c));
    LocalMux I__2176 (
            .O(N__9538),
            .I(CLK_CIA_c));
    CascadeMux I__2175 (
            .O(N__9531),
            .I(\U409_CIA.un1_CIA_CLK_COUNT_3_0_a2_0_cascade_ ));
    CascadeMux I__2174 (
            .O(N__9528),
            .I(N__9525));
    InMux I__2173 (
            .O(N__9525),
            .I(N__9521));
    InMux I__2172 (
            .O(N__9524),
            .I(N__9518));
    LocalMux I__2171 (
            .O(N__9521),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    LocalMux I__2170 (
            .O(N__9518),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    InMux I__2169 (
            .O(N__9513),
            .I(\U409_TICK.un3_COUNTER60_1_cry_6 ));
    InMux I__2168 (
            .O(N__9510),
            .I(\U409_TICK.un3_COUNTER60_1_cry_7 ));
    InMux I__2167 (
            .O(N__9507),
            .I(bfn_13_7_0_));
    InMux I__2166 (
            .O(N__9504),
            .I(N__9500));
    InMux I__2165 (
            .O(N__9503),
            .I(N__9497));
    LocalMux I__2164 (
            .O(N__9500),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    LocalMux I__2163 (
            .O(N__9497),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    InMux I__2162 (
            .O(N__9492),
            .I(\U409_TICK.un3_COUNTER60_1_cry_9 ));
    InMux I__2161 (
            .O(N__9489),
            .I(\U409_TICK.un3_COUNTER60_1_cry_10 ));
    InMux I__2160 (
            .O(N__9486),
            .I(N__9482));
    InMux I__2159 (
            .O(N__9485),
            .I(N__9479));
    LocalMux I__2158 (
            .O(N__9482),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    LocalMux I__2157 (
            .O(N__9479),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    InMux I__2156 (
            .O(N__9474),
            .I(\U409_TICK.un3_COUNTER60_1_cry_11 ));
    InMux I__2155 (
            .O(N__9471),
            .I(N__9467));
    InMux I__2154 (
            .O(N__9470),
            .I(N__9464));
    LocalMux I__2153 (
            .O(N__9467),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    LocalMux I__2152 (
            .O(N__9464),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    InMux I__2151 (
            .O(N__9459),
            .I(\U409_TICK.un3_COUNTER60_1_cry_12 ));
    InMux I__2150 (
            .O(N__9456),
            .I(\U409_TICK.un3_COUNTER60_1_cry_13 ));
    CascadeMux I__2149 (
            .O(N__9453),
            .I(N__9449));
    InMux I__2148 (
            .O(N__9452),
            .I(N__9446));
    InMux I__2147 (
            .O(N__9449),
            .I(N__9443));
    LocalMux I__2146 (
            .O(N__9446),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    LocalMux I__2145 (
            .O(N__9443),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    InMux I__2144 (
            .O(N__9438),
            .I(N__9435));
    LocalMux I__2143 (
            .O(N__9435),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ));
    InMux I__2142 (
            .O(N__9432),
            .I(\U409_TICK.un3_COUNTER60_1_cry_14 ));
    InMux I__2141 (
            .O(N__9429),
            .I(N__9426));
    LocalMux I__2140 (
            .O(N__9426),
            .I(N__9421));
    SRMux I__2139 (
            .O(N__9425),
            .I(N__9387));
    SRMux I__2138 (
            .O(N__9424),
            .I(N__9387));
    Glb2LocalMux I__2137 (
            .O(N__9421),
            .I(N__9387));
    SRMux I__2136 (
            .O(N__9420),
            .I(N__9387));
    SRMux I__2135 (
            .O(N__9419),
            .I(N__9387));
    SRMux I__2134 (
            .O(N__9418),
            .I(N__9387));
    SRMux I__2133 (
            .O(N__9417),
            .I(N__9387));
    SRMux I__2132 (
            .O(N__9416),
            .I(N__9387));
    SRMux I__2131 (
            .O(N__9415),
            .I(N__9387));
    SRMux I__2130 (
            .O(N__9414),
            .I(N__9387));
    SRMux I__2129 (
            .O(N__9413),
            .I(N__9387));
    SRMux I__2128 (
            .O(N__9412),
            .I(N__9387));
    GlobalMux I__2127 (
            .O(N__9387),
            .I(N__9384));
    gio2CtrlBuf I__2126 (
            .O(N__9384),
            .I(RESETn_c_i_g));
    InMux I__2125 (
            .O(N__9381),
            .I(N__9377));
    InMux I__2124 (
            .O(N__9380),
            .I(N__9374));
    LocalMux I__2123 (
            .O(N__9377),
            .I(N__9369));
    LocalMux I__2122 (
            .O(N__9374),
            .I(N__9369));
    Span4Mux_v I__2121 (
            .O(N__9369),
            .I(N__9366));
    Span4Mux_h I__2120 (
            .O(N__9366),
            .I(N__9362));
    InMux I__2119 (
            .O(N__9365),
            .I(N__9359));
    Sp12to4 I__2118 (
            .O(N__9362),
            .I(N__9356));
    LocalMux I__2117 (
            .O(N__9359),
            .I(N__9353));
    Span12Mux_h I__2116 (
            .O(N__9356),
            .I(N__9350));
    Span12Mux_v I__2115 (
            .O(N__9353),
            .I(N__9347));
    Span12Mux_v I__2114 (
            .O(N__9350),
            .I(N__9342));
    Span12Mux_h I__2113 (
            .O(N__9347),
            .I(N__9342));
    Odrv12 I__2112 (
            .O(N__9342),
            .I(OVL_c));
    InMux I__2111 (
            .O(N__9339),
            .I(N__9336));
    LocalMux I__2110 (
            .O(N__9336),
            .I(N__9332));
    CascadeMux I__2109 (
            .O(N__9335),
            .I(N__9329));
    Span4Mux_v I__2108 (
            .O(N__9332),
            .I(N__9325));
    InMux I__2107 (
            .O(N__9329),
            .I(N__9322));
    InMux I__2106 (
            .O(N__9328),
            .I(N__9319));
    Odrv4 I__2105 (
            .O(N__9325),
            .I(N_429));
    LocalMux I__2104 (
            .O(N__9322),
            .I(N_429));
    LocalMux I__2103 (
            .O(N__9319),
            .I(N_429));
    CascadeMux I__2102 (
            .O(N__9312),
            .I(N__9309));
    InMux I__2101 (
            .O(N__9309),
            .I(N__9305));
    InMux I__2100 (
            .O(N__9308),
            .I(N__9298));
    LocalMux I__2099 (
            .O(N__9305),
            .I(N__9295));
    InMux I__2098 (
            .O(N__9304),
            .I(N__9290));
    InMux I__2097 (
            .O(N__9303),
            .I(N__9290));
    InMux I__2096 (
            .O(N__9302),
            .I(N__9287));
    InMux I__2095 (
            .O(N__9301),
            .I(N__9284));
    LocalMux I__2094 (
            .O(N__9298),
            .I(N__9281));
    Span4Mux_h I__2093 (
            .O(N__9295),
            .I(N__9272));
    LocalMux I__2092 (
            .O(N__9290),
            .I(N__9272));
    LocalMux I__2091 (
            .O(N__9287),
            .I(N__9272));
    LocalMux I__2090 (
            .O(N__9284),
            .I(N__9272));
    Span4Mux_v I__2089 (
            .O(N__9281),
            .I(N__9267));
    Span4Mux_v I__2088 (
            .O(N__9272),
            .I(N__9264));
    InMux I__2087 (
            .O(N__9271),
            .I(N__9261));
    InMux I__2086 (
            .O(N__9270),
            .I(N__9258));
    Odrv4 I__2085 (
            .O(N__9267),
            .I(N_348));
    Odrv4 I__2084 (
            .O(N__9264),
            .I(N_348));
    LocalMux I__2083 (
            .O(N__9261),
            .I(N_348));
    LocalMux I__2082 (
            .O(N__9258),
            .I(N_348));
    CascadeMux I__2081 (
            .O(N__9249),
            .I(N__9243));
    InMux I__2080 (
            .O(N__9248),
            .I(N__9240));
    InMux I__2079 (
            .O(N__9247),
            .I(N__9237));
    InMux I__2078 (
            .O(N__9246),
            .I(N__9231));
    InMux I__2077 (
            .O(N__9243),
            .I(N__9231));
    LocalMux I__2076 (
            .O(N__9240),
            .I(N__9227));
    LocalMux I__2075 (
            .O(N__9237),
            .I(N__9224));
    InMux I__2074 (
            .O(N__9236),
            .I(N__9221));
    LocalMux I__2073 (
            .O(N__9231),
            .I(N__9218));
    InMux I__2072 (
            .O(N__9230),
            .I(N__9215));
    Span4Mux_h I__2071 (
            .O(N__9227),
            .I(N__9208));
    Span4Mux_v I__2070 (
            .O(N__9224),
            .I(N__9208));
    LocalMux I__2069 (
            .O(N__9221),
            .I(N__9208));
    Span12Mux_v I__2068 (
            .O(N__9218),
            .I(N__9205));
    LocalMux I__2067 (
            .O(N__9215),
            .I(N__9202));
    Span4Mux_v I__2066 (
            .O(N__9208),
            .I(N__9199));
    Odrv12 I__2065 (
            .O(N__9205),
            .I(N_156_i));
    Odrv12 I__2064 (
            .O(N__9202),
            .I(N_156_i));
    Odrv4 I__2063 (
            .O(N__9199),
            .I(N_156_i));
    IoInMux I__2062 (
            .O(N__9192),
            .I(N__9189));
    LocalMux I__2061 (
            .O(N__9189),
            .I(N__9186));
    Span12Mux_s11_v I__2060 (
            .O(N__9186),
            .I(N__9183));
    Odrv12 I__2059 (
            .O(N__9183),
            .I(N_264_i));
    InMux I__2058 (
            .O(N__9180),
            .I(N__9174));
    CascadeMux I__2057 (
            .O(N__9179),
            .I(N__9171));
    CascadeMux I__2056 (
            .O(N__9178),
            .I(N__9164));
    CascadeMux I__2055 (
            .O(N__9177),
            .I(N__9160));
    LocalMux I__2054 (
            .O(N__9174),
            .I(N__9155));
    InMux I__2053 (
            .O(N__9171),
            .I(N__9152));
    InMux I__2052 (
            .O(N__9170),
            .I(N__9149));
    InMux I__2051 (
            .O(N__9169),
            .I(N__9146));
    InMux I__2050 (
            .O(N__9168),
            .I(N__9137));
    InMux I__2049 (
            .O(N__9167),
            .I(N__9137));
    InMux I__2048 (
            .O(N__9164),
            .I(N__9137));
    InMux I__2047 (
            .O(N__9163),
            .I(N__9137));
    InMux I__2046 (
            .O(N__9160),
            .I(N__9132));
    InMux I__2045 (
            .O(N__9159),
            .I(N__9127));
    InMux I__2044 (
            .O(N__9158),
            .I(N__9127));
    Span4Mux_h I__2043 (
            .O(N__9155),
            .I(N__9122));
    LocalMux I__2042 (
            .O(N__9152),
            .I(N__9122));
    LocalMux I__2041 (
            .O(N__9149),
            .I(N__9119));
    LocalMux I__2040 (
            .O(N__9146),
            .I(N__9114));
    LocalMux I__2039 (
            .O(N__9137),
            .I(N__9114));
    InMux I__2038 (
            .O(N__9136),
            .I(N__9111));
    InMux I__2037 (
            .O(N__9135),
            .I(N__9108));
    LocalMux I__2036 (
            .O(N__9132),
            .I(N__9100));
    LocalMux I__2035 (
            .O(N__9127),
            .I(N__9100));
    Span4Mux_v I__2034 (
            .O(N__9122),
            .I(N__9090));
    Span4Mux_h I__2033 (
            .O(N__9119),
            .I(N__9090));
    Span4Mux_h I__2032 (
            .O(N__9114),
            .I(N__9090));
    LocalMux I__2031 (
            .O(N__9111),
            .I(N__9090));
    LocalMux I__2030 (
            .O(N__9108),
            .I(N__9087));
    InMux I__2029 (
            .O(N__9107),
            .I(N__9084));
    InMux I__2028 (
            .O(N__9106),
            .I(N__9079));
    InMux I__2027 (
            .O(N__9105),
            .I(N__9079));
    Span4Mux_h I__2026 (
            .O(N__9100),
            .I(N__9076));
    InMux I__2025 (
            .O(N__9099),
            .I(N__9073));
    Span4Mux_v I__2024 (
            .O(N__9090),
            .I(N__9067));
    Span4Mux_h I__2023 (
            .O(N__9087),
            .I(N__9062));
    LocalMux I__2022 (
            .O(N__9084),
            .I(N__9062));
    LocalMux I__2021 (
            .O(N__9079),
            .I(N__9059));
    Span4Mux_h I__2020 (
            .O(N__9076),
            .I(N__9056));
    LocalMux I__2019 (
            .O(N__9073),
            .I(N__9053));
    InMux I__2018 (
            .O(N__9072),
            .I(N__9050));
    InMux I__2017 (
            .O(N__9071),
            .I(N__9045));
    InMux I__2016 (
            .O(N__9070),
            .I(N__9045));
    Span4Mux_h I__2015 (
            .O(N__9067),
            .I(N__9037));
    Span4Mux_v I__2014 (
            .O(N__9062),
            .I(N__9037));
    Span4Mux_v I__2013 (
            .O(N__9059),
            .I(N__9037));
    Sp12to4 I__2012 (
            .O(N__9056),
            .I(N__9028));
    Span12Mux_s7_v I__2011 (
            .O(N__9053),
            .I(N__9028));
    LocalMux I__2010 (
            .O(N__9050),
            .I(N__9028));
    LocalMux I__2009 (
            .O(N__9045),
            .I(N__9028));
    InMux I__2008 (
            .O(N__9044),
            .I(N__9025));
    Sp12to4 I__2007 (
            .O(N__9037),
            .I(N__9018));
    Span12Mux_v I__2006 (
            .O(N__9028),
            .I(N__9018));
    LocalMux I__2005 (
            .O(N__9025),
            .I(N__9018));
    Span12Mux_v I__2004 (
            .O(N__9018),
            .I(N__9015));
    Span12Mux_h I__2003 (
            .O(N__9015),
            .I(N__9012));
    Odrv12 I__2002 (
            .O(N__9012),
            .I(RESETn_c));
    IoInMux I__2001 (
            .O(N__9009),
            .I(N__9006));
    LocalMux I__2000 (
            .O(N__9006),
            .I(N__9003));
    Odrv12 I__1999 (
            .O(N__9003),
            .I(RESETn_c_i));
    CascadeMux I__1998 (
            .O(N__9000),
            .I(N__8996));
    InMux I__1997 (
            .O(N__8999),
            .I(N__8991));
    InMux I__1996 (
            .O(N__8996),
            .I(N__8991));
    LocalMux I__1995 (
            .O(N__8991),
            .I(N__8987));
    InMux I__1994 (
            .O(N__8990),
            .I(N__8984));
    Odrv4 I__1993 (
            .O(N__8987),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__1992 (
            .O(N__8984),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    InMux I__1991 (
            .O(N__8979),
            .I(N__8975));
    InMux I__1990 (
            .O(N__8978),
            .I(N__8972));
    LocalMux I__1989 (
            .O(N__8975),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    LocalMux I__1988 (
            .O(N__8972),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    InMux I__1987 (
            .O(N__8967),
            .I(\U409_TICK.un3_COUNTER60_1_cry_1 ));
    InMux I__1986 (
            .O(N__8964),
            .I(\U409_TICK.un3_COUNTER60_1_cry_2 ));
    InMux I__1985 (
            .O(N__8961),
            .I(\U409_TICK.un3_COUNTER60_1_cry_3 ));
    InMux I__1984 (
            .O(N__8958),
            .I(\U409_TICK.un3_COUNTER60_1_cry_4 ));
    CascadeMux I__1983 (
            .O(N__8955),
            .I(N__8952));
    InMux I__1982 (
            .O(N__8952),
            .I(N__8949));
    LocalMux I__1981 (
            .O(N__8949),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ));
    InMux I__1980 (
            .O(N__8946),
            .I(\U409_TICK.un3_COUNTER60_1_cry_5 ));
    CascadeMux I__1979 (
            .O(N__8943),
            .I(\U409_TRANSFER_ACK.m12_i_0_cascade_ ));
    InMux I__1978 (
            .O(N__8940),
            .I(N__8937));
    LocalMux I__1977 (
            .O(N__8937),
            .I(\U409_TRANSFER_ACK.N_293 ));
    InMux I__1976 (
            .O(N__8934),
            .I(N__8931));
    LocalMux I__1975 (
            .O(N__8931),
            .I(\U409_TRANSFER_ACK.N_191 ));
    CascadeMux I__1974 (
            .O(N__8928),
            .I(\U409_TRANSFER_ACK.N_191_cascade_ ));
    InMux I__1973 (
            .O(N__8925),
            .I(N__8922));
    LocalMux I__1972 (
            .O(N__8922),
            .I(\U409_TRANSFER_ACK.N_223 ));
    CascadeMux I__1971 (
            .O(N__8919),
            .I(\U409_TRANSFER_ACK.i5_mux_cascade_ ));
    InMux I__1970 (
            .O(N__8916),
            .I(N__8913));
    LocalMux I__1969 (
            .O(N__8913),
            .I(N__8905));
    InMux I__1968 (
            .O(N__8912),
            .I(N__8900));
    InMux I__1967 (
            .O(N__8911),
            .I(N__8900));
    InMux I__1966 (
            .O(N__8910),
            .I(N__8897));
    InMux I__1965 (
            .O(N__8909),
            .I(N__8892));
    InMux I__1964 (
            .O(N__8908),
            .I(N__8892));
    Odrv4 I__1963 (
            .O(N__8905),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__1962 (
            .O(N__8900),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__1961 (
            .O(N__8897),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__1960 (
            .O(N__8892),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    CascadeMux I__1959 (
            .O(N__8883),
            .I(N__8880));
    InMux I__1958 (
            .O(N__8880),
            .I(N__8877));
    LocalMux I__1957 (
            .O(N__8877),
            .I(N__8870));
    InMux I__1956 (
            .O(N__8876),
            .I(N__8863));
    InMux I__1955 (
            .O(N__8875),
            .I(N__8863));
    InMux I__1954 (
            .O(N__8874),
            .I(N__8863));
    InMux I__1953 (
            .O(N__8873),
            .I(N__8860));
    Odrv4 I__1952 (
            .O(N__8870),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__1951 (
            .O(N__8863),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__1950 (
            .O(N__8860),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    InMux I__1949 (
            .O(N__8853),
            .I(N__8850));
    LocalMux I__1948 (
            .O(N__8850),
            .I(\U409_TRANSFER_ACK.N_290 ));
    InMux I__1947 (
            .O(N__8847),
            .I(N__8841));
    InMux I__1946 (
            .O(N__8846),
            .I(N__8834));
    InMux I__1945 (
            .O(N__8845),
            .I(N__8834));
    InMux I__1944 (
            .O(N__8844),
            .I(N__8834));
    LocalMux I__1943 (
            .O(N__8841),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__1942 (
            .O(N__8834),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    CascadeMux I__1941 (
            .O(N__8829),
            .I(N__8825));
    CascadeMux I__1940 (
            .O(N__8828),
            .I(N__8822));
    InMux I__1939 (
            .O(N__8825),
            .I(N__8814));
    InMux I__1938 (
            .O(N__8822),
            .I(N__8814));
    InMux I__1937 (
            .O(N__8821),
            .I(N__8814));
    LocalMux I__1936 (
            .O(N__8814),
            .I(N__8811));
    Odrv4 I__1935 (
            .O(N__8811),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    InMux I__1934 (
            .O(N__8808),
            .I(N__8802));
    InMux I__1933 (
            .O(N__8807),
            .I(N__8797));
    InMux I__1932 (
            .O(N__8806),
            .I(N__8797));
    InMux I__1931 (
            .O(N__8805),
            .I(N__8794));
    LocalMux I__1930 (
            .O(N__8802),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__1929 (
            .O(N__8797),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__1928 (
            .O(N__8794),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    InMux I__1927 (
            .O(N__8787),
            .I(N__8780));
    InMux I__1926 (
            .O(N__8786),
            .I(N__8780));
    InMux I__1925 (
            .O(N__8785),
            .I(N__8777));
    LocalMux I__1924 (
            .O(N__8780),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    LocalMux I__1923 (
            .O(N__8777),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    CascadeMux I__1922 (
            .O(N__8772),
            .I(CIA_ENABLE_cascade_));
    InMux I__1921 (
            .O(N__8769),
            .I(N__8766));
    LocalMux I__1920 (
            .O(N__8766),
            .I(N__8763));
    Span12Mux_h I__1919 (
            .O(N__8763),
            .I(N__8760));
    Odrv12 I__1918 (
            .O(N__8760),
            .I(A_c_12));
    IoInMux I__1917 (
            .O(N__8757),
            .I(N__8754));
    LocalMux I__1916 (
            .O(N__8754),
            .I(N__8751));
    Span4Mux_s0_h I__1915 (
            .O(N__8751),
            .I(N__8748));
    Span4Mux_h I__1914 (
            .O(N__8748),
            .I(N__8745));
    Sp12to4 I__1913 (
            .O(N__8745),
            .I(N__8742));
    Span12Mux_s8_v I__1912 (
            .O(N__8742),
            .I(N__8739));
    Span12Mux_h I__1911 (
            .O(N__8739),
            .I(N__8736));
    Odrv12 I__1910 (
            .O(N__8736),
            .I(U409_ADDRESS_DECODE_un1_CIACS0n_i));
    CascadeMux I__1909 (
            .O(N__8733),
            .I(\U409_TICK.TICK603_10_cascade_ ));
    CascadeMux I__1908 (
            .O(N__8730),
            .I(\U409_TRANSFER_ACK.m12_i_a2_1_0_cascade_ ));
    CascadeMux I__1907 (
            .O(N__8727),
            .I(N__8724));
    InMux I__1906 (
            .O(N__8724),
            .I(N__8721));
    LocalMux I__1905 (
            .O(N__8721),
            .I(\U409_TRANSFER_ACK.N_379 ));
    InMux I__1904 (
            .O(N__8718),
            .I(N__8715));
    LocalMux I__1903 (
            .O(N__8715),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0 ));
    InMux I__1902 (
            .O(N__8712),
            .I(N__8709));
    LocalMux I__1901 (
            .O(N__8709),
            .I(\U409_TRANSFER_ACK.N_307 ));
    CascadeMux I__1900 (
            .O(N__8706),
            .I(N__8703));
    InMux I__1899 (
            .O(N__8703),
            .I(N__8699));
    InMux I__1898 (
            .O(N__8702),
            .I(N__8695));
    LocalMux I__1897 (
            .O(N__8699),
            .I(N__8692));
    InMux I__1896 (
            .O(N__8698),
            .I(N__8689));
    LocalMux I__1895 (
            .O(N__8695),
            .I(N__8686));
    Span4Mux_v I__1894 (
            .O(N__8692),
            .I(N__8681));
    LocalMux I__1893 (
            .O(N__8689),
            .I(N__8681));
    Odrv4 I__1892 (
            .O(N__8686),
            .I(\U409_TRANSFER_ACK.N_381 ));
    Odrv4 I__1891 (
            .O(N__8681),
            .I(\U409_TRANSFER_ACK.N_381 ));
    InMux I__1890 (
            .O(N__8676),
            .I(N__8673));
    LocalMux I__1889 (
            .O(N__8673),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0 ));
    InMux I__1888 (
            .O(N__8670),
            .I(N__8667));
    LocalMux I__1887 (
            .O(N__8667),
            .I(\U409_TRANSFER_ACK.ROMENn_e_1 ));
    IoInMux I__1886 (
            .O(N__8664),
            .I(N__8661));
    LocalMux I__1885 (
            .O(N__8661),
            .I(N__8658));
    Span4Mux_s2_v I__1884 (
            .O(N__8658),
            .I(N__8655));
    Sp12to4 I__1883 (
            .O(N__8655),
            .I(N__8652));
    Span12Mux_h I__1882 (
            .O(N__8652),
            .I(N__8648));
    CascadeMux I__1881 (
            .O(N__8651),
            .I(N__8645));
    Span12Mux_v I__1880 (
            .O(N__8648),
            .I(N__8642));
    InMux I__1879 (
            .O(N__8645),
            .I(N__8639));
    Odrv12 I__1878 (
            .O(N__8642),
            .I(ROMENn_c));
    LocalMux I__1877 (
            .O(N__8639),
            .I(ROMENn_c));
    CascadeMux I__1876 (
            .O(N__8634),
            .I(N__8627));
    InMux I__1875 (
            .O(N__8633),
            .I(N__8620));
    InMux I__1874 (
            .O(N__8632),
            .I(N__8620));
    InMux I__1873 (
            .O(N__8631),
            .I(N__8617));
    InMux I__1872 (
            .O(N__8630),
            .I(N__8614));
    InMux I__1871 (
            .O(N__8627),
            .I(N__8611));
    InMux I__1870 (
            .O(N__8626),
            .I(N__8608));
    InMux I__1869 (
            .O(N__8625),
            .I(N__8605));
    LocalMux I__1868 (
            .O(N__8620),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1867 (
            .O(N__8617),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1866 (
            .O(N__8614),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1865 (
            .O(N__8611),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1864 (
            .O(N__8608),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1863 (
            .O(N__8605),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    CascadeMux I__1862 (
            .O(N__8592),
            .I(N__8587));
    CascadeMux I__1861 (
            .O(N__8591),
            .I(N__8582));
    InMux I__1860 (
            .O(N__8590),
            .I(N__8578));
    InMux I__1859 (
            .O(N__8587),
            .I(N__8575));
    InMux I__1858 (
            .O(N__8586),
            .I(N__8572));
    InMux I__1857 (
            .O(N__8585),
            .I(N__8569));
    InMux I__1856 (
            .O(N__8582),
            .I(N__8564));
    InMux I__1855 (
            .O(N__8581),
            .I(N__8564));
    LocalMux I__1854 (
            .O(N__8578),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1853 (
            .O(N__8575),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1852 (
            .O(N__8572),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1851 (
            .O(N__8569),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1850 (
            .O(N__8564),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    CascadeMux I__1849 (
            .O(N__8553),
            .I(N__8548));
    InMux I__1848 (
            .O(N__8552),
            .I(N__8540));
    InMux I__1847 (
            .O(N__8551),
            .I(N__8540));
    InMux I__1846 (
            .O(N__8548),
            .I(N__8535));
    InMux I__1845 (
            .O(N__8547),
            .I(N__8535));
    InMux I__1844 (
            .O(N__8546),
            .I(N__8532));
    InMux I__1843 (
            .O(N__8545),
            .I(N__8529));
    LocalMux I__1842 (
            .O(N__8540),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1841 (
            .O(N__8535),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1840 (
            .O(N__8532),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1839 (
            .O(N__8529),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    InMux I__1838 (
            .O(N__8520),
            .I(N__8512));
    InMux I__1837 (
            .O(N__8519),
            .I(N__8507));
    InMux I__1836 (
            .O(N__8518),
            .I(N__8507));
    InMux I__1835 (
            .O(N__8517),
            .I(N__8504));
    InMux I__1834 (
            .O(N__8516),
            .I(N__8499));
    InMux I__1833 (
            .O(N__8515),
            .I(N__8499));
    LocalMux I__1832 (
            .O(N__8512),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1831 (
            .O(N__8507),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1830 (
            .O(N__8504),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1829 (
            .O(N__8499),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    IoInMux I__1828 (
            .O(N__8490),
            .I(N__8487));
    LocalMux I__1827 (
            .O(N__8487),
            .I(N__8483));
    IoInMux I__1826 (
            .O(N__8486),
            .I(N__8480));
    IoSpan4Mux I__1825 (
            .O(N__8483),
            .I(N__8477));
    LocalMux I__1824 (
            .O(N__8480),
            .I(N__8474));
    Span4Mux_s2_v I__1823 (
            .O(N__8477),
            .I(N__8469));
    Span4Mux_s2_v I__1822 (
            .O(N__8474),
            .I(N__8469));
    Span4Mux_v I__1821 (
            .O(N__8469),
            .I(N__8466));
    Sp12to4 I__1820 (
            .O(N__8466),
            .I(N__8461));
    InMux I__1819 (
            .O(N__8465),
            .I(N__8458));
    CascadeMux I__1818 (
            .O(N__8464),
            .I(N__8455));
    Span12Mux_h I__1817 (
            .O(N__8461),
            .I(N__8450));
    LocalMux I__1816 (
            .O(N__8458),
            .I(N__8450));
    InMux I__1815 (
            .O(N__8455),
            .I(N__8447));
    Odrv12 I__1814 (
            .O(N__8450),
            .I(TACK_EN));
    LocalMux I__1813 (
            .O(N__8447),
            .I(TACK_EN));
    InMux I__1812 (
            .O(N__8442),
            .I(N__8439));
    LocalMux I__1811 (
            .O(N__8439),
            .I(N__8435));
    InMux I__1810 (
            .O(N__8438),
            .I(N__8432));
    Span4Mux_v I__1809 (
            .O(N__8435),
            .I(N__8429));
    LocalMux I__1808 (
            .O(N__8432),
            .I(N__8426));
    Odrv4 I__1807 (
            .O(N__8429),
            .I(N_357));
    Odrv4 I__1806 (
            .O(N__8426),
            .I(N_357));
    InMux I__1805 (
            .O(N__8421),
            .I(N__8418));
    LocalMux I__1804 (
            .O(N__8418),
            .I(N__8414));
    InMux I__1803 (
            .O(N__8417),
            .I(N__8411));
    Odrv4 I__1802 (
            .O(N__8414),
            .I(N_339));
    LocalMux I__1801 (
            .O(N__8411),
            .I(N_339));
    IoInMux I__1800 (
            .O(N__8406),
            .I(N__8403));
    LocalMux I__1799 (
            .O(N__8403),
            .I(N__8400));
    IoSpan4Mux I__1798 (
            .O(N__8400),
            .I(N__8397));
    IoSpan4Mux I__1797 (
            .O(N__8397),
            .I(N__8394));
    Sp12to4 I__1796 (
            .O(N__8394),
            .I(N__8391));
    Span12Mux_v I__1795 (
            .O(N__8391),
            .I(N__8388));
    Odrv12 I__1794 (
            .O(N__8388),
            .I(TCIn_1_i));
    CascadeMux I__1793 (
            .O(N__8385),
            .I(N__8377));
    CascadeMux I__1792 (
            .O(N__8384),
            .I(N__8374));
    InMux I__1791 (
            .O(N__8383),
            .I(N__8370));
    InMux I__1790 (
            .O(N__8382),
            .I(N__8365));
    InMux I__1789 (
            .O(N__8381),
            .I(N__8365));
    InMux I__1788 (
            .O(N__8380),
            .I(N__8362));
    InMux I__1787 (
            .O(N__8377),
            .I(N__8359));
    InMux I__1786 (
            .O(N__8374),
            .I(N__8354));
    InMux I__1785 (
            .O(N__8373),
            .I(N__8354));
    LocalMux I__1784 (
            .O(N__8370),
            .I(N__8351));
    LocalMux I__1783 (
            .O(N__8365),
            .I(N__8339));
    LocalMux I__1782 (
            .O(N__8362),
            .I(N__8336));
    LocalMux I__1781 (
            .O(N__8359),
            .I(N__8333));
    LocalMux I__1780 (
            .O(N__8354),
            .I(N__8330));
    Glb2LocalMux I__1779 (
            .O(N__8351),
            .I(N__8298));
    ClkMux I__1778 (
            .O(N__8350),
            .I(N__8298));
    ClkMux I__1777 (
            .O(N__8349),
            .I(N__8298));
    ClkMux I__1776 (
            .O(N__8348),
            .I(N__8298));
    ClkMux I__1775 (
            .O(N__8347),
            .I(N__8298));
    ClkMux I__1774 (
            .O(N__8346),
            .I(N__8298));
    ClkMux I__1773 (
            .O(N__8345),
            .I(N__8298));
    ClkMux I__1772 (
            .O(N__8344),
            .I(N__8298));
    ClkMux I__1771 (
            .O(N__8343),
            .I(N__8298));
    ClkMux I__1770 (
            .O(N__8342),
            .I(N__8298));
    Glb2LocalMux I__1769 (
            .O(N__8339),
            .I(N__8298));
    Glb2LocalMux I__1768 (
            .O(N__8336),
            .I(N__8298));
    Glb2LocalMux I__1767 (
            .O(N__8333),
            .I(N__8298));
    Glb2LocalMux I__1766 (
            .O(N__8330),
            .I(N__8298));
    ClkMux I__1765 (
            .O(N__8329),
            .I(N__8298));
    GlobalMux I__1764 (
            .O(N__8298),
            .I(N__8295));
    gio2CtrlBuf I__1763 (
            .O(N__8295),
            .I(CLK40_IN_c_g));
    IoInMux I__1762 (
            .O(N__8292),
            .I(N__8289));
    LocalMux I__1761 (
            .O(N__8289),
            .I(N__8286));
    Span4Mux_s2_v I__1760 (
            .O(N__8286),
            .I(N__8283));
    Span4Mux_v I__1759 (
            .O(N__8283),
            .I(N__8280));
    Odrv4 I__1758 (
            .O(N__8280),
            .I(GB_BUFFER_CLK40_IN_c_g_THRU_CO));
    InMux I__1757 (
            .O(N__8277),
            .I(N__8274));
    LocalMux I__1756 (
            .O(N__8274),
            .I(CIA_ENABLE));
    CascadeMux I__1755 (
            .O(N__8271),
            .I(\U409_TRANSFER_ACK.CIA_STATE_d_2_cascade_ ));
    InMux I__1754 (
            .O(N__8268),
            .I(N__8265));
    LocalMux I__1753 (
            .O(N__8265),
            .I(\U409_TRANSFER_ACK.N_289 ));
    CascadeMux I__1752 (
            .O(N__8262),
            .I(\U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ));
    IoInMux I__1751 (
            .O(N__8259),
            .I(N__8255));
    IoInMux I__1750 (
            .O(N__8258),
            .I(N__8252));
    LocalMux I__1749 (
            .O(N__8255),
            .I(N__8247));
    LocalMux I__1748 (
            .O(N__8252),
            .I(N__8247));
    IoSpan4Mux I__1747 (
            .O(N__8247),
            .I(N__8243));
    IoInMux I__1746 (
            .O(N__8246),
            .I(N__8240));
    Span4Mux_s1_v I__1745 (
            .O(N__8243),
            .I(N__8237));
    LocalMux I__1744 (
            .O(N__8240),
            .I(N__8234));
    Span4Mux_v I__1743 (
            .O(N__8237),
            .I(N__8229));
    Span4Mux_s1_v I__1742 (
            .O(N__8234),
            .I(N__8229));
    Sp12to4 I__1741 (
            .O(N__8229),
            .I(N__8226));
    Span12Mux_h I__1740 (
            .O(N__8226),
            .I(N__8223));
    Span12Mux_v I__1739 (
            .O(N__8223),
            .I(N__8218));
    InMux I__1738 (
            .O(N__8222),
            .I(N__8213));
    InMux I__1737 (
            .O(N__8221),
            .I(N__8213));
    Odrv12 I__1736 (
            .O(N__8218),
            .I(TACK_OUTn));
    LocalMux I__1735 (
            .O(N__8213),
            .I(TACK_OUTn));
    CascadeMux I__1734 (
            .O(N__8208),
            .I(N__8202));
    CascadeMux I__1733 (
            .O(N__8207),
            .I(N__8199));
    CascadeMux I__1732 (
            .O(N__8206),
            .I(N__8196));
    InMux I__1731 (
            .O(N__8205),
            .I(N__8193));
    InMux I__1730 (
            .O(N__8202),
            .I(N__8186));
    InMux I__1729 (
            .O(N__8199),
            .I(N__8186));
    InMux I__1728 (
            .O(N__8196),
            .I(N__8186));
    LocalMux I__1727 (
            .O(N__8193),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    LocalMux I__1726 (
            .O(N__8186),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    InMux I__1725 (
            .O(N__8181),
            .I(N__8175));
    InMux I__1724 (
            .O(N__8180),
            .I(N__8168));
    InMux I__1723 (
            .O(N__8179),
            .I(N__8168));
    InMux I__1722 (
            .O(N__8178),
            .I(N__8168));
    LocalMux I__1721 (
            .O(N__8175),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    LocalMux I__1720 (
            .O(N__8168),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    InMux I__1719 (
            .O(N__8163),
            .I(N__8158));
    InMux I__1718 (
            .O(N__8162),
            .I(N__8153));
    InMux I__1717 (
            .O(N__8161),
            .I(N__8153));
    LocalMux I__1716 (
            .O(N__8158),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    LocalMux I__1715 (
            .O(N__8153),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    InMux I__1714 (
            .O(N__8148),
            .I(N__8145));
    LocalMux I__1713 (
            .O(N__8145),
            .I(N__8141));
    InMux I__1712 (
            .O(N__8144),
            .I(N__8138));
    Odrv4 I__1711 (
            .O(N__8141),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    LocalMux I__1710 (
            .O(N__8138),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    CascadeMux I__1709 (
            .O(N__8133),
            .I(N__8130));
    InMux I__1708 (
            .O(N__8130),
            .I(N__8126));
    CascadeMux I__1707 (
            .O(N__8129),
            .I(N__8123));
    LocalMux I__1706 (
            .O(N__8126),
            .I(N__8120));
    InMux I__1705 (
            .O(N__8123),
            .I(N__8117));
    Span4Mux_h I__1704 (
            .O(N__8120),
            .I(N__8112));
    LocalMux I__1703 (
            .O(N__8117),
            .I(N__8112));
    Span4Mux_h I__1702 (
            .O(N__8112),
            .I(N__8109));
    Odrv4 I__1701 (
            .O(N__8109),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz ));
    InMux I__1700 (
            .O(N__8106),
            .I(N__8102));
    InMux I__1699 (
            .O(N__8105),
            .I(N__8099));
    LocalMux I__1698 (
            .O(N__8102),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    LocalMux I__1697 (
            .O(N__8099),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    CascadeMux I__1696 (
            .O(N__8094),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_ ));
    InMux I__1695 (
            .O(N__8091),
            .I(N__8087));
    InMux I__1694 (
            .O(N__8090),
            .I(N__8084));
    LocalMux I__1693 (
            .O(N__8087),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    LocalMux I__1692 (
            .O(N__8084),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    InMux I__1691 (
            .O(N__8079),
            .I(N__8075));
    InMux I__1690 (
            .O(N__8078),
            .I(N__8072));
    LocalMux I__1689 (
            .O(N__8075),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    LocalMux I__1688 (
            .O(N__8072),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    InMux I__1687 (
            .O(N__8067),
            .I(N__8061));
    InMux I__1686 (
            .O(N__8066),
            .I(N__8061));
    LocalMux I__1685 (
            .O(N__8061),
            .I(\U409_TRANSFER_ACK.N_159 ));
    InMux I__1684 (
            .O(N__8058),
            .I(N__8055));
    LocalMux I__1683 (
            .O(N__8055),
            .I(\U409_TRANSFER_ACK.N_380 ));
    CascadeMux I__1682 (
            .O(N__8052),
            .I(\U409_TRANSFER_ACK.N_380_cascade_ ));
    InMux I__1681 (
            .O(N__8049),
            .I(N__8046));
    LocalMux I__1680 (
            .O(N__8046),
            .I(N_190));
    InMux I__1679 (
            .O(N__8043),
            .I(N__8040));
    LocalMux I__1678 (
            .O(N__8040),
            .I(N__8036));
    InMux I__1677 (
            .O(N__8039),
            .I(N__8033));
    Span4Mux_v I__1676 (
            .O(N__8036),
            .I(N__8030));
    LocalMux I__1675 (
            .O(N__8033),
            .I(N__8027));
    Odrv4 I__1674 (
            .O(N__8030),
            .I(N_297));
    Odrv4 I__1673 (
            .O(N__8027),
            .I(N_297));
    IoInMux I__1672 (
            .O(N__8022),
            .I(N__8019));
    LocalMux I__1671 (
            .O(N__8019),
            .I(N__8016));
    Span12Mux_s7_v I__1670 (
            .O(N__8016),
            .I(N__8013));
    Span12Mux_h I__1669 (
            .O(N__8013),
            .I(N__8010));
    Odrv12 I__1668 (
            .O(N__8010),
            .I(N_94_i));
    InMux I__1667 (
            .O(N__8007),
            .I(N__8004));
    LocalMux I__1666 (
            .O(N__8004),
            .I(N__8001));
    Span4Mux_v I__1665 (
            .O(N__8001),
            .I(N__7998));
    Sp12to4 I__1664 (
            .O(N__7998),
            .I(N__7995));
    Span12Mux_h I__1663 (
            .O(N__7995),
            .I(N__7992));
    Odrv12 I__1662 (
            .O(N__7992),
            .I(A_c_13));
    IoInMux I__1661 (
            .O(N__7989),
            .I(N__7986));
    LocalMux I__1660 (
            .O(N__7986),
            .I(N__7983));
    Span4Mux_s1_h I__1659 (
            .O(N__7983),
            .I(N__7980));
    Sp12to4 I__1658 (
            .O(N__7980),
            .I(N__7977));
    Span12Mux_s9_v I__1657 (
            .O(N__7977),
            .I(N__7974));
    Span12Mux_h I__1656 (
            .O(N__7974),
            .I(N__7971));
    Odrv12 I__1655 (
            .O(N__7971),
            .I(U409_ADDRESS_DECODE_un1_CIACS1n_i));
    InMux I__1654 (
            .O(N__7968),
            .I(N__7965));
    LocalMux I__1653 (
            .O(N__7965),
            .I(N__7959));
    InMux I__1652 (
            .O(N__7964),
            .I(N__7956));
    InMux I__1651 (
            .O(N__7963),
            .I(N__7953));
    InMux I__1650 (
            .O(N__7962),
            .I(N__7949));
    Span4Mux_v I__1649 (
            .O(N__7959),
            .I(N__7944));
    LocalMux I__1648 (
            .O(N__7956),
            .I(N__7944));
    LocalMux I__1647 (
            .O(N__7953),
            .I(N__7941));
    InMux I__1646 (
            .O(N__7952),
            .I(N__7938));
    LocalMux I__1645 (
            .O(N__7949),
            .I(N__7933));
    Span4Mux_v I__1644 (
            .O(N__7944),
            .I(N__7926));
    Span4Mux_h I__1643 (
            .O(N__7941),
            .I(N__7926));
    LocalMux I__1642 (
            .O(N__7938),
            .I(N__7926));
    InMux I__1641 (
            .O(N__7937),
            .I(N__7923));
    InMux I__1640 (
            .O(N__7936),
            .I(N__7920));
    Span4Mux_v I__1639 (
            .O(N__7933),
            .I(N__7917));
    Span4Mux_h I__1638 (
            .O(N__7926),
            .I(N__7912));
    LocalMux I__1637 (
            .O(N__7923),
            .I(N__7912));
    LocalMux I__1636 (
            .O(N__7920),
            .I(N__7909));
    Span4Mux_v I__1635 (
            .O(N__7917),
            .I(N__7906));
    Span4Mux_v I__1634 (
            .O(N__7912),
            .I(N__7903));
    Span12Mux_h I__1633 (
            .O(N__7909),
            .I(N__7900));
    Span4Mux_v I__1632 (
            .O(N__7906),
            .I(N__7897));
    Span4Mux_v I__1631 (
            .O(N__7903),
            .I(N__7894));
    Span12Mux_v I__1630 (
            .O(N__7900),
            .I(N__7891));
    Sp12to4 I__1629 (
            .O(N__7897),
            .I(N__7886));
    Sp12to4 I__1628 (
            .O(N__7894),
            .I(N__7886));
    Odrv12 I__1627 (
            .O(N__7891),
            .I(A_c_22));
    Odrv12 I__1626 (
            .O(N__7886),
            .I(A_c_22));
    CascadeMux I__1625 (
            .O(N__7881),
            .I(N__7878));
    InMux I__1624 (
            .O(N__7878),
            .I(N__7875));
    LocalMux I__1623 (
            .O(N__7875),
            .I(N__7871));
    CascadeMux I__1622 (
            .O(N__7874),
            .I(N__7867));
    Span4Mux_v I__1621 (
            .O(N__7871),
            .I(N__7864));
    InMux I__1620 (
            .O(N__7870),
            .I(N__7861));
    InMux I__1619 (
            .O(N__7867),
            .I(N__7858));
    Sp12to4 I__1618 (
            .O(N__7864),
            .I(N__7850));
    LocalMux I__1617 (
            .O(N__7861),
            .I(N__7850));
    LocalMux I__1616 (
            .O(N__7858),
            .I(N__7850));
    InMux I__1615 (
            .O(N__7857),
            .I(N__7847));
    Odrv12 I__1614 (
            .O(N__7850),
            .I(N_401));
    LocalMux I__1613 (
            .O(N__7847),
            .I(N_401));
    CascadeMux I__1612 (
            .O(N__7842),
            .I(N_431_cascade_));
    InMux I__1611 (
            .O(N__7839),
            .I(N__7836));
    LocalMux I__1610 (
            .O(N__7836),
            .I(N__7832));
    InMux I__1609 (
            .O(N__7835),
            .I(N__7829));
    Span4Mux_h I__1608 (
            .O(N__7832),
            .I(N__7823));
    LocalMux I__1607 (
            .O(N__7829),
            .I(N__7823));
    InMux I__1606 (
            .O(N__7828),
            .I(N__7820));
    Sp12to4 I__1605 (
            .O(N__7823),
            .I(N__7815));
    LocalMux I__1604 (
            .O(N__7820),
            .I(N__7815));
    Odrv12 I__1603 (
            .O(N__7815),
            .I(N_422));
    InMux I__1602 (
            .O(N__7812),
            .I(N__7808));
    InMux I__1601 (
            .O(N__7811),
            .I(N__7805));
    LocalMux I__1600 (
            .O(N__7808),
            .I(N__7797));
    LocalMux I__1599 (
            .O(N__7805),
            .I(N__7797));
    InMux I__1598 (
            .O(N__7804),
            .I(N__7794));
    InMux I__1597 (
            .O(N__7803),
            .I(N__7791));
    InMux I__1596 (
            .O(N__7802),
            .I(N__7788));
    Span4Mux_v I__1595 (
            .O(N__7797),
            .I(N__7784));
    LocalMux I__1594 (
            .O(N__7794),
            .I(N__7781));
    LocalMux I__1593 (
            .O(N__7791),
            .I(N__7778));
    LocalMux I__1592 (
            .O(N__7788),
            .I(N__7775));
    InMux I__1591 (
            .O(N__7787),
            .I(N__7772));
    Span4Mux_h I__1590 (
            .O(N__7784),
            .I(N__7767));
    Span4Mux_v I__1589 (
            .O(N__7781),
            .I(N__7767));
    Span4Mux_v I__1588 (
            .O(N__7778),
            .I(N__7764));
    Span4Mux_v I__1587 (
            .O(N__7775),
            .I(N__7759));
    LocalMux I__1586 (
            .O(N__7772),
            .I(N__7759));
    Span4Mux_v I__1585 (
            .O(N__7767),
            .I(N__7756));
    Span4Mux_h I__1584 (
            .O(N__7764),
            .I(N__7751));
    Span4Mux_v I__1583 (
            .O(N__7759),
            .I(N__7751));
    Sp12to4 I__1582 (
            .O(N__7756),
            .I(N__7746));
    Sp12to4 I__1581 (
            .O(N__7751),
            .I(N__7746));
    Span12Mux_h I__1580 (
            .O(N__7746),
            .I(N__7743));
    Span12Mux_v I__1579 (
            .O(N__7743),
            .I(N__7740));
    Odrv12 I__1578 (
            .O(N__7740),
            .I(A_c_19));
    InMux I__1577 (
            .O(N__7737),
            .I(N__7733));
    InMux I__1576 (
            .O(N__7736),
            .I(N__7730));
    LocalMux I__1575 (
            .O(N__7733),
            .I(ATA_BASE_7));
    LocalMux I__1574 (
            .O(N__7730),
            .I(ATA_BASE_7));
    CascadeMux I__1573 (
            .O(N__7725),
            .I(N__7722));
    InMux I__1572 (
            .O(N__7722),
            .I(N__7719));
    LocalMux I__1571 (
            .O(N__7719),
            .I(N__7715));
    InMux I__1570 (
            .O(N__7718),
            .I(N__7712));
    Span4Mux_v I__1569 (
            .O(N__7715),
            .I(N__7708));
    LocalMux I__1568 (
            .O(N__7712),
            .I(N__7705));
    InMux I__1567 (
            .O(N__7711),
            .I(N__7702));
    Span4Mux_v I__1566 (
            .O(N__7708),
            .I(N__7696));
    Span4Mux_h I__1565 (
            .O(N__7705),
            .I(N__7691));
    LocalMux I__1564 (
            .O(N__7702),
            .I(N__7691));
    InMux I__1563 (
            .O(N__7701),
            .I(N__7688));
    CascadeMux I__1562 (
            .O(N__7700),
            .I(N__7685));
    CascadeMux I__1561 (
            .O(N__7699),
            .I(N__7682));
    Span4Mux_h I__1560 (
            .O(N__7696),
            .I(N__7679));
    Span4Mux_v I__1559 (
            .O(N__7691),
            .I(N__7676));
    LocalMux I__1558 (
            .O(N__7688),
            .I(N__7673));
    InMux I__1557 (
            .O(N__7685),
            .I(N__7668));
    InMux I__1556 (
            .O(N__7682),
            .I(N__7668));
    Sp12to4 I__1555 (
            .O(N__7679),
            .I(N__7659));
    Sp12to4 I__1554 (
            .O(N__7676),
            .I(N__7659));
    Span12Mux_h I__1553 (
            .O(N__7673),
            .I(N__7659));
    LocalMux I__1552 (
            .O(N__7668),
            .I(N__7659));
    Odrv12 I__1551 (
            .O(N__7659),
            .I(A_c_23));
    InMux I__1550 (
            .O(N__7656),
            .I(N__7650));
    InMux I__1549 (
            .O(N__7655),
            .I(N__7650));
    LocalMux I__1548 (
            .O(N__7650),
            .I(\U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_5 ));
    CascadeMux I__1547 (
            .O(N__7647),
            .I(N__7640));
    InMux I__1546 (
            .O(N__7646),
            .I(N__7629));
    InMux I__1545 (
            .O(N__7645),
            .I(N__7629));
    InMux I__1544 (
            .O(N__7644),
            .I(N__7629));
    InMux I__1543 (
            .O(N__7643),
            .I(N__7629));
    InMux I__1542 (
            .O(N__7640),
            .I(N__7626));
    CascadeMux I__1541 (
            .O(N__7639),
            .I(N__7620));
    CascadeMux I__1540 (
            .O(N__7638),
            .I(N__7615));
    LocalMux I__1539 (
            .O(N__7629),
            .I(N__7612));
    LocalMux I__1538 (
            .O(N__7626),
            .I(N__7609));
    InMux I__1537 (
            .O(N__7625),
            .I(N__7594));
    InMux I__1536 (
            .O(N__7624),
            .I(N__7594));
    InMux I__1535 (
            .O(N__7623),
            .I(N__7594));
    InMux I__1534 (
            .O(N__7620),
            .I(N__7594));
    InMux I__1533 (
            .O(N__7619),
            .I(N__7594));
    InMux I__1532 (
            .O(N__7618),
            .I(N__7594));
    InMux I__1531 (
            .O(N__7615),
            .I(N__7594));
    Span4Mux_v I__1530 (
            .O(N__7612),
            .I(N__7591));
    Span4Mux_v I__1529 (
            .O(N__7609),
            .I(N__7588));
    LocalMux I__1528 (
            .O(N__7594),
            .I(N__7585));
    Odrv4 I__1527 (
            .O(N__7591),
            .I(N_361));
    Odrv4 I__1526 (
            .O(N__7588),
            .I(N_361));
    Odrv12 I__1525 (
            .O(N__7585),
            .I(N_361));
    CascadeMux I__1524 (
            .O(N__7578),
            .I(N__7574));
    CascadeMux I__1523 (
            .O(N__7577),
            .I(N__7571));
    InMux I__1522 (
            .O(N__7574),
            .I(N__7568));
    InMux I__1521 (
            .O(N__7571),
            .I(N__7565));
    LocalMux I__1520 (
            .O(N__7568),
            .I(N__7562));
    LocalMux I__1519 (
            .O(N__7565),
            .I(N__7559));
    Span4Mux_v I__1518 (
            .O(N__7562),
            .I(N__7555));
    Span4Mux_v I__1517 (
            .O(N__7559),
            .I(N__7552));
    InMux I__1516 (
            .O(N__7558),
            .I(N__7549));
    Span4Mux_h I__1515 (
            .O(N__7555),
            .I(N__7546));
    Span4Mux_v I__1514 (
            .O(N__7552),
            .I(N__7543));
    LocalMux I__1513 (
            .O(N__7549),
            .I(N__7540));
    Sp12to4 I__1512 (
            .O(N__7546),
            .I(N__7535));
    Sp12to4 I__1511 (
            .O(N__7543),
            .I(N__7535));
    Span4Mux_v I__1510 (
            .O(N__7540),
            .I(N__7532));
    Span12Mux_h I__1509 (
            .O(N__7535),
            .I(N__7527));
    Sp12to4 I__1508 (
            .O(N__7532),
            .I(N__7527));
    Odrv12 I__1507 (
            .O(N__7527),
            .I(D_in_7));
    InMux I__1506 (
            .O(N__7524),
            .I(N__7518));
    InMux I__1505 (
            .O(N__7523),
            .I(N__7518));
    LocalMux I__1504 (
            .O(N__7518),
            .I(ATA_BASE_3));
    CEMux I__1503 (
            .O(N__7515),
            .I(N__7512));
    LocalMux I__1502 (
            .O(N__7512),
            .I(N__7509));
    Span4Mux_h I__1501 (
            .O(N__7509),
            .I(N__7506));
    Span4Mux_h I__1500 (
            .O(N__7506),
            .I(N__7502));
    CEMux I__1499 (
            .O(N__7505),
            .I(N__7499));
    Odrv4 I__1498 (
            .O(N__7502),
            .I(\U409_AUTOCONFIG.un1_STATE_1_0_0 ));
    LocalMux I__1497 (
            .O(N__7499),
            .I(\U409_AUTOCONFIG.un1_STATE_1_0_0 ));
    InMux I__1496 (
            .O(N__7494),
            .I(N__7482));
    InMux I__1495 (
            .O(N__7493),
            .I(N__7482));
    InMux I__1494 (
            .O(N__7492),
            .I(N__7482));
    InMux I__1493 (
            .O(N__7491),
            .I(N__7482));
    LocalMux I__1492 (
            .O(N__7482),
            .I(\U409_AUTOCONFIG.N_172 ));
    CascadeMux I__1491 (
            .O(N__7479),
            .I(N__7476));
    InMux I__1490 (
            .O(N__7476),
            .I(N__7472));
    InMux I__1489 (
            .O(N__7475),
            .I(N__7465));
    LocalMux I__1488 (
            .O(N__7472),
            .I(N__7461));
    InMux I__1487 (
            .O(N__7471),
            .I(N__7458));
    InMux I__1486 (
            .O(N__7470),
            .I(N__7455));
    CascadeMux I__1485 (
            .O(N__7469),
            .I(N__7452));
    InMux I__1484 (
            .O(N__7468),
            .I(N__7447));
    LocalMux I__1483 (
            .O(N__7465),
            .I(N__7444));
    CascadeMux I__1482 (
            .O(N__7464),
            .I(N__7440));
    Span4Mux_h I__1481 (
            .O(N__7461),
            .I(N__7435));
    LocalMux I__1480 (
            .O(N__7458),
            .I(N__7435));
    LocalMux I__1479 (
            .O(N__7455),
            .I(N__7432));
    InMux I__1478 (
            .O(N__7452),
            .I(N__7429));
    InMux I__1477 (
            .O(N__7451),
            .I(N__7424));
    InMux I__1476 (
            .O(N__7450),
            .I(N__7424));
    LocalMux I__1475 (
            .O(N__7447),
            .I(N__7421));
    Span4Mux_h I__1474 (
            .O(N__7444),
            .I(N__7418));
    InMux I__1473 (
            .O(N__7443),
            .I(N__7413));
    InMux I__1472 (
            .O(N__7440),
            .I(N__7413));
    Odrv4 I__1471 (
            .O(N__7435),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    Odrv12 I__1470 (
            .O(N__7432),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    LocalMux I__1469 (
            .O(N__7429),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    LocalMux I__1468 (
            .O(N__7424),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    Odrv12 I__1467 (
            .O(N__7421),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    Odrv4 I__1466 (
            .O(N__7418),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    LocalMux I__1465 (
            .O(N__7413),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    InMux I__1464 (
            .O(N__7398),
            .I(N__7395));
    LocalMux I__1463 (
            .O(N__7395),
            .I(N__7388));
    InMux I__1462 (
            .O(N__7394),
            .I(N__7383));
    InMux I__1461 (
            .O(N__7393),
            .I(N__7383));
    InMux I__1460 (
            .O(N__7392),
            .I(N__7378));
    InMux I__1459 (
            .O(N__7391),
            .I(N__7378));
    Odrv4 I__1458 (
            .O(N__7388),
            .I(\U409_AUTOCONFIG.un1_STATE_1_0_a2_0 ));
    LocalMux I__1457 (
            .O(N__7383),
            .I(\U409_AUTOCONFIG.un1_STATE_1_0_a2_0 ));
    LocalMux I__1456 (
            .O(N__7378),
            .I(\U409_AUTOCONFIG.un1_STATE_1_0_a2_0 ));
    InMux I__1455 (
            .O(N__7371),
            .I(N__7357));
    InMux I__1454 (
            .O(N__7370),
            .I(N__7357));
    InMux I__1453 (
            .O(N__7369),
            .I(N__7350));
    InMux I__1452 (
            .O(N__7368),
            .I(N__7350));
    InMux I__1451 (
            .O(N__7367),
            .I(N__7350));
    CascadeMux I__1450 (
            .O(N__7366),
            .I(N__7347));
    CascadeMux I__1449 (
            .O(N__7365),
            .I(N__7343));
    CascadeMux I__1448 (
            .O(N__7364),
            .I(N__7340));
    CascadeMux I__1447 (
            .O(N__7363),
            .I(N__7337));
    CascadeMux I__1446 (
            .O(N__7362),
            .I(N__7334));
    LocalMux I__1445 (
            .O(N__7357),
            .I(N__7320));
    LocalMux I__1444 (
            .O(N__7350),
            .I(N__7320));
    InMux I__1443 (
            .O(N__7347),
            .I(N__7317));
    InMux I__1442 (
            .O(N__7346),
            .I(N__7312));
    InMux I__1441 (
            .O(N__7343),
            .I(N__7312));
    InMux I__1440 (
            .O(N__7340),
            .I(N__7305));
    InMux I__1439 (
            .O(N__7337),
            .I(N__7305));
    InMux I__1438 (
            .O(N__7334),
            .I(N__7305));
    InMux I__1437 (
            .O(N__7333),
            .I(N__7294));
    InMux I__1436 (
            .O(N__7332),
            .I(N__7294));
    InMux I__1435 (
            .O(N__7331),
            .I(N__7294));
    InMux I__1434 (
            .O(N__7330),
            .I(N__7294));
    InMux I__1433 (
            .O(N__7329),
            .I(N__7294));
    InMux I__1432 (
            .O(N__7328),
            .I(N__7291));
    InMux I__1431 (
            .O(N__7327),
            .I(N__7286));
    InMux I__1430 (
            .O(N__7326),
            .I(N__7286));
    CascadeMux I__1429 (
            .O(N__7325),
            .I(N__7281));
    Span4Mux_v I__1428 (
            .O(N__7320),
            .I(N__7275));
    LocalMux I__1427 (
            .O(N__7317),
            .I(N__7275));
    LocalMux I__1426 (
            .O(N__7312),
            .I(N__7272));
    LocalMux I__1425 (
            .O(N__7305),
            .I(N__7263));
    LocalMux I__1424 (
            .O(N__7294),
            .I(N__7263));
    LocalMux I__1423 (
            .O(N__7291),
            .I(N__7263));
    LocalMux I__1422 (
            .O(N__7286),
            .I(N__7263));
    InMux I__1421 (
            .O(N__7285),
            .I(N__7258));
    InMux I__1420 (
            .O(N__7284),
            .I(N__7258));
    InMux I__1419 (
            .O(N__7281),
            .I(N__7255));
    InMux I__1418 (
            .O(N__7280),
            .I(N__7252));
    Span4Mux_v I__1417 (
            .O(N__7275),
            .I(N__7249));
    Span4Mux_v I__1416 (
            .O(N__7272),
            .I(N__7246));
    Span4Mux_v I__1415 (
            .O(N__7263),
            .I(N__7243));
    LocalMux I__1414 (
            .O(N__7258),
            .I(N__7236));
    LocalMux I__1413 (
            .O(N__7255),
            .I(N__7236));
    LocalMux I__1412 (
            .O(N__7252),
            .I(N__7236));
    Sp12to4 I__1411 (
            .O(N__7249),
            .I(N__7229));
    Sp12to4 I__1410 (
            .O(N__7246),
            .I(N__7229));
    Sp12to4 I__1409 (
            .O(N__7243),
            .I(N__7229));
    Span12Mux_h I__1408 (
            .O(N__7236),
            .I(N__7226));
    Span12Mux_h I__1407 (
            .O(N__7229),
            .I(N__7223));
    Span12Mux_v I__1406 (
            .O(N__7226),
            .I(N__7220));
    Span12Mux_v I__1405 (
            .O(N__7223),
            .I(N__7217));
    Odrv12 I__1404 (
            .O(N__7220),
            .I(A_c_1));
    Odrv12 I__1403 (
            .O(N__7217),
            .I(A_c_1));
    IoInMux I__1402 (
            .O(N__7212),
            .I(N__7209));
    LocalMux I__1401 (
            .O(N__7209),
            .I(N__7206));
    Span4Mux_s3_v I__1400 (
            .O(N__7206),
            .I(N__7203));
    Sp12to4 I__1399 (
            .O(N__7203),
            .I(N__7198));
    InMux I__1398 (
            .O(N__7202),
            .I(N__7195));
    InMux I__1397 (
            .O(N__7201),
            .I(N__7192));
    Span12Mux_h I__1396 (
            .O(N__7198),
            .I(N__7189));
    LocalMux I__1395 (
            .O(N__7195),
            .I(N__7183));
    LocalMux I__1394 (
            .O(N__7192),
            .I(N__7183));
    Span12Mux_v I__1393 (
            .O(N__7189),
            .I(N__7179));
    InMux I__1392 (
            .O(N__7188),
            .I(N__7176));
    Span4Mux_h I__1391 (
            .O(N__7183),
            .I(N__7173));
    InMux I__1390 (
            .O(N__7182),
            .I(N__7170));
    Odrv12 I__1389 (
            .O(N__7179),
            .I(CONFIGENn_c));
    LocalMux I__1388 (
            .O(N__7176),
            .I(CONFIGENn_c));
    Odrv4 I__1387 (
            .O(N__7173),
            .I(CONFIGENn_c));
    LocalMux I__1386 (
            .O(N__7170),
            .I(CONFIGENn_c));
    InMux I__1385 (
            .O(N__7161),
            .I(N__7157));
    InMux I__1384 (
            .O(N__7160),
            .I(N__7154));
    LocalMux I__1383 (
            .O(N__7157),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    LocalMux I__1382 (
            .O(N__7154),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    InMux I__1381 (
            .O(N__7149),
            .I(N__7146));
    LocalMux I__1380 (
            .O(N__7146),
            .I(N__7143));
    Odrv4 I__1379 (
            .O(N__7143),
            .I(AC_TACK));
    InMux I__1378 (
            .O(N__7140),
            .I(N__7136));
    InMux I__1377 (
            .O(N__7139),
            .I(N__7131));
    LocalMux I__1376 (
            .O(N__7136),
            .I(N__7128));
    InMux I__1375 (
            .O(N__7135),
            .I(N__7125));
    CascadeMux I__1374 (
            .O(N__7134),
            .I(N__7122));
    LocalMux I__1373 (
            .O(N__7131),
            .I(N__7118));
    Span4Mux_v I__1372 (
            .O(N__7128),
            .I(N__7113));
    LocalMux I__1371 (
            .O(N__7125),
            .I(N__7113));
    InMux I__1370 (
            .O(N__7122),
            .I(N__7110));
    InMux I__1369 (
            .O(N__7121),
            .I(N__7107));
    Span4Mux_v I__1368 (
            .O(N__7118),
            .I(N__7104));
    Span4Mux_h I__1367 (
            .O(N__7113),
            .I(N__7101));
    LocalMux I__1366 (
            .O(N__7110),
            .I(N__7094));
    LocalMux I__1365 (
            .O(N__7107),
            .I(N__7094));
    Sp12to4 I__1364 (
            .O(N__7104),
            .I(N__7094));
    Span4Mux_h I__1363 (
            .O(N__7101),
            .I(N__7091));
    Span12Mux_h I__1362 (
            .O(N__7094),
            .I(N__7088));
    Sp12to4 I__1361 (
            .O(N__7091),
            .I(N__7085));
    Span12Mux_v I__1360 (
            .O(N__7088),
            .I(N__7082));
    Span12Mux_v I__1359 (
            .O(N__7085),
            .I(N__7079));
    Odrv12 I__1358 (
            .O(N__7082),
            .I(RnW_c));
    Odrv12 I__1357 (
            .O(N__7079),
            .I(RnW_c));
    CascadeMux I__1356 (
            .O(N__7074),
            .I(N__7071));
    InMux I__1355 (
            .O(N__7071),
            .I(N__7068));
    LocalMux I__1354 (
            .O(N__7068),
            .I(N__7064));
    InMux I__1353 (
            .O(N__7067),
            .I(N__7061));
    Span4Mux_v I__1352 (
            .O(N__7064),
            .I(N__7056));
    LocalMux I__1351 (
            .O(N__7061),
            .I(N__7053));
    InMux I__1350 (
            .O(N__7060),
            .I(N__7048));
    InMux I__1349 (
            .O(N__7059),
            .I(N__7048));
    Odrv4 I__1348 (
            .O(N__7056),
            .I(N_356));
    Odrv4 I__1347 (
            .O(N__7053),
            .I(N_356));
    LocalMux I__1346 (
            .O(N__7048),
            .I(N_356));
    InMux I__1345 (
            .O(N__7041),
            .I(N__7032));
    InMux I__1344 (
            .O(N__7040),
            .I(N__7027));
    InMux I__1343 (
            .O(N__7039),
            .I(N__7027));
    InMux I__1342 (
            .O(N__7038),
            .I(N__7024));
    InMux I__1341 (
            .O(N__7037),
            .I(N__7017));
    InMux I__1340 (
            .O(N__7036),
            .I(N__7017));
    InMux I__1339 (
            .O(N__7035),
            .I(N__7017));
    LocalMux I__1338 (
            .O(N__7032),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1337 (
            .O(N__7027),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1336 (
            .O(N__7024),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1335 (
            .O(N__7017),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    InMux I__1334 (
            .O(N__7008),
            .I(N__7002));
    InMux I__1333 (
            .O(N__7007),
            .I(N__6999));
    InMux I__1332 (
            .O(N__7006),
            .I(N__6994));
    InMux I__1331 (
            .O(N__7005),
            .I(N__6994));
    LocalMux I__1330 (
            .O(N__7002),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1329 (
            .O(N__6999),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1328 (
            .O(N__6994),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    InMux I__1327 (
            .O(N__6987),
            .I(N__6980));
    InMux I__1326 (
            .O(N__6986),
            .I(N__6977));
    InMux I__1325 (
            .O(N__6985),
            .I(N__6974));
    InMux I__1324 (
            .O(N__6984),
            .I(N__6971));
    InMux I__1323 (
            .O(N__6983),
            .I(N__6968));
    LocalMux I__1322 (
            .O(N__6980),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1321 (
            .O(N__6977),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1320 (
            .O(N__6974),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1319 (
            .O(N__6971),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1318 (
            .O(N__6968),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    CascadeMux I__1317 (
            .O(N__6957),
            .I(N__6953));
    InMux I__1316 (
            .O(N__6956),
            .I(N__6949));
    InMux I__1315 (
            .O(N__6953),
            .I(N__6944));
    InMux I__1314 (
            .O(N__6952),
            .I(N__6944));
    LocalMux I__1313 (
            .O(N__6949),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ));
    LocalMux I__1312 (
            .O(N__6944),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ));
    CascadeMux I__1311 (
            .O(N__6939),
            .I(N__6936));
    InMux I__1310 (
            .O(N__6936),
            .I(N__6933));
    LocalMux I__1309 (
            .O(N__6933),
            .I(N__6928));
    InMux I__1308 (
            .O(N__6932),
            .I(N__6925));
    CascadeMux I__1307 (
            .O(N__6931),
            .I(N__6922));
    Span4Mux_h I__1306 (
            .O(N__6928),
            .I(N__6915));
    LocalMux I__1305 (
            .O(N__6925),
            .I(N__6915));
    InMux I__1304 (
            .O(N__6922),
            .I(N__6912));
    InMux I__1303 (
            .O(N__6921),
            .I(N__6906));
    InMux I__1302 (
            .O(N__6920),
            .I(N__6906));
    Span4Mux_v I__1301 (
            .O(N__6915),
            .I(N__6901));
    LocalMux I__1300 (
            .O(N__6912),
            .I(N__6901));
    CascadeMux I__1299 (
            .O(N__6911),
            .I(N__6897));
    LocalMux I__1298 (
            .O(N__6906),
            .I(N__6894));
    Span4Mux_v I__1297 (
            .O(N__6901),
            .I(N__6890));
    InMux I__1296 (
            .O(N__6900),
            .I(N__6887));
    InMux I__1295 (
            .O(N__6897),
            .I(N__6884));
    Span4Mux_v I__1294 (
            .O(N__6894),
            .I(N__6881));
    InMux I__1293 (
            .O(N__6893),
            .I(N__6878));
    Sp12to4 I__1292 (
            .O(N__6890),
            .I(N__6867));
    LocalMux I__1291 (
            .O(N__6887),
            .I(N__6867));
    LocalMux I__1290 (
            .O(N__6884),
            .I(N__6867));
    Sp12to4 I__1289 (
            .O(N__6881),
            .I(N__6867));
    LocalMux I__1288 (
            .O(N__6878),
            .I(N__6867));
    Span12Mux_h I__1287 (
            .O(N__6867),
            .I(N__6864));
    Odrv12 I__1286 (
            .O(N__6864),
            .I(A_c_20));
    CascadeMux I__1285 (
            .O(N__6861),
            .I(\U409_TRANSFER_ACK.N_346_cascade_ ));
    InMux I__1284 (
            .O(N__6858),
            .I(N__6855));
    LocalMux I__1283 (
            .O(N__6855),
            .I(N__6851));
    InMux I__1282 (
            .O(N__6854),
            .I(N__6848));
    Span4Mux_v I__1281 (
            .O(N__6851),
            .I(N__6843));
    LocalMux I__1280 (
            .O(N__6848),
            .I(N__6843));
    Span4Mux_h I__1279 (
            .O(N__6843),
            .I(N__6839));
    InMux I__1278 (
            .O(N__6842),
            .I(N__6836));
    Odrv4 I__1277 (
            .O(N__6839),
            .I(N_434));
    LocalMux I__1276 (
            .O(N__6836),
            .I(N_434));
    CascadeMux I__1275 (
            .O(N__6831),
            .I(N_190_cascade_));
    InMux I__1274 (
            .O(N__6828),
            .I(N__6825));
    LocalMux I__1273 (
            .O(N__6825),
            .I(N__6822));
    Span12Mux_h I__1272 (
            .O(N__6822),
            .I(N__6819));
    Span12Mux_h I__1271 (
            .O(N__6819),
            .I(N__6816));
    Span12Mux_v I__1270 (
            .O(N__6816),
            .I(N__6813));
    Odrv12 I__1269 (
            .O(N__6813),
            .I(TACKn_in));
    SRMux I__1268 (
            .O(N__6810),
            .I(N__6805));
    SRMux I__1267 (
            .O(N__6809),
            .I(N__6802));
    SRMux I__1266 (
            .O(N__6808),
            .I(N__6799));
    LocalMux I__1265 (
            .O(N__6805),
            .I(N__6792));
    LocalMux I__1264 (
            .O(N__6802),
            .I(N__6792));
    LocalMux I__1263 (
            .O(N__6799),
            .I(N__6792));
    Span4Mux_v I__1262 (
            .O(N__6792),
            .I(N__6789));
    Span4Mux_v I__1261 (
            .O(N__6789),
            .I(N__6786));
    Odrv4 I__1260 (
            .O(N__6786),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    InMux I__1259 (
            .O(N__6783),
            .I(N__6779));
    InMux I__1258 (
            .O(N__6782),
            .I(N__6776));
    LocalMux I__1257 (
            .O(N__6779),
            .I(N__6771));
    LocalMux I__1256 (
            .O(N__6776),
            .I(N__6768));
    InMux I__1255 (
            .O(N__6775),
            .I(N__6765));
    InMux I__1254 (
            .O(N__6774),
            .I(N__6760));
    Span4Mux_v I__1253 (
            .O(N__6771),
            .I(N__6753));
    Span4Mux_h I__1252 (
            .O(N__6768),
            .I(N__6753));
    LocalMux I__1251 (
            .O(N__6765),
            .I(N__6753));
    InMux I__1250 (
            .O(N__6764),
            .I(N__6750));
    InMux I__1249 (
            .O(N__6763),
            .I(N__6747));
    LocalMux I__1248 (
            .O(N__6760),
            .I(N__6738));
    Span4Mux_h I__1247 (
            .O(N__6753),
            .I(N__6738));
    LocalMux I__1246 (
            .O(N__6750),
            .I(N__6738));
    LocalMux I__1245 (
            .O(N__6747),
            .I(N__6738));
    Span4Mux_v I__1244 (
            .O(N__6738),
            .I(N__6732));
    InMux I__1243 (
            .O(N__6737),
            .I(N__6727));
    InMux I__1242 (
            .O(N__6736),
            .I(N__6727));
    InMux I__1241 (
            .O(N__6735),
            .I(N__6724));
    Sp12to4 I__1240 (
            .O(N__6732),
            .I(N__6717));
    LocalMux I__1239 (
            .O(N__6727),
            .I(N__6717));
    LocalMux I__1238 (
            .O(N__6724),
            .I(N__6714));
    InMux I__1237 (
            .O(N__6723),
            .I(N__6709));
    InMux I__1236 (
            .O(N__6722),
            .I(N__6709));
    Span12Mux_h I__1235 (
            .O(N__6717),
            .I(N__6702));
    Sp12to4 I__1234 (
            .O(N__6714),
            .I(N__6702));
    LocalMux I__1233 (
            .O(N__6709),
            .I(N__6702));
    Odrv12 I__1232 (
            .O(N__6702),
            .I(A_c_21));
    InMux I__1231 (
            .O(N__6699),
            .I(N__6689));
    InMux I__1230 (
            .O(N__6698),
            .I(N__6689));
    InMux I__1229 (
            .O(N__6697),
            .I(N__6686));
    InMux I__1228 (
            .O(N__6696),
            .I(N__6683));
    InMux I__1227 (
            .O(N__6695),
            .I(N__6680));
    CascadeMux I__1226 (
            .O(N__6694),
            .I(N__6677));
    LocalMux I__1225 (
            .O(N__6689),
            .I(N__6674));
    LocalMux I__1224 (
            .O(N__6686),
            .I(N__6671));
    LocalMux I__1223 (
            .O(N__6683),
            .I(N__6666));
    LocalMux I__1222 (
            .O(N__6680),
            .I(N__6666));
    InMux I__1221 (
            .O(N__6677),
            .I(N__6663));
    Span4Mux_v I__1220 (
            .O(N__6674),
            .I(N__6654));
    Span4Mux_v I__1219 (
            .O(N__6671),
            .I(N__6654));
    Span4Mux_v I__1218 (
            .O(N__6666),
            .I(N__6654));
    LocalMux I__1217 (
            .O(N__6663),
            .I(N__6651));
    InMux I__1216 (
            .O(N__6662),
            .I(N__6646));
    InMux I__1215 (
            .O(N__6661),
            .I(N__6646));
    Odrv4 I__1214 (
            .O(N__6654),
            .I(N_351));
    Odrv12 I__1213 (
            .O(N__6651),
            .I(N_351));
    LocalMux I__1212 (
            .O(N__6646),
            .I(N_351));
    IoInMux I__1211 (
            .O(N__6639),
            .I(N__6636));
    LocalMux I__1210 (
            .O(N__6636),
            .I(N__6633));
    IoSpan4Mux I__1209 (
            .O(N__6633),
            .I(N__6630));
    Sp12to4 I__1208 (
            .O(N__6630),
            .I(N__6627));
    Span12Mux_s7_h I__1207 (
            .O(N__6627),
            .I(N__6624));
    Span12Mux_h I__1206 (
            .O(N__6624),
            .I(N__6621));
    Span12Mux_v I__1205 (
            .O(N__6621),
            .I(N__6618));
    Odrv12 I__1204 (
            .O(N__6618),
            .I(N_436_i));
    InMux I__1203 (
            .O(N__6615),
            .I(N__6609));
    InMux I__1202 (
            .O(N__6614),
            .I(N__6603));
    InMux I__1201 (
            .O(N__6613),
            .I(N__6600));
    InMux I__1200 (
            .O(N__6612),
            .I(N__6597));
    LocalMux I__1199 (
            .O(N__6609),
            .I(N__6594));
    CascadeMux I__1198 (
            .O(N__6608),
            .I(N__6591));
    CascadeMux I__1197 (
            .O(N__6607),
            .I(N__6587));
    CascadeMux I__1196 (
            .O(N__6606),
            .I(N__6583));
    LocalMux I__1195 (
            .O(N__6603),
            .I(N__6578));
    LocalMux I__1194 (
            .O(N__6600),
            .I(N__6578));
    LocalMux I__1193 (
            .O(N__6597),
            .I(N__6573));
    Span4Mux_v I__1192 (
            .O(N__6594),
            .I(N__6573));
    InMux I__1191 (
            .O(N__6591),
            .I(N__6570));
    InMux I__1190 (
            .O(N__6590),
            .I(N__6567));
    InMux I__1189 (
            .O(N__6587),
            .I(N__6564));
    InMux I__1188 (
            .O(N__6586),
            .I(N__6561));
    InMux I__1187 (
            .O(N__6583),
            .I(N__6558));
    Span4Mux_v I__1186 (
            .O(N__6578),
            .I(N__6551));
    Span4Mux_h I__1185 (
            .O(N__6573),
            .I(N__6551));
    LocalMux I__1184 (
            .O(N__6570),
            .I(N__6551));
    LocalMux I__1183 (
            .O(N__6567),
            .I(N__6548));
    LocalMux I__1182 (
            .O(N__6564),
            .I(N__6541));
    LocalMux I__1181 (
            .O(N__6561),
            .I(N__6541));
    LocalMux I__1180 (
            .O(N__6558),
            .I(N__6541));
    Sp12to4 I__1179 (
            .O(N__6551),
            .I(N__6538));
    Span4Mux_v I__1178 (
            .O(N__6548),
            .I(N__6533));
    Span4Mux_v I__1177 (
            .O(N__6541),
            .I(N__6533));
    Span12Mux_v I__1176 (
            .O(N__6538),
            .I(N__6528));
    Sp12to4 I__1175 (
            .O(N__6533),
            .I(N__6528));
    Span12Mux_h I__1174 (
            .O(N__6528),
            .I(N__6525));
    Span12Mux_v I__1173 (
            .O(N__6525),
            .I(N__6522));
    Odrv12 I__1172 (
            .O(N__6522),
            .I(A_c_17));
    InMux I__1171 (
            .O(N__6519),
            .I(N__6516));
    LocalMux I__1170 (
            .O(N__6516),
            .I(N__6512));
    InMux I__1169 (
            .O(N__6515),
            .I(N__6509));
    Odrv4 I__1168 (
            .O(N__6512),
            .I(N_431));
    LocalMux I__1167 (
            .O(N__6509),
            .I(N_431));
    CascadeMux I__1166 (
            .O(N__6504),
            .I(N__6501));
    InMux I__1165 (
            .O(N__6501),
            .I(N__6498));
    LocalMux I__1164 (
            .O(N__6498),
            .I(\U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_7 ));
    CascadeMux I__1163 (
            .O(N__6495),
            .I(N__6491));
    InMux I__1162 (
            .O(N__6494),
            .I(N__6488));
    InMux I__1161 (
            .O(N__6491),
            .I(N__6485));
    LocalMux I__1160 (
            .O(N__6488),
            .I(\U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_o2dupZ0 ));
    LocalMux I__1159 (
            .O(N__6485),
            .I(\U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_o2dupZ0 ));
    CascadeMux I__1158 (
            .O(N__6480),
            .I(\U409_ADDRESS_DECODE.un1_ATA_ENn_i_0Z0Z_3_cascade_ ));
    InMux I__1157 (
            .O(N__6477),
            .I(N__6471));
    InMux I__1156 (
            .O(N__6476),
            .I(N__6471));
    LocalMux I__1155 (
            .O(N__6471),
            .I(\U409_ADDRESS_DECODE.ATA_ENZ0 ));
    IoInMux I__1154 (
            .O(N__6468),
            .I(N__6465));
    LocalMux I__1153 (
            .O(N__6465),
            .I(N__6462));
    Span12Mux_s10_h I__1152 (
            .O(N__6462),
            .I(N__6459));
    Odrv12 I__1151 (
            .O(N__6459),
            .I(N_107));
    InMux I__1150 (
            .O(N__6456),
            .I(N__6452));
    InMux I__1149 (
            .O(N__6455),
            .I(N__6449));
    LocalMux I__1148 (
            .O(N__6452),
            .I(N__6443));
    LocalMux I__1147 (
            .O(N__6449),
            .I(N__6443));
    InMux I__1146 (
            .O(N__6448),
            .I(N__6440));
    Span4Mux_v I__1145 (
            .O(N__6443),
            .I(N__6437));
    LocalMux I__1144 (
            .O(N__6440),
            .I(N__6434));
    Span4Mux_v I__1143 (
            .O(N__6437),
            .I(N__6431));
    Span4Mux_v I__1142 (
            .O(N__6434),
            .I(N__6428));
    Span4Mux_v I__1141 (
            .O(N__6431),
            .I(N__6425));
    Sp12to4 I__1140 (
            .O(N__6428),
            .I(N__6422));
    Sp12to4 I__1139 (
            .O(N__6425),
            .I(N__6417));
    Span12Mux_v I__1138 (
            .O(N__6422),
            .I(N__6417));
    Odrv12 I__1137 (
            .O(N__6417),
            .I(A_c_16));
    InMux I__1136 (
            .O(N__6414),
            .I(N__6411));
    LocalMux I__1135 (
            .O(N__6411),
            .I(N__6407));
    CascadeMux I__1134 (
            .O(N__6410),
            .I(N__6404));
    Span4Mux_v I__1133 (
            .O(N__6407),
            .I(N__6401));
    InMux I__1132 (
            .O(N__6404),
            .I(N__6398));
    Odrv4 I__1131 (
            .O(N__6401),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ1Z_2 ));
    LocalMux I__1130 (
            .O(N__6398),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ1Z_2 ));
    InMux I__1129 (
            .O(N__6393),
            .I(N__6390));
    LocalMux I__1128 (
            .O(N__6390),
            .I(N__6386));
    InMux I__1127 (
            .O(N__6389),
            .I(N__6383));
    Odrv4 I__1126 (
            .O(N__6386),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ));
    LocalMux I__1125 (
            .O(N__6383),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ));
    CascadeMux I__1124 (
            .O(N__6378),
            .I(N__6373));
    InMux I__1123 (
            .O(N__6377),
            .I(N__6370));
    InMux I__1122 (
            .O(N__6376),
            .I(N__6367));
    InMux I__1121 (
            .O(N__6373),
            .I(N__6364));
    LocalMux I__1120 (
            .O(N__6370),
            .I(N__6359));
    LocalMux I__1119 (
            .O(N__6367),
            .I(N__6354));
    LocalMux I__1118 (
            .O(N__6364),
            .I(N__6354));
    InMux I__1117 (
            .O(N__6363),
            .I(N__6351));
    InMux I__1116 (
            .O(N__6362),
            .I(N__6348));
    Odrv4 I__1115 (
            .O(N__6359),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    Odrv4 I__1114 (
            .O(N__6354),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    LocalMux I__1113 (
            .O(N__6351),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    LocalMux I__1112 (
            .O(N__6348),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    IoInMux I__1111 (
            .O(N__6339),
            .I(N__6336));
    LocalMux I__1110 (
            .O(N__6336),
            .I(N__6333));
    IoSpan4Mux I__1109 (
            .O(N__6333),
            .I(N__6330));
    Sp12to4 I__1108 (
            .O(N__6330),
            .I(N__6327));
    Span12Mux_s9_v I__1107 (
            .O(N__6327),
            .I(N__6324));
    Odrv12 I__1106 (
            .O(N__6324),
            .I(N_128));
    InMux I__1105 (
            .O(N__6321),
            .I(N__6313));
    InMux I__1104 (
            .O(N__6320),
            .I(N__6313));
    InMux I__1103 (
            .O(N__6319),
            .I(N__6310));
    InMux I__1102 (
            .O(N__6318),
            .I(N__6307));
    LocalMux I__1101 (
            .O(N__6313),
            .I(N__6303));
    LocalMux I__1100 (
            .O(N__6310),
            .I(N__6300));
    LocalMux I__1099 (
            .O(N__6307),
            .I(N__6297));
    InMux I__1098 (
            .O(N__6306),
            .I(N__6294));
    Span4Mux_v I__1097 (
            .O(N__6303),
            .I(N__6291));
    Span4Mux_h I__1096 (
            .O(N__6300),
            .I(N__6284));
    Span4Mux_v I__1095 (
            .O(N__6297),
            .I(N__6284));
    LocalMux I__1094 (
            .O(N__6294),
            .I(N__6284));
    Span4Mux_v I__1093 (
            .O(N__6291),
            .I(N__6281));
    Span4Mux_v I__1092 (
            .O(N__6284),
            .I(N__6278));
    Sp12to4 I__1091 (
            .O(N__6281),
            .I(N__6275));
    Span4Mux_h I__1090 (
            .O(N__6278),
            .I(N__6272));
    Span12Mux_h I__1089 (
            .O(N__6275),
            .I(N__6267));
    Sp12to4 I__1088 (
            .O(N__6272),
            .I(N__6267));
    Odrv12 I__1087 (
            .O(N__6267),
            .I(TSn_c));
    CascadeMux I__1086 (
            .O(N__6264),
            .I(N__6257));
    InMux I__1085 (
            .O(N__6263),
            .I(N__6253));
    InMux I__1084 (
            .O(N__6262),
            .I(N__6248));
    InMux I__1083 (
            .O(N__6261),
            .I(N__6248));
    InMux I__1082 (
            .O(N__6260),
            .I(N__6241));
    InMux I__1081 (
            .O(N__6257),
            .I(N__6241));
    InMux I__1080 (
            .O(N__6256),
            .I(N__6241));
    LocalMux I__1079 (
            .O(N__6253),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__1078 (
            .O(N__6248),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__1077 (
            .O(N__6241),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    InMux I__1076 (
            .O(N__6234),
            .I(N__6230));
    InMux I__1075 (
            .O(N__6233),
            .I(N__6227));
    LocalMux I__1074 (
            .O(N__6230),
            .I(\U409_TRANSFER_ACK.N_268 ));
    LocalMux I__1073 (
            .O(N__6227),
            .I(\U409_TRANSFER_ACK.N_268 ));
    InMux I__1072 (
            .O(N__6222),
            .I(N__6218));
    InMux I__1071 (
            .O(N__6221),
            .I(N__6215));
    LocalMux I__1070 (
            .O(N__6218),
            .I(\U409_TRANSFER_ACK.N_237 ));
    LocalMux I__1069 (
            .O(N__6215),
            .I(\U409_TRANSFER_ACK.N_237 ));
    CascadeMux I__1068 (
            .O(N__6210),
            .I(N__6206));
    CascadeMux I__1067 (
            .O(N__6209),
            .I(N__6203));
    InMux I__1066 (
            .O(N__6206),
            .I(N__6200));
    InMux I__1065 (
            .O(N__6203),
            .I(N__6197));
    LocalMux I__1064 (
            .O(N__6200),
            .I(N__6192));
    LocalMux I__1063 (
            .O(N__6197),
            .I(N__6192));
    Span4Mux_v I__1062 (
            .O(N__6192),
            .I(N__6188));
    CascadeMux I__1061 (
            .O(N__6191),
            .I(N__6185));
    Span4Mux_v I__1060 (
            .O(N__6188),
            .I(N__6182));
    InMux I__1059 (
            .O(N__6185),
            .I(N__6179));
    Sp12to4 I__1058 (
            .O(N__6182),
            .I(N__6176));
    LocalMux I__1057 (
            .O(N__6179),
            .I(N__6173));
    Span12Mux_h I__1056 (
            .O(N__6176),
            .I(N__6168));
    Span12Mux_v I__1055 (
            .O(N__6173),
            .I(N__6168));
    Odrv12 I__1054 (
            .O(N__6168),
            .I(D_in_6));
    InMux I__1053 (
            .O(N__6165),
            .I(N__6161));
    InMux I__1052 (
            .O(N__6164),
            .I(N__6158));
    LocalMux I__1051 (
            .O(N__6161),
            .I(ATA_BASE_6));
    LocalMux I__1050 (
            .O(N__6158),
            .I(ATA_BASE_6));
    CascadeMux I__1049 (
            .O(N__6153),
            .I(N__6150));
    InMux I__1048 (
            .O(N__6150),
            .I(N__6146));
    InMux I__1047 (
            .O(N__6149),
            .I(N__6143));
    LocalMux I__1046 (
            .O(N__6146),
            .I(ATA_BASE_1));
    LocalMux I__1045 (
            .O(N__6143),
            .I(ATA_BASE_1));
    InMux I__1044 (
            .O(N__6138),
            .I(N__6134));
    InMux I__1043 (
            .O(N__6137),
            .I(N__6131));
    LocalMux I__1042 (
            .O(N__6134),
            .I(ATA_BASE_0));
    LocalMux I__1041 (
            .O(N__6131),
            .I(ATA_BASE_0));
    CascadeMux I__1040 (
            .O(N__6126),
            .I(\U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_7Z0Z_0_cascade_ ));
    CascadeMux I__1039 (
            .O(N__6123),
            .I(\U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_7_cascade_ ));
    CascadeMux I__1038 (
            .O(N__6120),
            .I(\U409_ADDRESS_DECODE.ATA_EN_2_0_o2_3_cascade_ ));
    InMux I__1037 (
            .O(N__6117),
            .I(N__6113));
    InMux I__1036 (
            .O(N__6116),
            .I(N__6108));
    LocalMux I__1035 (
            .O(N__6113),
            .I(N__6105));
    InMux I__1034 (
            .O(N__6112),
            .I(N__6102));
    InMux I__1033 (
            .O(N__6111),
            .I(N__6099));
    LocalMux I__1032 (
            .O(N__6108),
            .I(N__6092));
    Span4Mux_h I__1031 (
            .O(N__6105),
            .I(N__6092));
    LocalMux I__1030 (
            .O(N__6102),
            .I(N__6092));
    LocalMux I__1029 (
            .O(N__6099),
            .I(N__6089));
    Span4Mux_v I__1028 (
            .O(N__6092),
            .I(N__6085));
    Span4Mux_v I__1027 (
            .O(N__6089),
            .I(N__6082));
    InMux I__1026 (
            .O(N__6088),
            .I(N__6079));
    Sp12to4 I__1025 (
            .O(N__6085),
            .I(N__6072));
    Sp12to4 I__1024 (
            .O(N__6082),
            .I(N__6072));
    LocalMux I__1023 (
            .O(N__6079),
            .I(N__6072));
    Span12Mux_h I__1022 (
            .O(N__6072),
            .I(N__6069));
    Span12Mux_v I__1021 (
            .O(N__6069),
            .I(N__6066));
    Odrv12 I__1020 (
            .O(N__6066),
            .I(A_c_18));
    InMux I__1019 (
            .O(N__6063),
            .I(N__6059));
    InMux I__1018 (
            .O(N__6062),
            .I(N__6056));
    LocalMux I__1017 (
            .O(N__6059),
            .I(ATA_BASE_2));
    LocalMux I__1016 (
            .O(N__6056),
            .I(ATA_BASE_2));
    InMux I__1015 (
            .O(N__6051),
            .I(N__6048));
    LocalMux I__1014 (
            .O(N__6048),
            .I(\U409_ADDRESS_DECODE.N_183_i ));
    InMux I__1013 (
            .O(N__6045),
            .I(N__6042));
    LocalMux I__1012 (
            .O(N__6042),
            .I(\U409_ADDRESS_DECODE.ATA_EN_2_0_o2_2 ));
    InMux I__1011 (
            .O(N__6039),
            .I(N__6033));
    InMux I__1010 (
            .O(N__6038),
            .I(N__6033));
    LocalMux I__1009 (
            .O(N__6033),
            .I(\U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_2 ));
    InMux I__1008 (
            .O(N__6030),
            .I(N__6024));
    InMux I__1007 (
            .O(N__6029),
            .I(N__6024));
    LocalMux I__1006 (
            .O(N__6024),
            .I(N__6021));
    Span4Mux_v I__1005 (
            .O(N__6021),
            .I(N__6018));
    Span4Mux_v I__1004 (
            .O(N__6018),
            .I(N__6015));
    Odrv4 I__1003 (
            .O(N__6015),
            .I(\U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_0 ));
    CascadeMux I__1002 (
            .O(N__6012),
            .I(N__6008));
    InMux I__1001 (
            .O(N__6011),
            .I(N__6003));
    InMux I__1000 (
            .O(N__6008),
            .I(N__5996));
    InMux I__999 (
            .O(N__6007),
            .I(N__5996));
    InMux I__998 (
            .O(N__6006),
            .I(N__5993));
    LocalMux I__997 (
            .O(N__6003),
            .I(N__5990));
    InMux I__996 (
            .O(N__6002),
            .I(N__5985));
    InMux I__995 (
            .O(N__6001),
            .I(N__5985));
    LocalMux I__994 (
            .O(N__5996),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__993 (
            .O(N__5993),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    Odrv12 I__992 (
            .O(N__5990),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__991 (
            .O(N__5985),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    InMux I__990 (
            .O(N__5976),
            .I(N__5971));
    InMux I__989 (
            .O(N__5975),
            .I(N__5966));
    InMux I__988 (
            .O(N__5974),
            .I(N__5963));
    LocalMux I__987 (
            .O(N__5971),
            .I(N__5960));
    InMux I__986 (
            .O(N__5970),
            .I(N__5955));
    InMux I__985 (
            .O(N__5969),
            .I(N__5955));
    LocalMux I__984 (
            .O(N__5966),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__983 (
            .O(N__5963),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    Odrv4 I__982 (
            .O(N__5960),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__981 (
            .O(N__5955),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    InMux I__980 (
            .O(N__5946),
            .I(N__5943));
    LocalMux I__979 (
            .O(N__5943),
            .I(N__5939));
    CascadeMux I__978 (
            .O(N__5942),
            .I(N__5936));
    Span4Mux_v I__977 (
            .O(N__5939),
            .I(N__5933));
    InMux I__976 (
            .O(N__5936),
            .I(N__5930));
    Odrv4 I__975 (
            .O(N__5933),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ));
    LocalMux I__974 (
            .O(N__5930),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ));
    InMux I__973 (
            .O(N__5925),
            .I(N__5922));
    LocalMux I__972 (
            .O(N__5922),
            .I(N__5919));
    Span4Mux_v I__971 (
            .O(N__5919),
            .I(N__5915));
    InMux I__970 (
            .O(N__5918),
            .I(N__5912));
    Odrv4 I__969 (
            .O(N__5915),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ));
    LocalMux I__968 (
            .O(N__5912),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ));
    IoInMux I__967 (
            .O(N__5907),
            .I(N__5904));
    LocalMux I__966 (
            .O(N__5904),
            .I(N__5901));
    IoSpan4Mux I__965 (
            .O(N__5901),
            .I(N__5898));
    Span4Mux_s2_v I__964 (
            .O(N__5898),
            .I(N__5895));
    Sp12to4 I__963 (
            .O(N__5895),
            .I(N__5892));
    Odrv12 I__962 (
            .O(N__5892),
            .I(N_130));
    InMux I__961 (
            .O(N__5889),
            .I(N__5883));
    InMux I__960 (
            .O(N__5888),
            .I(N__5883));
    LocalMux I__959 (
            .O(N__5883),
            .I(ATA_BASE_4));
    InMux I__958 (
            .O(N__5880),
            .I(N__5874));
    InMux I__957 (
            .O(N__5879),
            .I(N__5874));
    LocalMux I__956 (
            .O(N__5874),
            .I(ATA_BASE_5));
    CascadeMux I__955 (
            .O(N__5871),
            .I(N__5866));
    InMux I__954 (
            .O(N__5870),
            .I(N__5861));
    InMux I__953 (
            .O(N__5869),
            .I(N__5861));
    InMux I__952 (
            .O(N__5866),
            .I(N__5858));
    LocalMux I__951 (
            .O(N__5861),
            .I(N__5855));
    LocalMux I__950 (
            .O(N__5858),
            .I(N__5852));
    Span4Mux_v I__949 (
            .O(N__5855),
            .I(N__5849));
    Span4Mux_v I__948 (
            .O(N__5852),
            .I(N__5846));
    Sp12to4 I__947 (
            .O(N__5849),
            .I(N__5841));
    Sp12to4 I__946 (
            .O(N__5846),
            .I(N__5841));
    Span12Mux_h I__945 (
            .O(N__5841),
            .I(N__5838));
    Odrv12 I__944 (
            .O(N__5838),
            .I(D_in_4));
    CascadeMux I__943 (
            .O(N__5835),
            .I(N__5832));
    InMux I__942 (
            .O(N__5832),
            .I(N__5826));
    InMux I__941 (
            .O(N__5831),
            .I(N__5826));
    LocalMux I__940 (
            .O(N__5826),
            .I(N__5823));
    Span4Mux_v I__939 (
            .O(N__5823),
            .I(N__5819));
    CascadeMux I__938 (
            .O(N__5822),
            .I(N__5816));
    Span4Mux_v I__937 (
            .O(N__5819),
            .I(N__5813));
    InMux I__936 (
            .O(N__5816),
            .I(N__5810));
    Sp12to4 I__935 (
            .O(N__5813),
            .I(N__5807));
    LocalMux I__934 (
            .O(N__5810),
            .I(N__5804));
    Span12Mux_h I__933 (
            .O(N__5807),
            .I(N__5799));
    Span12Mux_v I__932 (
            .O(N__5804),
            .I(N__5799));
    Odrv12 I__931 (
            .O(N__5799),
            .I(D_in_5));
    InMux I__930 (
            .O(N__5796),
            .I(N__5793));
    LocalMux I__929 (
            .O(N__5793),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3 ));
    InMux I__928 (
            .O(N__5790),
            .I(N__5782));
    InMux I__927 (
            .O(N__5789),
            .I(N__5782));
    InMux I__926 (
            .O(N__5788),
            .I(N__5777));
    InMux I__925 (
            .O(N__5787),
            .I(N__5777));
    LocalMux I__924 (
            .O(N__5782),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__923 (
            .O(N__5777),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    CascadeMux I__922 (
            .O(N__5772),
            .I(N__5768));
    InMux I__921 (
            .O(N__5771),
            .I(N__5764));
    InMux I__920 (
            .O(N__5768),
            .I(N__5759));
    InMux I__919 (
            .O(N__5767),
            .I(N__5759));
    LocalMux I__918 (
            .O(N__5764),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    LocalMux I__917 (
            .O(N__5759),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    CascadeMux I__916 (
            .O(N__5754),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_a2_3_cascade_ ));
    CascadeMux I__915 (
            .O(N__5751),
            .I(\U409_TRANSFER_ACK.N_268_cascade_ ));
    CascadeMux I__914 (
            .O(N__5748),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1_cascade_ ));
    CascadeMux I__913 (
            .O(N__5745),
            .I(N__5742));
    InMux I__912 (
            .O(N__5742),
            .I(N__5736));
    InMux I__911 (
            .O(N__5741),
            .I(N__5736));
    LocalMux I__910 (
            .O(N__5736),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ));
    CascadeMux I__909 (
            .O(N__5733),
            .I(N__5729));
    InMux I__908 (
            .O(N__5732),
            .I(N__5724));
    InMux I__907 (
            .O(N__5729),
            .I(N__5724));
    LocalMux I__906 (
            .O(N__5724),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ));
    InMux I__905 (
            .O(N__5721),
            .I(N__5718));
    LocalMux I__904 (
            .O(N__5718),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out ));
    CascadeMux I__903 (
            .O(N__5715),
            .I(N__5710));
    CascadeMux I__902 (
            .O(N__5714),
            .I(N__5707));
    InMux I__901 (
            .O(N__5713),
            .I(N__5703));
    InMux I__900 (
            .O(N__5710),
            .I(N__5696));
    InMux I__899 (
            .O(N__5707),
            .I(N__5696));
    InMux I__898 (
            .O(N__5706),
            .I(N__5696));
    LocalMux I__897 (
            .O(N__5703),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__896 (
            .O(N__5696),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    InMux I__895 (
            .O(N__5691),
            .I(N__5688));
    LocalMux I__894 (
            .O(N__5688),
            .I(N__5685));
    Span4Mux_h I__893 (
            .O(N__5685),
            .I(N__5680));
    InMux I__892 (
            .O(N__5684),
            .I(N__5677));
    InMux I__891 (
            .O(N__5683),
            .I(N__5674));
    Span4Mux_h I__890 (
            .O(N__5680),
            .I(N__5669));
    LocalMux I__889 (
            .O(N__5677),
            .I(N__5669));
    LocalMux I__888 (
            .O(N__5674),
            .I(N__5666));
    Span4Mux_h I__887 (
            .O(N__5669),
            .I(N__5663));
    Span12Mux_v I__886 (
            .O(N__5666),
            .I(N__5660));
    Span4Mux_v I__885 (
            .O(N__5663),
            .I(N__5657));
    Odrv12 I__884 (
            .O(N__5660),
            .I(A_c_31));
    Odrv4 I__883 (
            .O(N__5657),
            .I(A_c_31));
    InMux I__882 (
            .O(N__5652),
            .I(N__5648));
    InMux I__881 (
            .O(N__5651),
            .I(N__5645));
    LocalMux I__880 (
            .O(N__5648),
            .I(BRIDGE_BASE_3));
    LocalMux I__879 (
            .O(N__5645),
            .I(BRIDGE_BASE_3));
    CascadeMux I__878 (
            .O(N__5640),
            .I(N__5637));
    InMux I__877 (
            .O(N__5637),
            .I(N__5633));
    InMux I__876 (
            .O(N__5636),
            .I(N__5630));
    LocalMux I__875 (
            .O(N__5633),
            .I(BRIDGE_BASE_2));
    LocalMux I__874 (
            .O(N__5630),
            .I(BRIDGE_BASE_2));
    InMux I__873 (
            .O(N__5625),
            .I(N__5621));
    InMux I__872 (
            .O(N__5624),
            .I(N__5618));
    LocalMux I__871 (
            .O(N__5621),
            .I(N__5615));
    LocalMux I__870 (
            .O(N__5618),
            .I(N__5611));
    Span4Mux_h I__869 (
            .O(N__5615),
            .I(N__5608));
    InMux I__868 (
            .O(N__5614),
            .I(N__5605));
    Span4Mux_h I__867 (
            .O(N__5611),
            .I(N__5602));
    Span4Mux_h I__866 (
            .O(N__5608),
            .I(N__5597));
    LocalMux I__865 (
            .O(N__5605),
            .I(N__5597));
    Sp12to4 I__864 (
            .O(N__5602),
            .I(N__5594));
    Span4Mux_h I__863 (
            .O(N__5597),
            .I(N__5591));
    Span12Mux_v I__862 (
            .O(N__5594),
            .I(N__5588));
    Span4Mux_v I__861 (
            .O(N__5591),
            .I(N__5585));
    Odrv12 I__860 (
            .O(N__5588),
            .I(A_c_30));
    Odrv4 I__859 (
            .O(N__5585),
            .I(A_c_30));
    InMux I__858 (
            .O(N__5580),
            .I(N__5577));
    LocalMux I__857 (
            .O(N__5577),
            .I(\U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0Z0Z_1 ));
    InMux I__856 (
            .O(N__5574),
            .I(N__5562));
    InMux I__855 (
            .O(N__5573),
            .I(N__5562));
    InMux I__854 (
            .O(N__5572),
            .I(N__5562));
    InMux I__853 (
            .O(N__5571),
            .I(N__5562));
    LocalMux I__852 (
            .O(N__5562),
            .I(\U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa ));
    InMux I__851 (
            .O(N__5559),
            .I(N__5553));
    InMux I__850 (
            .O(N__5558),
            .I(N__5548));
    InMux I__849 (
            .O(N__5557),
            .I(N__5548));
    InMux I__848 (
            .O(N__5556),
            .I(N__5545));
    LocalMux I__847 (
            .O(N__5553),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    LocalMux I__846 (
            .O(N__5548),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    LocalMux I__845 (
            .O(N__5545),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    InMux I__844 (
            .O(N__5538),
            .I(N__5529));
    InMux I__843 (
            .O(N__5537),
            .I(N__5529));
    InMux I__842 (
            .O(N__5536),
            .I(N__5529));
    LocalMux I__841 (
            .O(N__5529),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_o2_5));
    InMux I__840 (
            .O(N__5526),
            .I(N__5522));
    CascadeMux I__839 (
            .O(N__5525),
            .I(N__5519));
    LocalMux I__838 (
            .O(N__5522),
            .I(N__5516));
    InMux I__837 (
            .O(N__5519),
            .I(N__5513));
    Span4Mux_v I__836 (
            .O(N__5516),
            .I(N__5508));
    LocalMux I__835 (
            .O(N__5513),
            .I(N__5508));
    Odrv4 I__834 (
            .O(N__5508),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ));
    InMux I__833 (
            .O(N__5505),
            .I(N__5502));
    LocalMux I__832 (
            .O(N__5502),
            .I(N__5499));
    Span4Mux_v I__831 (
            .O(N__5499),
            .I(N__5495));
    InMux I__830 (
            .O(N__5498),
            .I(N__5492));
    Odrv4 I__829 (
            .O(N__5495),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ));
    LocalMux I__828 (
            .O(N__5492),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ));
    IoInMux I__827 (
            .O(N__5487),
            .I(N__5484));
    LocalMux I__826 (
            .O(N__5484),
            .I(N__5481));
    Sp12to4 I__825 (
            .O(N__5481),
            .I(N__5478));
    Span12Mux_s10_v I__824 (
            .O(N__5478),
            .I(N__5475));
    Odrv12 I__823 (
            .O(N__5475),
            .I(N_126));
    IoInMux I__822 (
            .O(N__5472),
            .I(N__5469));
    LocalMux I__821 (
            .O(N__5469),
            .I(N__5466));
    IoSpan4Mux I__820 (
            .O(N__5466),
            .I(N__5463));
    Span4Mux_s1_h I__819 (
            .O(N__5463),
            .I(N__5460));
    Sp12to4 I__818 (
            .O(N__5460),
            .I(N__5457));
    Span12Mux_h I__817 (
            .O(N__5457),
            .I(N__5454));
    Odrv12 I__816 (
            .O(N__5454),
            .I(N_96));
    CascadeMux I__815 (
            .O(N__5451),
            .I(N__5448));
    InMux I__814 (
            .O(N__5448),
            .I(N__5443));
    InMux I__813 (
            .O(N__5447),
            .I(N__5440));
    InMux I__812 (
            .O(N__5446),
            .I(N__5437));
    LocalMux I__811 (
            .O(N__5443),
            .I(N__5432));
    LocalMux I__810 (
            .O(N__5440),
            .I(N__5432));
    LocalMux I__809 (
            .O(N__5437),
            .I(N__5429));
    Span4Mux_v I__808 (
            .O(N__5432),
            .I(N__5426));
    Span12Mux_h I__807 (
            .O(N__5429),
            .I(N__5423));
    Span4Mux_v I__806 (
            .O(N__5426),
            .I(N__5420));
    Span12Mux_v I__805 (
            .O(N__5423),
            .I(N__5417));
    Sp12to4 I__804 (
            .O(N__5420),
            .I(N__5414));
    Odrv12 I__803 (
            .O(N__5417),
            .I(A_c_29));
    Odrv12 I__802 (
            .O(N__5414),
            .I(A_c_29));
    InMux I__801 (
            .O(N__5409),
            .I(N__5405));
    InMux I__800 (
            .O(N__5408),
            .I(N__5402));
    LocalMux I__799 (
            .O(N__5405),
            .I(BRIDGE_BASE_1));
    LocalMux I__798 (
            .O(N__5402),
            .I(BRIDGE_BASE_1));
    InMux I__797 (
            .O(N__5397),
            .I(N__5392));
    CascadeMux I__796 (
            .O(N__5396),
            .I(N__5389));
    CascadeMux I__795 (
            .O(N__5395),
            .I(N__5386));
    LocalMux I__794 (
            .O(N__5392),
            .I(N__5383));
    InMux I__793 (
            .O(N__5389),
            .I(N__5380));
    InMux I__792 (
            .O(N__5386),
            .I(N__5377));
    Span4Mux_v I__791 (
            .O(N__5383),
            .I(N__5374));
    LocalMux I__790 (
            .O(N__5380),
            .I(N__5371));
    LocalMux I__789 (
            .O(N__5377),
            .I(N__5368));
    Span4Mux_v I__788 (
            .O(N__5374),
            .I(N__5365));
    Span12Mux_v I__787 (
            .O(N__5371),
            .I(N__5360));
    Sp12to4 I__786 (
            .O(N__5368),
            .I(N__5360));
    Span4Mux_v I__785 (
            .O(N__5365),
            .I(N__5357));
    Span12Mux_v I__784 (
            .O(N__5360),
            .I(N__5354));
    Span4Mux_h I__783 (
            .O(N__5357),
            .I(N__5351));
    Odrv12 I__782 (
            .O(N__5354),
            .I(A_c_28));
    Odrv4 I__781 (
            .O(N__5351),
            .I(A_c_28));
    InMux I__780 (
            .O(N__5346),
            .I(N__5342));
    InMux I__779 (
            .O(N__5345),
            .I(N__5339));
    LocalMux I__778 (
            .O(N__5342),
            .I(BRIDGE_BASE_0));
    LocalMux I__777 (
            .O(N__5339),
            .I(BRIDGE_BASE_0));
    InMux I__776 (
            .O(N__5334),
            .I(N__5331));
    LocalMux I__775 (
            .O(N__5331),
            .I(\U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0Z0Z_0 ));
    IoInMux I__774 (
            .O(N__5328),
            .I(N__5325));
    LocalMux I__773 (
            .O(N__5325),
            .I(N__5320));
    IoInMux I__772 (
            .O(N__5324),
            .I(N__5317));
    IoInMux I__771 (
            .O(N__5323),
            .I(N__5314));
    IoSpan4Mux I__770 (
            .O(N__5320),
            .I(N__5307));
    LocalMux I__769 (
            .O(N__5317),
            .I(N__5307));
    LocalMux I__768 (
            .O(N__5314),
            .I(N__5307));
    IoSpan4Mux I__767 (
            .O(N__5307),
            .I(N__5303));
    IoInMux I__766 (
            .O(N__5306),
            .I(N__5300));
    Span4Mux_s2_v I__765 (
            .O(N__5303),
            .I(N__5297));
    LocalMux I__764 (
            .O(N__5300),
            .I(N__5294));
    Sp12to4 I__763 (
            .O(N__5297),
            .I(N__5289));
    Span12Mux_s4_v I__762 (
            .O(N__5294),
            .I(N__5289));
    Odrv12 I__761 (
            .O(N__5289),
            .I(D_1_i));
    InMux I__760 (
            .O(N__5286),
            .I(N__5283));
    LocalMux I__759 (
            .O(N__5283),
            .I(N__5280));
    Span4Mux_v I__758 (
            .O(N__5280),
            .I(N__5277));
    Sp12to4 I__757 (
            .O(N__5277),
            .I(N__5274));
    Span12Mux_h I__756 (
            .O(N__5274),
            .I(N__5271));
    Span12Mux_h I__755 (
            .O(N__5271),
            .I(N__5268));
    Span12Mux_v I__754 (
            .O(N__5268),
            .I(N__5265));
    Odrv12 I__753 (
            .O(N__5265),
            .I(AUTOBOOT_c));
    InMux I__752 (
            .O(N__5262),
            .I(N__5258));
    InMux I__751 (
            .O(N__5261),
            .I(N__5255));
    LocalMux I__750 (
            .O(N__5258),
            .I(\U409_AUTOCONFIG.N_360 ));
    LocalMux I__749 (
            .O(N__5255),
            .I(\U409_AUTOCONFIG.N_360 ));
    CascadeMux I__748 (
            .O(N__5250),
            .I(N__5244));
    InMux I__747 (
            .O(N__5249),
            .I(N__5241));
    InMux I__746 (
            .O(N__5248),
            .I(N__5236));
    InMux I__745 (
            .O(N__5247),
            .I(N__5236));
    InMux I__744 (
            .O(N__5244),
            .I(N__5233));
    LocalMux I__743 (
            .O(N__5241),
            .I(N__5224));
    LocalMux I__742 (
            .O(N__5236),
            .I(N__5221));
    LocalMux I__741 (
            .O(N__5233),
            .I(N__5218));
    InMux I__740 (
            .O(N__5232),
            .I(N__5211));
    InMux I__739 (
            .O(N__5231),
            .I(N__5211));
    InMux I__738 (
            .O(N__5230),
            .I(N__5211));
    CascadeMux I__737 (
            .O(N__5229),
            .I(N__5208));
    CascadeMux I__736 (
            .O(N__5228),
            .I(N__5205));
    CascadeMux I__735 (
            .O(N__5227),
            .I(N__5201));
    Span4Mux_v I__734 (
            .O(N__5224),
            .I(N__5196));
    Span4Mux_v I__733 (
            .O(N__5221),
            .I(N__5196));
    Span4Mux_v I__732 (
            .O(N__5218),
            .I(N__5191));
    LocalMux I__731 (
            .O(N__5211),
            .I(N__5191));
    InMux I__730 (
            .O(N__5208),
            .I(N__5182));
    InMux I__729 (
            .O(N__5205),
            .I(N__5182));
    InMux I__728 (
            .O(N__5204),
            .I(N__5182));
    InMux I__727 (
            .O(N__5201),
            .I(N__5182));
    Sp12to4 I__726 (
            .O(N__5196),
            .I(N__5175));
    Sp12to4 I__725 (
            .O(N__5191),
            .I(N__5175));
    LocalMux I__724 (
            .O(N__5182),
            .I(N__5175));
    Odrv12 I__723 (
            .O(N__5175),
            .I(A_c_5));
    InMux I__722 (
            .O(N__5172),
            .I(N__5169));
    LocalMux I__721 (
            .O(N__5169),
            .I(N__5162));
    InMux I__720 (
            .O(N__5168),
            .I(N__5155));
    InMux I__719 (
            .O(N__5167),
            .I(N__5155));
    InMux I__718 (
            .O(N__5166),
            .I(N__5155));
    InMux I__717 (
            .O(N__5165),
            .I(N__5148));
    Span4Mux_h I__716 (
            .O(N__5162),
            .I(N__5143));
    LocalMux I__715 (
            .O(N__5155),
            .I(N__5143));
    InMux I__714 (
            .O(N__5154),
            .I(N__5140));
    InMux I__713 (
            .O(N__5153),
            .I(N__5137));
    InMux I__712 (
            .O(N__5152),
            .I(N__5132));
    InMux I__711 (
            .O(N__5151),
            .I(N__5132));
    LocalMux I__710 (
            .O(N__5148),
            .I(N__5125));
    Span4Mux_h I__709 (
            .O(N__5143),
            .I(N__5125));
    LocalMux I__708 (
            .O(N__5140),
            .I(N__5125));
    LocalMux I__707 (
            .O(N__5137),
            .I(N__5120));
    LocalMux I__706 (
            .O(N__5132),
            .I(N__5120));
    Sp12to4 I__705 (
            .O(N__5125),
            .I(N__5117));
    Span12Mux_h I__704 (
            .O(N__5120),
            .I(N__5114));
    Span12Mux_v I__703 (
            .O(N__5117),
            .I(N__5111));
    Span12Mux_v I__702 (
            .O(N__5114),
            .I(N__5108));
    Odrv12 I__701 (
            .O(N__5111),
            .I(A_c_3));
    Odrv12 I__700 (
            .O(N__5108),
            .I(A_c_3));
    CascadeMux I__699 (
            .O(N__5103),
            .I(N__5100));
    InMux I__698 (
            .O(N__5100),
            .I(N__5097));
    LocalMux I__697 (
            .O(N__5097),
            .I(N__5094));
    Span4Mux_v I__696 (
            .O(N__5094),
            .I(N__5091));
    Odrv4 I__695 (
            .O(N__5091),
            .I(\U409_AUTOCONFIG.N_276 ));
    CascadeMux I__694 (
            .O(N__5088),
            .I(\U409_ADDRESS_DECODE.PORTSIZE_iZ0Z_1_cascade_ ));
    IoInMux I__693 (
            .O(N__5085),
            .I(N__5082));
    LocalMux I__692 (
            .O(N__5082),
            .I(N__5079));
    IoSpan4Mux I__691 (
            .O(N__5079),
            .I(N__5076));
    Span4Mux_s2_v I__690 (
            .O(N__5076),
            .I(N__5073));
    Sp12to4 I__689 (
            .O(N__5073),
            .I(N__5070));
    Odrv12 I__688 (
            .O(N__5070),
            .I(N_139));
    InMux I__687 (
            .O(N__5067),
            .I(N__5064));
    LocalMux I__686 (
            .O(N__5064),
            .I(N__5061));
    Span4Mux_v I__685 (
            .O(N__5061),
            .I(N__5058));
    Odrv4 I__684 (
            .O(N__5058),
            .I(\U409_ADDRESS_DECODE.N_343 ));
    InMux I__683 (
            .O(N__5055),
            .I(N__5051));
    InMux I__682 (
            .O(N__5054),
            .I(N__5048));
    LocalMux I__681 (
            .O(N__5051),
            .I(N__5043));
    LocalMux I__680 (
            .O(N__5048),
            .I(N__5043));
    Span4Mux_v I__679 (
            .O(N__5043),
            .I(N__5039));
    InMux I__678 (
            .O(N__5042),
            .I(N__5036));
    Span4Mux_h I__677 (
            .O(N__5039),
            .I(N__5033));
    LocalMux I__676 (
            .O(N__5036),
            .I(N__5030));
    Sp12to4 I__675 (
            .O(N__5033),
            .I(N__5027));
    Span12Mux_h I__674 (
            .O(N__5030),
            .I(N__5024));
    Odrv12 I__673 (
            .O(N__5027),
            .I(TM_c_1));
    Odrv12 I__672 (
            .O(N__5024),
            .I(TM_c_1));
    InMux I__671 (
            .O(N__5019),
            .I(N__5015));
    InMux I__670 (
            .O(N__5018),
            .I(N__5012));
    LocalMux I__669 (
            .O(N__5015),
            .I(N__5006));
    LocalMux I__668 (
            .O(N__5012),
            .I(N__5006));
    InMux I__667 (
            .O(N__5011),
            .I(N__5003));
    Span4Mux_v I__666 (
            .O(N__5006),
            .I(N__4998));
    LocalMux I__665 (
            .O(N__5003),
            .I(N__4998));
    Span4Mux_h I__664 (
            .O(N__4998),
            .I(N__4995));
    Sp12to4 I__663 (
            .O(N__4995),
            .I(N__4992));
    Odrv12 I__662 (
            .O(N__4992),
            .I(TM_c_0));
    IoInMux I__661 (
            .O(N__4989),
            .I(N__4986));
    LocalMux I__660 (
            .O(N__4986),
            .I(N__4983));
    Span12Mux_s11_v I__659 (
            .O(N__4983),
            .I(N__4980));
    Span12Mux_h I__658 (
            .O(N__4980),
            .I(N__4977));
    Odrv12 I__657 (
            .O(N__4977),
            .I(N_265_i));
    CascadeMux I__656 (
            .O(N__4974),
            .I(N__4969));
    CascadeMux I__655 (
            .O(N__4973),
            .I(N__4966));
    InMux I__654 (
            .O(N__4972),
            .I(N__4959));
    InMux I__653 (
            .O(N__4969),
            .I(N__4959));
    InMux I__652 (
            .O(N__4966),
            .I(N__4959));
    LocalMux I__651 (
            .O(N__4959),
            .I(N__4956));
    Odrv12 I__650 (
            .O(N__4956),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_o2_4));
    InMux I__649 (
            .O(N__4953),
            .I(N__4949));
    InMux I__648 (
            .O(N__4952),
            .I(N__4946));
    LocalMux I__647 (
            .O(N__4949),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ1Z_0 ));
    LocalMux I__646 (
            .O(N__4946),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ1Z_0 ));
    CascadeMux I__645 (
            .O(N__4941),
            .I(N__4938));
    InMux I__644 (
            .O(N__4938),
            .I(N__4935));
    LocalMux I__643 (
            .O(N__4935),
            .I(N__4931));
    InMux I__642 (
            .O(N__4934),
            .I(N__4928));
    Odrv4 I__641 (
            .O(N__4931),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ1Z_0 ));
    LocalMux I__640 (
            .O(N__4928),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ1Z_0 ));
    IoInMux I__639 (
            .O(N__4923),
            .I(N__4920));
    LocalMux I__638 (
            .O(N__4920),
            .I(N__4917));
    Span12Mux_s2_v I__637 (
            .O(N__4917),
            .I(N__4914));
    Odrv12 I__636 (
            .O(N__4914),
            .I(N_124));
    CascadeMux I__635 (
            .O(N__4911),
            .I(N__4908));
    InMux I__634 (
            .O(N__4908),
            .I(N__4905));
    LocalMux I__633 (
            .O(N__4905),
            .I(\U409_AUTOCONFIG.un1_STATE_1_0_a2_0Z0Z_2 ));
    CascadeMux I__632 (
            .O(N__4902),
            .I(N__4899));
    InMux I__631 (
            .O(N__4899),
            .I(N__4896));
    LocalMux I__630 (
            .O(N__4896),
            .I(N__4892));
    InMux I__629 (
            .O(N__4895),
            .I(N__4889));
    Sp12to4 I__628 (
            .O(N__4892),
            .I(N__4884));
    LocalMux I__627 (
            .O(N__4889),
            .I(N__4884));
    Span12Mux_v I__626 (
            .O(N__4884),
            .I(N__4881));
    Odrv12 I__625 (
            .O(N__4881),
            .I(CPUCONFn_c));
    InMux I__624 (
            .O(N__4878),
            .I(N__4874));
    InMux I__623 (
            .O(N__4877),
            .I(N__4871));
    LocalMux I__622 (
            .O(N__4874),
            .I(\U409_AUTOCONFIG.AC_STARTZ0 ));
    LocalMux I__621 (
            .O(N__4871),
            .I(\U409_AUTOCONFIG.AC_STARTZ0 ));
    CascadeMux I__620 (
            .O(N__4866),
            .I(N_354_cascade_));
    InMux I__619 (
            .O(N__4863),
            .I(N__4860));
    LocalMux I__618 (
            .O(N__4860),
            .I(N__4857));
    Odrv4 I__617 (
            .O(N__4857),
            .I(\U409_AUTOCONFIG.N_273 ));
    CascadeMux I__616 (
            .O(N__4854),
            .I(N__4850));
    InMux I__615 (
            .O(N__4853),
            .I(N__4845));
    InMux I__614 (
            .O(N__4850),
            .I(N__4845));
    LocalMux I__613 (
            .O(N__4845),
            .I(\U409_AUTOCONFIG.N_400 ));
    CascadeMux I__612 (
            .O(N__4842),
            .I(N__4837));
    InMux I__611 (
            .O(N__4841),
            .I(N__4831));
    InMux I__610 (
            .O(N__4840),
            .I(N__4827));
    InMux I__609 (
            .O(N__4837),
            .I(N__4818));
    InMux I__608 (
            .O(N__4836),
            .I(N__4818));
    InMux I__607 (
            .O(N__4835),
            .I(N__4818));
    InMux I__606 (
            .O(N__4834),
            .I(N__4818));
    LocalMux I__605 (
            .O(N__4831),
            .I(N__4813));
    InMux I__604 (
            .O(N__4830),
            .I(N__4806));
    LocalMux I__603 (
            .O(N__4827),
            .I(N__4801));
    LocalMux I__602 (
            .O(N__4818),
            .I(N__4801));
    InMux I__601 (
            .O(N__4817),
            .I(N__4796));
    InMux I__600 (
            .O(N__4816),
            .I(N__4796));
    Span4Mux_v I__599 (
            .O(N__4813),
            .I(N__4793));
    InMux I__598 (
            .O(N__4812),
            .I(N__4786));
    InMux I__597 (
            .O(N__4811),
            .I(N__4786));
    InMux I__596 (
            .O(N__4810),
            .I(N__4786));
    InMux I__595 (
            .O(N__4809),
            .I(N__4783));
    LocalMux I__594 (
            .O(N__4806),
            .I(N__4780));
    Span4Mux_v I__593 (
            .O(N__4801),
            .I(N__4775));
    LocalMux I__592 (
            .O(N__4796),
            .I(N__4775));
    Sp12to4 I__591 (
            .O(N__4793),
            .I(N__4768));
    LocalMux I__590 (
            .O(N__4786),
            .I(N__4768));
    LocalMux I__589 (
            .O(N__4783),
            .I(N__4768));
    Span4Mux_v I__588 (
            .O(N__4780),
            .I(N__4765));
    Span4Mux_v I__587 (
            .O(N__4775),
            .I(N__4762));
    Span12Mux_h I__586 (
            .O(N__4768),
            .I(N__4759));
    Sp12to4 I__585 (
            .O(N__4765),
            .I(N__4754));
    Sp12to4 I__584 (
            .O(N__4762),
            .I(N__4754));
    Span12Mux_v I__583 (
            .O(N__4759),
            .I(N__4751));
    Span12Mux_h I__582 (
            .O(N__4754),
            .I(N__4748));
    Odrv12 I__581 (
            .O(N__4751),
            .I(A_c_2));
    Odrv12 I__580 (
            .O(N__4748),
            .I(A_c_2));
    CascadeMux I__579 (
            .O(N__4743),
            .I(N__4733));
    CascadeMux I__578 (
            .O(N__4742),
            .I(N__4729));
    CascadeMux I__577 (
            .O(N__4741),
            .I(N__4726));
    CascadeMux I__576 (
            .O(N__4740),
            .I(N__4722));
    InMux I__575 (
            .O(N__4739),
            .I(N__4718));
    InMux I__574 (
            .O(N__4738),
            .I(N__4711));
    InMux I__573 (
            .O(N__4737),
            .I(N__4711));
    InMux I__572 (
            .O(N__4736),
            .I(N__4711));
    InMux I__571 (
            .O(N__4733),
            .I(N__4704));
    InMux I__570 (
            .O(N__4732),
            .I(N__4704));
    InMux I__569 (
            .O(N__4729),
            .I(N__4704));
    InMux I__568 (
            .O(N__4726),
            .I(N__4699));
    InMux I__567 (
            .O(N__4725),
            .I(N__4699));
    InMux I__566 (
            .O(N__4722),
            .I(N__4696));
    InMux I__565 (
            .O(N__4721),
            .I(N__4693));
    LocalMux I__564 (
            .O(N__4718),
            .I(N__4687));
    LocalMux I__563 (
            .O(N__4711),
            .I(N__4687));
    LocalMux I__562 (
            .O(N__4704),
            .I(N__4684));
    LocalMux I__561 (
            .O(N__4699),
            .I(N__4677));
    LocalMux I__560 (
            .O(N__4696),
            .I(N__4677));
    LocalMux I__559 (
            .O(N__4693),
            .I(N__4677));
    CascadeMux I__558 (
            .O(N__4692),
            .I(N__4673));
    Span4Mux_v I__557 (
            .O(N__4687),
            .I(N__4669));
    Span4Mux_v I__556 (
            .O(N__4684),
            .I(N__4664));
    Span4Mux_v I__555 (
            .O(N__4677),
            .I(N__4664));
    InMux I__554 (
            .O(N__4676),
            .I(N__4661));
    InMux I__553 (
            .O(N__4673),
            .I(N__4658));
    InMux I__552 (
            .O(N__4672),
            .I(N__4655));
    Sp12to4 I__551 (
            .O(N__4669),
            .I(N__4644));
    Sp12to4 I__550 (
            .O(N__4664),
            .I(N__4644));
    LocalMux I__549 (
            .O(N__4661),
            .I(N__4644));
    LocalMux I__548 (
            .O(N__4658),
            .I(N__4644));
    LocalMux I__547 (
            .O(N__4655),
            .I(N__4644));
    Odrv12 I__546 (
            .O(N__4644),
            .I(A_c_4));
    InMux I__545 (
            .O(N__4641),
            .I(N__4638));
    LocalMux I__544 (
            .O(N__4638),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_10 ));
    InMux I__543 (
            .O(N__4635),
            .I(N__4632));
    LocalMux I__542 (
            .O(N__4632),
            .I(N__4629));
    Span4Mux_h I__541 (
            .O(N__4629),
            .I(N__4626));
    Span4Mux_h I__540 (
            .O(N__4626),
            .I(N__4623));
    Odrv4 I__539 (
            .O(N__4623),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_11 ));
    CascadeMux I__538 (
            .O(N__4620),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_9_cascade_ ));
    CascadeMux I__537 (
            .O(N__4617),
            .I(N__4613));
    InMux I__536 (
            .O(N__4616),
            .I(N__4608));
    InMux I__535 (
            .O(N__4613),
            .I(N__4608));
    LocalMux I__534 (
            .O(N__4608),
            .I(N__4605));
    Odrv4 I__533 (
            .O(N__4605),
            .I(N_374));
    CascadeMux I__532 (
            .O(N__4602),
            .I(N_401_cascade_));
    InMux I__531 (
            .O(N__4599),
            .I(N__4596));
    LocalMux I__530 (
            .O(N__4596),
            .I(N_436));
    InMux I__529 (
            .O(N__4593),
            .I(N__4590));
    LocalMux I__528 (
            .O(N__4590),
            .I(\U409_AUTOCONFIG.N_285 ));
    InMux I__527 (
            .O(N__4587),
            .I(N__4584));
    LocalMux I__526 (
            .O(N__4584),
            .I(\U409_AUTOCONFIG.N_9 ));
    InMux I__525 (
            .O(N__4581),
            .I(N__4578));
    LocalMux I__524 (
            .O(N__4578),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_0_1 ));
    InMux I__523 (
            .O(N__4575),
            .I(N__4563));
    InMux I__522 (
            .O(N__4574),
            .I(N__4563));
    InMux I__521 (
            .O(N__4573),
            .I(N__4563));
    InMux I__520 (
            .O(N__4572),
            .I(N__4563));
    LocalMux I__519 (
            .O(N__4563),
            .I(\U409_AUTOCONFIG.N_405 ));
    InMux I__518 (
            .O(N__4560),
            .I(N__4557));
    LocalMux I__517 (
            .O(N__4557),
            .I(N__4554));
    Odrv4 I__516 (
            .O(N__4554),
            .I(\U409_AUTOCONFIG.LIDE_OUTc_0_1 ));
    CascadeMux I__515 (
            .O(N__4551),
            .I(N__4548));
    InMux I__514 (
            .O(N__4548),
            .I(N__4545));
    LocalMux I__513 (
            .O(N__4545),
            .I(N__4542));
    Odrv4 I__512 (
            .O(N__4542),
            .I(\U409_AUTOCONFIG.LIDE_OUTc_0_0 ));
    InMux I__511 (
            .O(N__4539),
            .I(N__4536));
    LocalMux I__510 (
            .O(N__4536),
            .I(\U409_AUTOCONFIG.N_286 ));
    InMux I__509 (
            .O(N__4533),
            .I(N__4521));
    InMux I__508 (
            .O(N__4532),
            .I(N__4521));
    InMux I__507 (
            .O(N__4531),
            .I(N__4521));
    InMux I__506 (
            .O(N__4530),
            .I(N__4521));
    LocalMux I__505 (
            .O(N__4521),
            .I(\U409_AUTOCONFIG.AC_START_RNI3D7VZ0Z2 ));
    InMux I__504 (
            .O(N__4518),
            .I(N__4515));
    LocalMux I__503 (
            .O(N__4515),
            .I(\U409_AUTOCONFIG.N_287 ));
    InMux I__502 (
            .O(N__4512),
            .I(N__4508));
    CascadeMux I__501 (
            .O(N__4511),
            .I(N__4505));
    LocalMux I__500 (
            .O(N__4508),
            .I(N__4501));
    InMux I__499 (
            .O(N__4505),
            .I(N__4498));
    InMux I__498 (
            .O(N__4504),
            .I(N__4495));
    Span4Mux_v I__497 (
            .O(N__4501),
            .I(N__4489));
    LocalMux I__496 (
            .O(N__4498),
            .I(N__4484));
    LocalMux I__495 (
            .O(N__4495),
            .I(N__4484));
    InMux I__494 (
            .O(N__4494),
            .I(N__4477));
    InMux I__493 (
            .O(N__4493),
            .I(N__4477));
    InMux I__492 (
            .O(N__4492),
            .I(N__4477));
    Sp12to4 I__491 (
            .O(N__4489),
            .I(N__4470));
    Sp12to4 I__490 (
            .O(N__4484),
            .I(N__4470));
    LocalMux I__489 (
            .O(N__4477),
            .I(N__4470));
    Odrv12 I__488 (
            .O(N__4470),
            .I(A_c_6));
    InMux I__487 (
            .O(N__4467),
            .I(N__4454));
    InMux I__486 (
            .O(N__4466),
            .I(N__4454));
    InMux I__485 (
            .O(N__4465),
            .I(N__4454));
    InMux I__484 (
            .O(N__4464),
            .I(N__4454));
    InMux I__483 (
            .O(N__4463),
            .I(N__4451));
    LocalMux I__482 (
            .O(N__4454),
            .I(N__4448));
    LocalMux I__481 (
            .O(N__4451),
            .I(N__4444));
    Span4Mux_v I__480 (
            .O(N__4448),
            .I(N__4441));
    InMux I__479 (
            .O(N__4447),
            .I(N__4438));
    Span12Mux_v I__478 (
            .O(N__4444),
            .I(N__4431));
    Sp12to4 I__477 (
            .O(N__4441),
            .I(N__4431));
    LocalMux I__476 (
            .O(N__4438),
            .I(N__4431));
    Odrv12 I__475 (
            .O(N__4431),
            .I(A_c_7));
    InMux I__474 (
            .O(N__4428),
            .I(N__4425));
    LocalMux I__473 (
            .O(N__4425),
            .I(\U409_AUTOCONFIG.N_274 ));
    CascadeMux I__472 (
            .O(N__4422),
            .I(\U409_AUTOCONFIG.N_383_cascade_ ));
    InMux I__471 (
            .O(N__4419),
            .I(N__4416));
    LocalMux I__470 (
            .O(N__4416),
            .I(N__4413));
    Span4Mux_h I__469 (
            .O(N__4413),
            .I(N__4410));
    Sp12to4 I__468 (
            .O(N__4410),
            .I(N__4407));
    Odrv12 I__467 (
            .O(N__4407),
            .I(TT_c_0));
    InMux I__466 (
            .O(N__4404),
            .I(N__4401));
    LocalMux I__465 (
            .O(N__4401),
            .I(N__4398));
    Span12Mux_h I__464 (
            .O(N__4398),
            .I(N__4395));
    Odrv12 I__463 (
            .O(N__4395),
            .I(TT_c_1));
    CascadeMux I__462 (
            .O(N__4392),
            .I(N__4389));
    InMux I__461 (
            .O(N__4389),
            .I(N__4386));
    LocalMux I__460 (
            .O(N__4386),
            .I(\U409_ADDRESS_DECODE.N_345 ));
    InMux I__459 (
            .O(N__4383),
            .I(N__4380));
    LocalMux I__458 (
            .O(N__4380),
            .I(\U409_ADDRESS_DECODE.N_344 ));
    CascadeMux I__457 (
            .O(N__4377),
            .I(\U409_AUTOCONFIG.N_288_cascade_ ));
    InMux I__456 (
            .O(N__4374),
            .I(N__4371));
    LocalMux I__455 (
            .O(N__4371),
            .I(N__4368));
    Odrv4 I__454 (
            .O(N__4368),
            .I(\U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_0_0_a2Z0Z_1 ));
    CascadeMux I__453 (
            .O(N__4365),
            .I(\U409_AUTOCONFIG.N_405_cascade_ ));
    InMux I__452 (
            .O(N__4362),
            .I(N__4354));
    InMux I__451 (
            .O(N__4361),
            .I(N__4354));
    InMux I__450 (
            .O(N__4360),
            .I(N__4351));
    CascadeMux I__449 (
            .O(N__4359),
            .I(N__4348));
    LocalMux I__448 (
            .O(N__4354),
            .I(N__4345));
    LocalMux I__447 (
            .O(N__4351),
            .I(N__4342));
    InMux I__446 (
            .O(N__4348),
            .I(N__4339));
    Odrv4 I__445 (
            .O(N__4345),
            .I(\U409_AUTOCONFIG.N_414 ));
    Odrv4 I__444 (
            .O(N__4342),
            .I(\U409_AUTOCONFIG.N_414 ));
    LocalMux I__443 (
            .O(N__4339),
            .I(\U409_AUTOCONFIG.N_414 ));
    InMux I__442 (
            .O(N__4332),
            .I(N__4328));
    InMux I__441 (
            .O(N__4331),
            .I(N__4325));
    LocalMux I__440 (
            .O(N__4328),
            .I(\U409_AUTOCONFIG.N_373 ));
    LocalMux I__439 (
            .O(N__4325),
            .I(\U409_AUTOCONFIG.N_373 ));
    CascadeMux I__438 (
            .O(N__4320),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_2_3_0_cascade_ ));
    InMux I__437 (
            .O(N__4317),
            .I(N__4314));
    LocalMux I__436 (
            .O(N__4314),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_0_0 ));
    InMux I__435 (
            .O(N__4311),
            .I(N__4305));
    InMux I__434 (
            .O(N__4310),
            .I(N__4305));
    LocalMux I__433 (
            .O(N__4305),
            .I(\U409_AUTOCONFIG.N_269 ));
    InMux I__432 (
            .O(N__4302),
            .I(N__4299));
    LocalMux I__431 (
            .O(N__4299),
            .I(N__4295));
    InMux I__430 (
            .O(N__4298),
            .I(N__4292));
    Odrv4 I__429 (
            .O(N__4295),
            .I(\U409_AUTOCONFIG.N_370 ));
    LocalMux I__428 (
            .O(N__4292),
            .I(\U409_AUTOCONFIG.N_370 ));
    CascadeMux I__427 (
            .O(N__4287),
            .I(\U409_AUTOCONFIG.N_195_cascade_ ));
    InMux I__426 (
            .O(N__4284),
            .I(N__4281));
    LocalMux I__425 (
            .O(N__4281),
            .I(N__4277));
    InMux I__424 (
            .O(N__4280),
            .I(N__4274));
    Odrv4 I__423 (
            .O(N__4277),
            .I(\U409_AUTOCONFIG.N_383 ));
    LocalMux I__422 (
            .O(N__4274),
            .I(\U409_AUTOCONFIG.N_383 ));
    CascadeMux I__421 (
            .O(N__4269),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_8_cascade_ ));
    InMux I__420 (
            .O(N__4266),
            .I(N__4262));
    InMux I__419 (
            .O(N__4265),
            .I(N__4259));
    LocalMux I__418 (
            .O(N__4262),
            .I(N__4254));
    LocalMux I__417 (
            .O(N__4259),
            .I(N__4254));
    Span4Mux_v I__416 (
            .O(N__4254),
            .I(N__4251));
    Span4Mux_v I__415 (
            .O(N__4251),
            .I(N__4248));
    Span4Mux_h I__414 (
            .O(N__4248),
            .I(N__4245));
    Odrv4 I__413 (
            .O(N__4245),
            .I(A_c_24));
    CascadeMux I__412 (
            .O(N__4242),
            .I(N__4239));
    InMux I__411 (
            .O(N__4239),
            .I(N__4236));
    LocalMux I__410 (
            .O(N__4236),
            .I(\U409_AUTOCONFIG.N_270 ));
    InMux I__409 (
            .O(N__4233),
            .I(N__4230));
    LocalMux I__408 (
            .O(N__4230),
            .I(\U409_AUTOCONFIG.N_271 ));
    CascadeMux I__407 (
            .O(N__4227),
            .I(\U409_AUTOCONFIG.N_433_cascade_ ));
    InMux I__406 (
            .O(N__4224),
            .I(N__4221));
    LocalMux I__405 (
            .O(N__4221),
            .I(\U409_AUTOCONFIG.N_433 ));
    CascadeMux I__404 (
            .O(N__4218),
            .I(N__4215));
    InMux I__403 (
            .O(N__4215),
            .I(N__4209));
    InMux I__402 (
            .O(N__4214),
            .I(N__4209));
    LocalMux I__401 (
            .O(N__4209),
            .I(N__4206));
    Span4Mux_v I__400 (
            .O(N__4206),
            .I(N__4203));
    Sp12to4 I__399 (
            .O(N__4203),
            .I(N__4200));
    Odrv12 I__398 (
            .O(N__4200),
            .I(A_c_25));
    InMux I__397 (
            .O(N__4197),
            .I(N__4191));
    InMux I__396 (
            .O(N__4196),
            .I(N__4191));
    LocalMux I__395 (
            .O(N__4191),
            .I(N__4188));
    Span4Mux_v I__394 (
            .O(N__4188),
            .I(N__4185));
    Span4Mux_h I__393 (
            .O(N__4185),
            .I(N__4182));
    Odrv4 I__392 (
            .O(N__4182),
            .I(A_c_27));
    CascadeMux I__391 (
            .O(N__4179),
            .I(N__4175));
    InMux I__390 (
            .O(N__4178),
            .I(N__4170));
    InMux I__389 (
            .O(N__4175),
            .I(N__4170));
    LocalMux I__388 (
            .O(N__4170),
            .I(N__4167));
    Span4Mux_v I__387 (
            .O(N__4167),
            .I(N__4164));
    Span4Mux_v I__386 (
            .O(N__4164),
            .I(N__4161));
    Sp12to4 I__385 (
            .O(N__4161),
            .I(N__4158));
    Odrv12 I__384 (
            .O(N__4158),
            .I(A_c_26));
    IoInMux I__383 (
            .O(N__4155),
            .I(N__4152));
    LocalMux I__382 (
            .O(N__4152),
            .I(N__4149));
    Span4Mux_s2_h I__381 (
            .O(N__4149),
            .I(N__4146));
    Sp12to4 I__380 (
            .O(N__4146),
            .I(N__4143));
    Span12Mux_v I__379 (
            .O(N__4143),
            .I(N__4140));
    Span12Mux_v I__378 (
            .O(N__4140),
            .I(N__4137));
    Odrv12 I__377 (
            .O(N__4137),
            .I(PIO_P0_c));
    IoInMux I__376 (
            .O(N__4134),
            .I(N__4131));
    LocalMux I__375 (
            .O(N__4131),
            .I(N__4128));
    IoSpan4Mux I__374 (
            .O(N__4128),
            .I(N__4125));
    Span4Mux_s2_h I__373 (
            .O(N__4125),
            .I(N__4122));
    Sp12to4 I__372 (
            .O(N__4122),
            .I(N__4119));
    Span12Mux_v I__371 (
            .O(N__4119),
            .I(N__4116));
    Span12Mux_v I__370 (
            .O(N__4116),
            .I(N__4113));
    Odrv12 I__369 (
            .O(N__4113),
            .I(PIO_S0_c));
    ClkMux I__368 (
            .O(N__4110),
            .I(N__4077));
    ClkMux I__367 (
            .O(N__4109),
            .I(N__4077));
    ClkMux I__366 (
            .O(N__4108),
            .I(N__4077));
    ClkMux I__365 (
            .O(N__4107),
            .I(N__4077));
    ClkMux I__364 (
            .O(N__4106),
            .I(N__4077));
    ClkMux I__363 (
            .O(N__4105),
            .I(N__4077));
    ClkMux I__362 (
            .O(N__4104),
            .I(N__4077));
    ClkMux I__361 (
            .O(N__4103),
            .I(N__4077));
    ClkMux I__360 (
            .O(N__4102),
            .I(N__4077));
    ClkMux I__359 (
            .O(N__4101),
            .I(N__4077));
    ClkMux I__358 (
            .O(N__4100),
            .I(N__4077));
    GlobalMux I__357 (
            .O(N__4077),
            .I(CLK80_OUT));
    INV \INVU409_TRANSFER_ACK.CIA_ENABLED_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .I(N__4101));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .I(N__4100));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .I(N__4107));
    INV \INVU409_TRANSFER_ACK.TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.TACK_ENC_net ),
            .I(N__4104));
    INV \INVU409_TRANSFER_ACK.TACK_OUTnC  (
            .O(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .I(N__4102));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net ),
            .I(N__4106));
    INV \INVU409_AUTOCONFIG.CONFIGENnC  (
            .O(\INVU409_AUTOCONFIG.CONFIGENnC_net ),
            .I(N__8329));
    INV \INVU409_TRANSFER_ACK.CIA_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .I(N__4103));
    INV \INVU409_AUTOCONFIG.ATA_BASE_ness_3C  (
            .O(\INVU409_AUTOCONFIG.ATA_BASE_ness_3C_net ),
            .I(N__8344));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .I(N__4108));
    INV \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC  (
            .O(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .I(N__4105));
    INV \INVU409_AUTOCONFIG.ATA_BASE_ness_4C  (
            .O(\INVU409_AUTOCONFIG.ATA_BASE_ness_4C_net ),
            .I(N__8346));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net ),
            .I(N__4110));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .I(N__4109));
    INV \INVU409_AUTOCONFIG.AC_TACKC  (
            .O(\INVU409_AUTOCONFIG.AC_TACKC_net ),
            .I(N__8342));
    INV \INVU409_AUTOCONFIG.BRIDGE_BASE_3C  (
            .O(\INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net ),
            .I(N__8349));
    INV \INVU409_AUTOCONFIG.STATE_0C  (
            .O(\INVU409_AUTOCONFIG.STATE_0C_net ),
            .I(N__8345));
    INV \INVU409_AUTOCONFIG.LIDE_OUT_0C  (
            .O(\INVU409_AUTOCONFIG.LIDE_OUT_0C_net ),
            .I(N__8347));
    INV \INVU409_AUTOCONFIG.BRIDGE_OUT_3C  (
            .O(\INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net ),
            .I(N__8350));
    defparam IN_MUX_bfv_13_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_6_0_));
    defparam IN_MUX_bfv_13_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_7_0_ (
            .carryinitin(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .carryinitout(bfn_13_7_0_));
    defparam IN_MUX_bfv_14_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_5_0_));
    defparam IN_MUX_bfv_14_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_6_0_ (
            .carryinitin(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .carryinitout(bfn_14_6_0_));
    defparam IN_MUX_bfv_14_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_9_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__9009),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_o2_4_LC_1_15_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_o2_4_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_o2_4_LC_1_15_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_o2_4_LC_1_15_1  (
            .in0(N__4214),
            .in1(N__4196),
            .in2(N__4179),
            .in3(N__4265),
            .lcout(U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_o2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_8_LC_1_15_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_8_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_8_LC_1_15_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_8_LC_1_15_5  (
            .in0(N__5684),
            .in1(N__5614),
            .in2(N__4218),
            .in3(N__5397),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_11_LC_1_15_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_11_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_11_LC_1_15_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_11_LC_1_15_6  (
            .in0(N__4197),
            .in1(N__4178),
            .in2(N__4269),
            .in3(N__4266),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_5_9_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_5_9_0 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_5_9_0  (
            .in0(N__4233),
            .in1(N__9169),
            .in2(N__4242),
            .in3(N__4317),
            .lcout(\U409_AUTOCONFIG.N_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_5_9_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_5_9_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_5_9_1  (
            .in0(N__4725),
            .in1(N__4840),
            .in2(_gnd_net_),
            .in3(N__4360),
            .lcout(\U409_AUTOCONFIG.N_270 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_5_9_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_5_9_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_5_9_7  (
            .in0(N__4302),
            .in1(N__4332),
            .in2(N__4741),
            .in3(N__7280),
            .lcout(\U409_AUTOCONFIG.N_271 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_5_10_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_5_10_0 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_5_10_0  (
            .in0(N__4310),
            .in1(N__4834),
            .in2(N__4359),
            .in3(N__7329),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_5_0_LC_5_10_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_5_0_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_5_0_LC_5_10_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_5_0_LC_5_10_1  (
            .in0(N__4835),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5166),
            .lcout(\U409_AUTOCONFIG.N_373 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_0_71_i_i_0_a2_1_LC_5_10_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_0_71_i_i_0_a2_1_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_0_71_i_i_0_a2_1_LC_5_10_2 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_7_0_71_i_i_0_a2_1_LC_5_10_2  (
            .in0(N__5167),
            .in1(N__4836),
            .in2(N__4742),
            .in3(N__7331),
            .lcout(\U409_AUTOCONFIG.N_433 ),
            .ltout(\U409_AUTOCONFIG.N_433_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_2_LC_5_10_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_2_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_2_LC_5_10_3 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_2_LC_5_10_3  (
            .in0(N__4298),
            .in1(_gnd_net_),
            .in2(N__4227),
            .in3(N__4284),
            .lcout(\U409_AUTOCONFIG.N_285 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_5_10_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_5_10_4 .LUT_INIT=16'b1100110111001100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_5_10_4  (
            .in0(N__5248),
            .in1(N__4224),
            .in2(N__4743),
            .in3(N__7333),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTc_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_4_0_LC_5_10_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_4_0_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_4_0_LC_5_10_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_4_0_LC_5_10_5  (
            .in0(N__7330),
            .in1(N__4447),
            .in2(N__4740),
            .in3(N__5247),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_2_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_3_0_LC_5_10_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_3_0_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_3_0_LC_5_10_6 .LUT_INIT=16'b1010101011101010;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_3_0_LC_5_10_6  (
            .in0(N__4311),
            .in1(N__4331),
            .in2(N__4320),
            .in3(N__4512),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_5_10_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_5_10_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_5_10_7  (
            .in0(N__7332),
            .in1(N__4732),
            .in2(N__4842),
            .in3(N__5168),
            .lcout(\U409_AUTOCONFIG.N_286 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_0_LC_5_11_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_0_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_0_LC_5_11_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_0_LC_5_11_0  (
            .in0(N__4280),
            .in1(N__4464),
            .in2(N__5227),
            .in3(N__4492),
            .lcout(\U409_AUTOCONFIG.N_269 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_7_0_LC_5_11_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_7_0_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_7_0_LC_5_11_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_7_0_LC_5_11_2  (
            .in0(N__5154),
            .in1(N__4466),
            .in2(N__5228),
            .in3(N__4494),
            .lcout(\U409_AUTOCONFIG.N_414 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_4_0_LC_5_11_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_4_0_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_4_0_LC_5_11_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_4_0_LC_5_11_4  (
            .in0(N__5204),
            .in1(N__4465),
            .in2(_gnd_net_),
            .in3(N__4493),
            .lcout(\U409_AUTOCONFIG.N_370 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_0_0_o2_LC_5_11_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_0_0_o2_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_0_0_o2_LC_5_11_6 .LUT_INIT=16'b0000111111110001;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_0_0_o2_LC_5_11_6  (
            .in0(N__4809),
            .in1(N__7328),
            .in2(N__5229),
            .in3(N__4721),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.N_195_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_0_0_a2_1_LC_5_11_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_0_0_a2_1_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_0_0_a2_1_LC_5_11_7 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_0_0_a2_1_LC_5_11_7  (
            .in0(N__4467),
            .in1(_gnd_net_),
            .in2(N__4287),
            .in3(N__4504),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_0_0_a2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_5_12_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_5_12_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_5_12_1  (
            .in0(N__7327),
            .in1(N__4817),
            .in2(N__4692),
            .in3(N__5152),
            .lcout(\U409_AUTOCONFIG.N_274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_6_0_LC_5_12_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_6_0_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_6_0_LC_5_12_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_6_0_LC_5_12_5  (
            .in0(N__7326),
            .in1(N__4816),
            .in2(_gnd_net_),
            .in3(N__4672),
            .lcout(\U409_AUTOCONFIG.N_383 ),
            .ltout(\U409_AUTOCONFIG.N_383_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_5_12_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_5_12_6 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_5_12_6  (
            .in0(N__5151),
            .in1(N__4428),
            .in2(N__4422),
            .in3(N__5249),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTc_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_4_LC_5_14_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_4_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_4_LC_5_14_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_4_LC_5_14_2  (
            .in0(N__6723),
            .in1(N__6921),
            .in2(N__7700),
            .in3(N__7804),
            .lcout(\U409_ADDRESS_DECODE.N_344 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_2_LC_5_14_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_2_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_2_LC_5_14_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_2_LC_5_14_6  (
            .in0(N__6722),
            .in1(N__6920),
            .in2(N__7699),
            .in3(N__6117),
            .lcout(\U409_ADDRESS_DECODE.N_345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_10_LC_5_15_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_10_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_10_LC_5_15_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_10_LC_5_15_0  (
            .in0(N__4419),
            .in1(N__4404),
            .in2(N__9177),
            .in3(N__6615),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_1_LC_5_15_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_1_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_1_LC_5_15_4 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_1_LC_5_15_4  (
            .in0(N__7937),
            .in1(N__5067),
            .in2(N__4392),
            .in3(N__4383),
            .lcout(N_434),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_6_9_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_6_9_1 .LUT_INIT=16'b1000000000100000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_6_9_1  (
            .in0(N__4362),
            .in1(N__4841),
            .in2(N__7325),
            .in3(N__4739),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.N_288_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_6_9_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_6_9_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_6_9_2 .LUT_INIT=16'b0100110000001000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_6_9_2  (
            .in0(N__4575),
            .in1(N__9170),
            .in2(N__4377),
            .in3(N__5918),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_START_RNIJJLA1_LC_6_9_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_START_RNIJJLA1_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.AC_START_RNIJJLA1_LC_6_9_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_AUTOCONFIG.AC_START_RNIJJLA1_LC_6_9_3  (
            .in0(N__7121),
            .in1(N__5556),
            .in2(N__4902),
            .in3(N__4877),
            .lcout(\U409_AUTOCONFIG.N_405 ),
            .ltout(\U409_AUTOCONFIG.N_405_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_START_RNI3D7V2_LC_6_9_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_START_RNI3D7V2_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.AC_START_RNI3D7V2_LC_6_9_4 .LUT_INIT=16'b1111010111010101;
    LogicCell40 \U409_AUTOCONFIG.AC_START_RNI3D7V2_LC_6_9_4  (
            .in0(N__9163),
            .in1(N__4374),
            .in2(N__4365),
            .in3(N__4361),
            .lcout(\U409_AUTOCONFIG.AC_START_RNI3D7VZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_6_9_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_6_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_6_9_5 .LUT_INIT=16'b0100010011000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_6_9_5  (
            .in0(N__4593),
            .in1(N__9168),
            .in2(N__6410),
            .in3(N__4574),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_6_9_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_6_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_6_9_6 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_6_9_6  (
            .in0(N__4573),
            .in1(N__4587),
            .in2(N__9178),
            .in3(N__4952),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_6_9_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_6_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_6_9_7 .LUT_INIT=16'b0100010011000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_6_9_7  (
            .in0(N__4581),
            .in1(N__9167),
            .in2(N__5525),
            .in3(N__4572),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_6_10_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_6_10_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_6_10_1 .LUT_INIT=16'b0000010111001100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_0_LC_6_10_1  (
            .in0(N__4560),
            .in1(N__4934),
            .in2(N__5103),
            .in3(N__4530),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_0C_net ),
            .ce(),
            .sr(N__9424));
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_6_10_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_6_10_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_6_10_2 .LUT_INIT=16'b0101011100000010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_1_LC_6_10_2  (
            .in0(N__4531),
            .in1(N__4863),
            .in2(N__4551),
            .in3(N__5498),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_0C_net ),
            .ce(),
            .sr(N__9424));
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_6_10_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_6_10_3 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_6_10_3 .LUT_INIT=16'b0000010111001100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_2_LC_6_10_3  (
            .in0(N__4539),
            .in1(N__6389),
            .in2(N__4854),
            .in3(N__4532),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_0C_net ),
            .ce(),
            .sr(N__9424));
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_6_10_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_6_10_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_6_10_4 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_3_LC_6_10_4  (
            .in0(N__4533),
            .in1(N__4518),
            .in2(N__5942),
            .in3(N__4853),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_0C_net ),
            .ce(),
            .sr(N__9424));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_6_11_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_6_11_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_6_11_2  (
            .in0(N__4737),
            .in1(N__4811),
            .in2(N__7363),
            .in3(N__5165),
            .lcout(\U409_AUTOCONFIG.N_287 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_STATE_1_0_a2_0_2_LC_6_11_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_STATE_1_0_a2_0_2_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_STATE_1_0_a2_0_2_LC_6_11_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_AUTOCONFIG.un1_STATE_1_0_a2_0_2_LC_6_11_3  (
            .in0(N__5232),
            .in1(N__5262),
            .in2(N__4511),
            .in3(N__4463),
            .lcout(\U409_AUTOCONFIG.un1_STATE_1_0_a2_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_6_11_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_6_11_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_6_11_4  (
            .in0(N__4736),
            .in1(N__4810),
            .in2(N__7362),
            .in3(N__5230),
            .lcout(\U409_AUTOCONFIG.N_273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_1_129_i_i_0_a2_0_LC_6_11_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_1_129_i_i_0_a2_0_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_1_129_i_i_0_a2_0_LC_6_11_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_1_129_i_i_0_a2_0_LC_6_11_6  (
            .in0(N__4738),
            .in1(N__4812),
            .in2(N__7364),
            .in3(N__5231),
            .lcout(\U409_AUTOCONFIG.N_400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_2_LC_6_12_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_2_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_2_LC_6_12_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_2_LC_6_12_5  (
            .in0(N__6112),
            .in1(N__6893),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_374),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_3_0_LC_6_12_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_3_0_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_3_0_LC_6_12_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_3_0_LC_6_12_6  (
            .in0(_gnd_net_),
            .in1(N__4830),
            .in2(_gnd_net_),
            .in3(N__4676),
            .lcout(\U409_AUTOCONFIG.N_360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_9_LC_6_14_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_9_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_9_LC_6_14_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_9_LC_6_14_0  (
            .in0(N__6699),
            .in1(N__7839),
            .in2(N__5451),
            .in3(N__4616),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_6_14_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_6_14_1 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_6_14_1  (
            .in0(N__4641),
            .in1(N__4635),
            .in2(N__4620),
            .in3(N__4599),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_i_a2_1_LC_6_14_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_i_a2_1_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_i_a2_1_LC_6_14_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_i_a2_1_LC_6_14_5  (
            .in0(N__5018),
            .in1(N__5054),
            .in2(N__4617),
            .in3(N__9270),
            .lcout(N_401),
            .ltout(N_401_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_6_14_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_6_14_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_6_14_6  (
            .in0(N__6698),
            .in1(N__6735),
            .in2(N__4602),
            .in3(N__6590),
            .lcout(N_436),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_0_LC_6_15_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_0_LC_6_15_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_0_LC_6_15_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_0_LC_6_15_2  (
            .in0(N__9159),
            .in1(N__5538),
            .in2(_gnd_net_),
            .in3(N__4972),
            .lcout(N_348),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.N_265_i_LC_6_15_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.N_265_i_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.N_265_i_LC_6_15_3 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \U409_ADDRESS_DECODE.N_265_i_LC_6_15_3  (
            .in0(N__5536),
            .in1(N__9158),
            .in2(N__4973),
            .in3(N__6842),
            .lcout(N_265_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_0_LC_6_15_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_0_LC_6_15_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_0_LC_6_15_7 .LUT_INIT=16'b1111111011111011;
    LogicCell40 \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_0_LC_6_15_7  (
            .in0(N__5537),
            .in1(N__5011),
            .in2(N__4974),
            .in3(N__5042),
            .lcout(\U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIMM061_0_LC_7_8_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIMM061_0_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIMM061_0_LC_7_8_1 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNIMM061_0_LC_7_8_1  (
            .in0(N__4953),
            .in1(N__6376),
            .in2(N__4941),
            .in3(N__7471),
            .lcout(N_124),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_START_LC_7_9_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_START_LC_7_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.AC_START_LC_7_9_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U409_AUTOCONFIG.AC_START_LC_7_9_7  (
            .in0(N__8438),
            .in1(N__6318),
            .in2(_gnd_net_),
            .in3(N__7201),
            .lcout(\U409_AUTOCONFIG.AC_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8348),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNI2IAK1_0_LC_7_10_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNI2IAK1_0_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNI2IAK1_0_LC_7_10_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNI2IAK1_0_LC_7_10_0  (
            .in0(N__5172),
            .in1(N__7140),
            .in2(N__4911),
            .in3(N__5557),
            .lcout(\U409_AUTOCONFIG.un1_STATE_1_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_0_LC_7_10_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_0_LC_7_10_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.STATE_0_LC_7_10_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_AUTOCONFIG.STATE_0_LC_7_10_1  (
            .in0(N__5558),
            .in1(N__4895),
            .in2(N__9179),
            .in3(N__4878),
            .lcout(\U409_AUTOCONFIG.STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_5_LC_7_10_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_5_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_5_LC_7_10_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_5_LC_7_10_2  (
            .in0(N__6932),
            .in1(N__6775),
            .in2(_gnd_net_),
            .in3(N__6088),
            .lcout(),
            .ltout(N_354_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_a2_1_LC_7_10_3 .C_ON=1'b0;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_a2_1_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_a2_1_LC_7_10_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_DATA_BUFFERS.un1_BUFENn_i_a2_1_LC_7_10_3  (
            .in0(N__9230),
            .in1(N__6448),
            .in2(N__4866),
            .in3(N__9308),
            .lcout(N_356),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_1_LC_7_10_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_1_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_1_LC_7_10_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_1_LC_7_10_7  (
            .in0(N__7787),
            .in1(N__7936),
            .in2(_gnd_net_),
            .in3(N__7718),
            .lcout(N_351),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_7_11_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_7_11_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.D_1_i_LC_7_11_0  (
            .in0(N__6661),
            .in1(N__7135),
            .in2(N__6606),
            .in3(N__7059),
            .lcout(D_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_1_i_a2_LC_7_11_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_1_i_a2_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_1_i_a2_LC_7_11_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_1_i_a2_LC_7_11_2  (
            .in0(N__6662),
            .in1(N__6586),
            .in2(_gnd_net_),
            .in3(N__7060),
            .lcout(N_357),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_a2_0_LC_7_12_2 .C_ON=1'b0;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_a2_0_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_a2_0_LC_7_12_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_DATA_BUFFERS.un1_BUFENn_i_a2_0_LC_7_12_2  (
            .in0(N__7962),
            .in1(N__7802),
            .in2(N__6607),
            .in3(N__7067),
            .lcout(N_297),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_7_12_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_7_12_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_7_12_7  (
            .in0(N__5286),
            .in1(N__5261),
            .in2(N__5250),
            .in3(N__5153),
            .lcout(\U409_AUTOCONFIG.N_276 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_7_13_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_7_13_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(N__6006),
            .in2(_gnd_net_),
            .in3(N__5974),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_i_1_LC_7_14_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_i_1_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_i_1_LC_7_14_2 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_i_1_LC_7_14_2  (
            .in0(N__6736),
            .in1(N__7857),
            .in2(N__6694),
            .in3(N__8417),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.PORTSIZE_iZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_i_LC_7_14_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_i_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_i_LC_7_14_3 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_i_LC_7_14_3  (
            .in0(N__6854),
            .in1(N__9271),
            .in2(N__5088),
            .in3(N__8039),
            .lcout(N_139),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_3_LC_7_14_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_3_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_3_LC_7_14_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_3_LC_7_14_5  (
            .in0(N__6116),
            .in1(N__6737),
            .in2(N__6931),
            .in3(N__6519),
            .lcout(\U409_ADDRESS_DECODE.N_343 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_x2_LC_7_15_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_x2_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_x2_LC_7_15_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_x2_LC_7_15_5  (
            .in0(N__5055),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5019),
            .lcout(N_156_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_o2_5_LC_7_15_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_o2_5_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_o2_5_LC_7_15_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_o2_5_LC_7_15_6  (
            .in0(N__5691),
            .in1(N__5625),
            .in2(N__5395),
            .in3(N__5447),
            .lcout(U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_o2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIOO061_1_LC_8_7_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIOO061_1_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIOO061_1_LC_8_7_2 .LUT_INIT=16'b1111101011001100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNIOO061_1_LC_8_7_2  (
            .in0(N__5526),
            .in1(N__5505),
            .in2(N__6378),
            .in3(N__7470),
            .lcout(N_126),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_8_8_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_8_8_1 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_8_8_1 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_8_8_1  (
            .in0(N__7646),
            .in1(N__5651),
            .in2(N__7578),
            .in3(N__5574),
            .lcout(BRIDGE_BASE_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net ),
            .ce(),
            .sr(N__9425));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_8_8_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_8_8_2 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_8_8_2 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_8_8_2  (
            .in0(N__5572),
            .in1(N__7644),
            .in2(N__5822),
            .in3(N__5408),
            .lcout(BRIDGE_BASE_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net ),
            .ce(),
            .sr(N__9425));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_8_8_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_8_8_3 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_8_8_3 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_8_8_3  (
            .in0(N__7643),
            .in1(N__5345),
            .in2(N__5871),
            .in3(N__5571),
            .lcout(BRIDGE_BASE_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net ),
            .ce(),
            .sr(N__9425));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_8_8_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_8_8_5 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_8_8_5 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_8_8_5  (
            .in0(N__7645),
            .in1(N__5636),
            .in2(N__6191),
            .in3(N__5573),
            .lcout(BRIDGE_BASE_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net ),
            .ce(),
            .sr(N__9425));
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0_LC_8_9_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0_LC_8_9_0 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0_LC_8_9_0  (
            .in0(N__5334),
            .in1(N__5580),
            .in2(N__6495),
            .in3(N__9247),
            .lcout(N_96),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0_0_LC_8_9_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0_0_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0_0_LC_8_9_1 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0_0_LC_8_9_1  (
            .in0(N__5446),
            .in1(N__5409),
            .in2(N__5396),
            .in3(N__5346),
            .lcout(\U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIOE6K2_LC_8_9_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIOE6K2_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIOE6K2_LC_8_9_2 .LUT_INIT=16'b1100111011101110;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNIOE6K2_LC_8_9_2  (
            .in0(N__7392),
            .in1(N__9429),
            .in2(N__7464),
            .in3(N__7285),
            .lcout(\U409_AUTOCONFIG.un1_STATE_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0_1_LC_8_9_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0_1_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0_1_LC_8_9_4 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0_1_LC_8_9_4  (
            .in0(N__5683),
            .in1(N__5652),
            .in2(N__5640),
            .in3(N__5624),
            .lcout(\U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI25A42_LC_8_9_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI25A42_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI25A42_LC_8_9_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNI25A42_LC_8_9_5  (
            .in0(N__7284),
            .in1(N__7443),
            .in2(_gnd_net_),
            .in3(N__7391),
            .lcout(\U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_o2dup_LC_8_9_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_o2dup_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_o2dup_LC_8_9_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_o2dup_LC_8_9_7  (
            .in0(N__9136),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7202),
            .lcout(\U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_o2dupZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_TACK_LC_8_10_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_TACK_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.AC_TACK_LC_8_10_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \U409_AUTOCONFIG.AC_TACK_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__5559),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(AC_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.AC_TACKC_net ),
            .ce(),
            .sr(N__9418));
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_LC_8_10_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_LC_8_10_3 .LUT_INIT=16'b1010111010101010;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_CONF_LC_8_10_3  (
            .in0(N__6362),
            .in1(N__7393),
            .in2(N__7365),
            .in3(N__7451),
            .lcout(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.AC_TACKC_net ),
            .ce(),
            .sr(N__9418));
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_8_10_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_8_10_7 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_LC_8_10_7  (
            .in0(N__7346),
            .in1(N__7394),
            .in2(_gnd_net_),
            .in3(N__7450),
            .lcout(\U409_AUTOCONFIG.LIDE_CONFZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.AC_TACKC_net ),
            .ce(),
            .sr(N__9418));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_8_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_8_11_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_8_11_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_8_11_0  (
            .in0(N__7041),
            .in1(N__7008),
            .in2(_gnd_net_),
            .in3(N__6987),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__6810));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_8_11_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_8_11_5 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_8_11_5 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_8_11_5  (
            .in0(N__5771),
            .in1(N__5790),
            .in2(N__5745),
            .in3(N__6262),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__6810));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_8_11_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_8_11_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_8_11_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_8_11_7  (
            .in0(N__5741),
            .in1(N__5789),
            .in2(_gnd_net_),
            .in3(N__6261),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__6810));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_8_12_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_8_12_0 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_8_12_0  (
            .in0(N__7035),
            .in1(N__6001),
            .in2(N__5733),
            .in3(N__5796),
            .lcout(\U409_TRANSFER_ACK.N_237 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_8_12_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_8_12_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_8_12_1  (
            .in0(N__5969),
            .in1(N__5787),
            .in2(N__5714),
            .in3(N__5767),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_8_12_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_8_12_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_8_12_2  (
            .in0(N__5788),
            .in1(N__5970),
            .in2(N__5772),
            .in3(N__5706),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_8_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_8_12_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_8_12_3  (
            .in0(N__6002),
            .in1(N__7036),
            .in2(N__5754),
            .in3(N__5732),
            .lcout(\U409_TRANSFER_ACK.N_268 ),
            .ltout(\U409_TRANSFER_ACK.N_268_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_3_LC_8_12_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_3_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_3_LC_8_12_4 .LUT_INIT=16'b0010000011111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_3_LC_8_12_4  (
            .in0(N__8380),
            .in1(N__6306),
            .in2(N__5751),
            .in3(N__6221),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_8_12_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_8_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_8_12_5  (
            .in0(N__7006),
            .in1(N__6011),
            .in2(N__5715),
            .in3(N__5976),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_8_12_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_8_12_6 .LUT_INIT=16'b1000000010000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_8_12_6  (
            .in0(N__7037),
            .in1(N__6984),
            .in2(N__5748),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_8_12_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_8_12_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_8_12_7  (
            .in0(N__7005),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6983),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_8_13_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_8_13_5 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_8_13_5 .LUT_INIT=16'b0000000001011010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_8_13_5  (
            .in0(N__6952),
            .in1(_gnd_net_),
            .in2(N__6012),
            .in3(N__6256),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net ),
            .ce(),
            .sr(N__6808));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_8_13_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_8_13_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_8_13_6 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_8_13_6  (
            .in0(N__6956),
            .in1(N__5721),
            .in2(N__6264),
            .in3(N__5713),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net ),
            .ce(),
            .sr(N__6808));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_8_13_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_8_13_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_8_13_7 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_8_13_7  (
            .in0(N__6007),
            .in1(N__5975),
            .in2(N__6957),
            .in3(N__6260),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net ),
            .ce(),
            .sr(N__6808));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_i_a2_0_LC_8_14_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_i_a2_0_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_i_a2_0_LC_8_14_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_i_a2_0_LC_8_14_2  (
            .in0(N__7952),
            .in1(N__6515),
            .in2(N__7874),
            .in3(N__7835),
            .lcout(N_339),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNISS061_3_LC_9_7_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNISS061_3_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNISS061_3_LC_9_7_4 .LUT_INIT=16'b1111101011001010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNISS061_3_LC_9_7_4  (
            .in0(N__5946),
            .in1(N__5925),
            .in2(N__7479),
            .in3(N__6377),
            .lcout(N_130),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_2_LC_9_8_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_2_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_2_LC_9_8_0 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_2_LC_9_8_0  (
            .in0(N__6783),
            .in1(N__5879),
            .in2(N__6939),
            .in3(N__5888),
            .lcout(\U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_4_LC_9_8_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_4_LC_9_8_1 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_4_LC_9_8_1 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_ness_4_LC_9_8_1  (
            .in0(N__5889),
            .in1(N__5870),
            .in2(N__7639),
            .in3(N__7491),
            .lcout(ATA_BASE_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_ness_4C_net ),
            .ce(N__7505),
            .sr(N__9420));
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_5_LC_9_8_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_5_LC_9_8_2 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_5_LC_9_8_2 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_ness_5_LC_9_8_2  (
            .in0(N__7492),
            .in1(N__7623),
            .in2(N__5835),
            .in3(N__5880),
            .lcout(ATA_BASE_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_ness_4C_net ),
            .ce(N__7505),
            .sr(N__9420));
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_0_LC_9_8_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_0_LC_9_8_3 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_0_LC_9_8_3 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_ness_0_LC_9_8_3  (
            .in0(N__7367),
            .in1(N__5869),
            .in2(N__7638),
            .in3(N__6138),
            .lcout(ATA_BASE_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_ness_4C_net ),
            .ce(N__7505),
            .sr(N__9420));
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_1_LC_9_8_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_1_LC_9_8_4 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_1_LC_9_8_4 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_ness_1_LC_9_8_4  (
            .in0(N__5831),
            .in1(N__7368),
            .in2(N__6153),
            .in3(N__7618),
            .lcout(ATA_BASE_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_ness_4C_net ),
            .ce(N__7505),
            .sr(N__9420));
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_6_LC_9_8_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_6_LC_9_8_5 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_6_LC_9_8_5 .LUT_INIT=16'b1110110000100000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_ness_6_LC_9_8_5  (
            .in0(N__7624),
            .in1(N__7493),
            .in2(N__6210),
            .in3(N__6165),
            .lcout(ATA_BASE_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_ness_4C_net ),
            .ce(N__7505),
            .sr(N__9420));
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_2_LC_9_8_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_2_LC_9_8_6 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_2_LC_9_8_6 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_ness_2_LC_9_8_6  (
            .in0(N__6063),
            .in1(N__7619),
            .in2(N__6209),
            .in3(N__7369),
            .lcout(ATA_BASE_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_ness_4C_net ),
            .ce(N__7505),
            .sr(N__9420));
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_7_LC_9_8_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_7_LC_9_8_7 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_7_LC_9_8_7 .LUT_INIT=16'b1110110000100000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_ness_7_LC_9_8_7  (
            .in0(N__7625),
            .in1(N__7494),
            .in2(N__7577),
            .in3(N__7737),
            .lcout(ATA_BASE_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_ness_4C_net ),
            .ce(N__7505),
            .sr(N__9420));
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_7_0_LC_9_9_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_7_0_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_7_0_LC_9_9_0 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_7_0_LC_9_9_0  (
            .in0(N__7968),
            .in1(N__6164),
            .in2(N__6608),
            .in3(N__6149),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_7Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_7_LC_9_9_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_7_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_7_LC_9_9_1 .LUT_INIT=16'b1111111111110110;
    LogicCell40 \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_7_LC_9_9_1  (
            .in0(N__6455),
            .in1(N__6137),
            .in2(N__6126),
            .in3(N__6051),
            .lcout(\U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_7 ),
            .ltout(\U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNO_1_LC_9_9_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNO_1_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNO_1_LC_9_9_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_RNO_1_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6123),
            .in3(N__7655),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.ATA_EN_2_0_o2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_LC_9_9_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_LC_9_9_3 .LUT_INIT=16'b1000100010001010;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_LC_9_9_3  (
            .in0(N__9135),
            .in1(N__6476),
            .in2(N__6120),
            .in3(N__6045),
            .lcout(\U409_ADDRESS_DECODE.ATA_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8343),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_x2_LC_9_9_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_x2_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_x2_LC_9_9_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_ADDRESS_DECODE.un1_ATA_ENn_i_x2_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__6111),
            .in2(_gnd_net_),
            .in3(N__6062),
            .lcout(\U409_ADDRESS_DECODE.N_183_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNO_0_LC_9_9_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNO_0_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNO_0_LC_9_9_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_RNO_0_LC_9_9_5  (
            .in0(N__6029),
            .in1(N__6038),
            .in2(N__7134),
            .in3(N__7182),
            .lcout(\U409_ADDRESS_DECODE.ATA_EN_2_0_o2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_0_3_LC_9_9_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_0_3_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_0_3_LC_9_9_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U409_ADDRESS_DECODE.un1_ATA_ENn_i_0_3_LC_9_9_6  (
            .in0(N__6039),
            .in1(N__6030),
            .in2(N__6504),
            .in3(N__6494),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.un1_ATA_ENn_i_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNIU5437_LC_9_9_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNIU5437_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNIU5437_LC_9_9_7 .LUT_INIT=16'b1111101011111111;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_RNIU5437_LC_9_9_7  (
            .in0(N__7656),
            .in1(_gnd_net_),
            .in2(N__6480),
            .in3(N__6477),
            .lcout(N_107),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_3_LC_9_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_3_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_3_LC_9_10_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_3_LC_9_10_0  (
            .in0(N__6782),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6456),
            .lcout(N_422),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_3_LC_9_10_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_3_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_3_LC_9_10_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_3_LC_9_10_1  (
            .in0(N__6321),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8382),
            .lcout(\U409_TRANSFER_ACK.N_381 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_9_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_9_10_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_9_10_5  (
            .in0(N__6320),
            .in1(N__8381),
            .in2(N__8129),
            .in3(N__8144),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIQQ061_2_LC_9_10_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIQQ061_2_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIQQ061_2_LC_9_10_6 .LUT_INIT=16'b1111110010101100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNIQQ061_2_LC_9_10_6  (
            .in0(N__6414),
            .in1(N__6393),
            .in2(N__7469),
            .in3(N__6363),
            .lcout(N_128),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_9_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_9_11_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_9_11_0 .LUT_INIT=16'b1101110000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_9_11_0  (
            .in0(N__6319),
            .in1(N__7040),
            .in2(N__8385),
            .in3(N__6233),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__6809));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_9_11_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_9_11_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_9_11_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_9_11_1  (
            .in0(N__7039),
            .in1(N__6986),
            .in2(_gnd_net_),
            .in3(N__6263),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__6809));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_9_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_9_11_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_9_11_2 .LUT_INIT=16'b0100010011111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_9_11_2  (
            .in0(N__6234),
            .in1(N__7161),
            .in2(_gnd_net_),
            .in3(N__6222),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__6809));
    defparam \U409_ADDRESS_DECODE.D_IN_0_a2_0_0_LC_9_12_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.D_IN_0_a2_0_0_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.D_IN_0_a2_0_0_LC_9_12_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.D_IN_0_a2_0_0_LC_9_12_2  (
            .in0(N__7139),
            .in1(N__6612),
            .in2(N__7074),
            .in3(N__6695),
            .lcout(N_361),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_9_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_9_12_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_9_12_3  (
            .in0(N__7038),
            .in1(N__7007),
            .in2(_gnd_net_),
            .in3(N__6985),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_LC_9_12_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_LC_9_12_4 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_LC_9_12_4  (
            .in0(N__9328),
            .in1(N__9380),
            .in2(N__6911),
            .in3(N__7811),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.N_346_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_9_12_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_9_12_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_9_12_5  (
            .in0(N__6900),
            .in1(N__6697),
            .in2(N__6861),
            .in3(N__6774),
            .lcout(\U409_TRANSFER_ACK.N_159 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a2_1_LC_9_12_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a2_1_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a2_1_LC_9_12_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a2_1_LC_9_12_7  (
            .in0(N__6764),
            .in1(N__7964),
            .in2(_gnd_net_),
            .in3(N__7711),
            .lcout(N_429),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_o2_LC_9_13_0 .C_ON=1'b0;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_o2_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_o2_LC_9_13_0 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \U409_DATA_BUFFERS.un1_BUFENn_i_o2_LC_9_13_0  (
            .in0(N__6858),
            .in1(N__9381),
            .in2(N__9335),
            .in3(N__9236),
            .lcout(N_190),
            .ltout(N_190_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_13_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_13_1 .LUT_INIT=16'b1011001111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_13_1  (
            .in0(N__9302),
            .in1(N__9180),
            .in2(N__6831),
            .in3(N__6828),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.N_436_i_LC_9_13_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.N_436_i_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.N_436_i_LC_9_13_3 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \U409_ADDRESS_DECODE.N_436_i_LC_9_13_3  (
            .in0(N__6763),
            .in1(N__6696),
            .in2(N__7881),
            .in3(N__6613),
            .lcout(N_436_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_i_a2_2_LC_9_14_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_i_a2_2_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_i_a2_2_LC_9_14_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_i_a2_2_LC_9_14_1  (
            .in0(N__7812),
            .in1(N__6614),
            .in2(_gnd_net_),
            .in3(N__7701),
            .lcout(N_431),
            .ltout(N_431_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_0_LC_9_14_2 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_0_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_0_LC_9_14_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_CIA.VMA_RNO_0_LC_9_14_2  (
            .in0(N__7963),
            .in1(N__7870),
            .in2(N__7842),
            .in3(N__7828),
            .lcout(\U409_CIA.VMA_3_0_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_5_LC_10_8_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_5_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_5_LC_10_8_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_5_LC_10_8_0  (
            .in0(N__7803),
            .in1(N__7736),
            .in2(N__7725),
            .in3(N__7523),
            .lcout(\U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_3_LC_10_8_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_3_LC_10_8_1 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.ATA_BASE_ness_3_LC_10_8_1 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_ness_3_LC_10_8_1  (
            .in0(N__7524),
            .in1(N__7370),
            .in2(N__7647),
            .in3(N__7558),
            .lcout(ATA_BASE_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_ness_3C_net ),
            .ce(N__7515),
            .sr(N__9419));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0JVF_LC_10_8_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0JVF_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0JVF_LC_10_8_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNI0JVF_LC_10_8_4  (
            .in0(N__7371),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7475),
            .lcout(\U409_AUTOCONFIG.N_172 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_9_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_9_2 .LUT_INIT=16'b0000110000101010;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_9_2  (
            .in0(N__8091),
            .in1(N__8916),
            .in2(N__8883),
            .in3(N__8268),
            .lcout(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__9417));
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_10_10_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_10_10_4 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_10_10_4 .LUT_INIT=16'b1111011100000000;
    LogicCell40 \U409_AUTOCONFIG.CONFIGENn_LC_10_10_4  (
            .in0(N__7468),
            .in1(N__7398),
            .in2(N__7366),
            .in3(N__7188),
            .lcout(CONFIGENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.CONFIGENnC_net ),
            .ce(),
            .sr(N__9416));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_10_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_10_10_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(N__7160),
            .in2(_gnd_net_),
            .in3(N__8105),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_10_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_10_10_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_10_10_6  (
            .in0(N__7149),
            .in1(N__8078),
            .in2(N__8094),
            .in3(N__8090),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_10_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_10_11_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_10_11_2 .LUT_INIT=16'b0111100011010000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_10_11_2  (
            .in0(N__8520),
            .in1(N__8551),
            .in2(N__8592),
            .in3(N__8632),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net ),
            .ce(),
            .sr(N__9414));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_10_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_10_11_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_10_11_6 .LUT_INIT=16'b1000101010111010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_LC_10_11_6  (
            .in0(N__8079),
            .in1(N__8552),
            .in2(N__8727),
            .in3(N__8633),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net ),
            .ce(),
            .sr(N__9414));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_1_0_LC_10_12_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_1_0_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_1_0_LC_10_12_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_1_0_LC_10_12_2  (
            .in0(N__8067),
            .in1(N__9304),
            .in2(N__8634),
            .in3(N__9246),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_10_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_10_12_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_10_12_3  (
            .in0(N__9303),
            .in1(N__8066),
            .in2(N__9249),
            .in3(N__8058),
            .lcout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_1_LC_10_12_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_1_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_1_LC_10_12_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_1_LC_10_12_4  (
            .in0(_gnd_net_),
            .in1(N__8545),
            .in2(_gnd_net_),
            .in3(N__8625),
            .lcout(\U409_TRANSFER_ACK.N_380 ),
            .ltout(\U409_TRANSFER_ACK.N_380_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_10_12_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_10_12_5 .LUT_INIT=16'b0000110011101110;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_10_12_5  (
            .in0(N__8702),
            .in1(N__8585),
            .in2(N__8052),
            .in3(N__8517),
            .lcout(\U409_TRANSFER_ACK.ROMENn_e_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_DATA_BUFFERS.N_94_i_LC_10_14_5 .C_ON=1'b0;
    defparam \U409_DATA_BUFFERS.N_94_i_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \U409_DATA_BUFFERS.N_94_i_LC_10_14_5 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \U409_DATA_BUFFERS.N_94_i_LC_10_14_5  (
            .in0(N__8049),
            .in1(N__9301),
            .in2(_gnd_net_),
            .in3(N__8043),
            .lcout(N_94_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_11_4_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_11_4_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_11_4_4 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_11_4_4  (
            .in0(_gnd_net_),
            .in1(N__8007),
            .in2(_gnd_net_),
            .in3(N__8277),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS1n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_3_0_LC_11_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_3_0_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_3_0_LC_11_9_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_3_0_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__8908),
            .in2(_gnd_net_),
            .in3(N__8873),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.CIA_STATE_d_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_11_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_11_9_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_11_9_1  (
            .in0(N__8787),
            .in1(N__8373),
            .in2(N__8271),
            .in3(N__8807),
            .lcout(\U409_TRANSFER_ACK.N_293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_9_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_9_2  (
            .in0(N__8806),
            .in1(N__8786),
            .in2(N__8384),
            .in3(N__8909),
            .lcout(\U409_TRANSFER_ACK.N_289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_9_3 .LUT_INIT=16'b0010001100100111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_9_3  (
            .in0(N__8178),
            .in1(N__8221),
            .in2(N__8206),
            .in3(N__8161),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_11_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_11_9_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_11_9_4 .LUT_INIT=16'b0000111110101010;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_LC_11_9_4  (
            .in0(N__8222),
            .in1(_gnd_net_),
            .in2(N__8262),
            .in3(N__9107),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_9_5 .LUT_INIT=16'b0100000001000100;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_9_5  (
            .in0(N__8180),
            .in1(N__9105),
            .in2(N__8208),
            .in3(N__8162),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_9_7 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_9_7  (
            .in0(N__8179),
            .in1(_gnd_net_),
            .in2(N__8207),
            .in3(N__9106),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_11_10_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_11_10_2 .LUT_INIT=16'b0111000001110001;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_LC_11_10_2  (
            .in0(N__8205),
            .in1(N__8181),
            .in2(N__8464),
            .in3(N__8163),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_ENC_net ),
            .ce(),
            .sr(N__9415));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_11_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_11_10_6 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_11_10_6  (
            .in0(N__8698),
            .in1(N__8148),
            .in2(N__8133),
            .in3(N__8106),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_ENC_net ),
            .ce(),
            .sr(N__9415));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_11_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_11_11_0 .LUT_INIT=16'b0011001100010010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_11_11_0  (
            .in0(N__8516),
            .in1(N__8626),
            .in2(N__8591),
            .in3(N__8546),
            .lcout(\U409_TRANSFER_ACK.N_307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_11_11_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_11_11_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__8581),
            .in2(_gnd_net_),
            .in3(N__8515),
            .lcout(\U409_TRANSFER_ACK.N_379 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_11_12_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_11_12_1 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_11_12_1  (
            .in0(N__8718),
            .in1(N__8712),
            .in2(N__8706),
            .in3(N__8518),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__9412));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_11_12_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_11_12_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(N__8547),
            .in2(_gnd_net_),
            .in3(N__8631),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__9412));
    defparam \U409_TRANSFER_ACK.ROMENn_LC_11_12_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_11_12_5 .SEQ_MODE=4'b1001;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_11_12_5 .LUT_INIT=16'b1011000011111010;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_LC_11_12_5  (
            .in0(N__8586),
            .in1(N__8676),
            .in2(N__8651),
            .in3(N__8670),
            .lcout(ROMENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__9412));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_11_12_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_11_12_7 .LUT_INIT=16'b0101101110100000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_11_12_7  (
            .in0(N__8630),
            .in1(N__8590),
            .in2(N__8553),
            .in3(N__8519),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__9412));
    defparam \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_11_14_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_11_14_7 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_11_14_7  (
            .in0(N__8465),
            .in1(N__8442),
            .in2(_gnd_net_),
            .in3(N__8421),
            .lcout(TCIn_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_4.C_ON=1'b0;
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_4.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8383),
            .lcout(GB_BUFFER_CLK40_IN_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNI692L_0_LC_12_5_1 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNI692L_0_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNI692L_0_LC_12_5_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_CIA.VMA_RNI692L_0_LC_12_5_1  (
            .in0(N__9696),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9044),
            .lcout(CIA_ENABLE),
            .ltout(CIA_ENABLE_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_12_5_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_12_5_2 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_12_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8772),
            .in3(N__8769),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS0n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_6_LC_12_7_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_6_LC_12_7_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_6_LC_12_7_0 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_6_LC_12_7_0  (
            .in0(N__9878),
            .in1(N__9801),
            .in2(N__8955),
            .in3(N__9849),
            .lcout(\U409_TICK.COUNTER60Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10654),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_12_7_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_12_7_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_TICK.COUNTER60_RNI2USG_10_LC_12_7_1  (
            .in0(N__9471),
            .in1(N__9504),
            .in2(N__9528),
            .in3(N__9452),
            .lcout(\U409_TICK.TICK603_10 ),
            .ltout(\U409_TICK.TICK603_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_15_LC_12_7_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_15_LC_12_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_15_LC_12_7_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_15_LC_12_7_2  (
            .in0(N__9877),
            .in1(N__9848),
            .in2(N__8733),
            .in3(N__9438),
            .lcout(\U409_TICK.COUNTER60Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10654),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_12_7_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_12_7_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER60_RNIDB4S_16_LC_12_7_3  (
            .in0(N__9486),
            .in1(N__8979),
            .in2(N__9000),
            .in3(N__9647),
            .lcout(\U409_TICK.TICK603_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_1_LC_12_7_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_1_LC_12_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_1_LC_12_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER60_1_LC_12_7_4  (
            .in0(_gnd_net_),
            .in1(N__8999),
            .in2(_gnd_net_),
            .in3(N__9978),
            .lcout(\U409_TICK.COUNTER60Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10654),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_1_LC_12_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_1_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_1_LC_12_9_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_1_1_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__8821),
            .in2(_gnd_net_),
            .in3(N__8844),
            .lcout(\U409_TRANSFER_ACK.N_223 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_4_0_LC_12_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_4_0_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_4_0_LC_12_9_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_4_0_LC_12_9_1  (
            .in0(N__8845),
            .in1(_gnd_net_),
            .in2(N__8828),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.m12_i_a2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_2_0_LC_12_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_2_0_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_2_0_LC_12_9_2 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_2_0_LC_12_9_2  (
            .in0(N__8875),
            .in1(N__8934),
            .in2(N__8730),
            .in3(N__8912),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.m12_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_12_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_12_9_3 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_0_LC_12_9_3  (
            .in0(N__9070),
            .in1(N__8853),
            .in2(N__8943),
            .in3(N__8940),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_12_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_12_9_4 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(N__8785),
            .in2(_gnd_net_),
            .in3(N__8805),
            .lcout(\U409_TRANSFER_ACK.N_191 ),
            .ltout(\U409_TRANSFER_ACK.N_191_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_9_5 .LUT_INIT=16'b0101000111011001;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_9_5  (
            .in0(N__8911),
            .in1(N__8876),
            .in2(N__8928),
            .in3(N__8925),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.i5_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_9_6 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8919),
            .in3(N__9071),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_12_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_12_9_7 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_12_9_7  (
            .in0(N__8846),
            .in1(N__8910),
            .in2(N__8829),
            .in3(N__8874),
            .lcout(\U409_TRANSFER_ACK.N_290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_10_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__9072),
            .in2(_gnd_net_),
            .in3(N__9689),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__9413));
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_12_10_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_12_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_0_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9548),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__9413));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_10_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8847),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__9413));
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_12_10_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_12_10_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_12_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_1_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8808),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__9413));
    defparam \U409_ADDRESS_DECODE.N_264_i_LC_12_11_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.N_264_i_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.N_264_i_LC_12_11_7 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \U409_ADDRESS_DECODE.N_264_i_LC_12_11_7  (
            .in0(N__9365),
            .in1(N__9339),
            .in2(N__9312),
            .in3(N__9248),
            .lcout(N_264_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_20_3.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_20_3.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_20_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9099),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_6_0 .C_ON=1'b1;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_6_0  (
            .in0(_gnd_net_),
            .in1(N__8990),
            .in2(N__9977),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_6_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_2_LC_13_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_2_LC_13_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_2_LC_13_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_2_LC_13_6_1  (
            .in0(_gnd_net_),
            .in1(N__8978),
            .in2(_gnd_net_),
            .in3(N__8967),
            .lcout(\U409_TICK.COUNTER60Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .clk(N__10648),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_3_LC_13_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_3_LC_13_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_3_LC_13_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_3_LC_13_6_2  (
            .in0(_gnd_net_),
            .in1(N__9617),
            .in2(_gnd_net_),
            .in3(N__8964),
            .lcout(\U409_TICK.COUNTER60Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .clk(N__10648),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_13_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_13_6_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_13_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_4_LC_13_6_3  (
            .in0(_gnd_net_),
            .in1(N__9944),
            .in2(_gnd_net_),
            .in3(N__8961),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_5_LC_13_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_5_LC_13_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_5_LC_13_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_5_LC_13_6_4  (
            .in0(_gnd_net_),
            .in1(N__9728),
            .in2(_gnd_net_),
            .in3(N__8958),
            .lcout(\U409_TICK.COUNTER60Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .clk(N__10648),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_13_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_13_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_13_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_6_LC_13_6_5  (
            .in0(_gnd_net_),
            .in1(N__9914),
            .in2(_gnd_net_),
            .in3(N__8946),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_7_LC_13_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_7_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_7_LC_13_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_7_LC_13_6_6  (
            .in0(_gnd_net_),
            .in1(N__9524),
            .in2(_gnd_net_),
            .in3(N__9513),
            .lcout(\U409_TICK.COUNTER60Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .clk(N__10648),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_13_6_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_13_6_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_13_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_8_LC_13_6_7  (
            .in0(_gnd_net_),
            .in1(N__9767),
            .in2(_gnd_net_),
            .in3(N__9510),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_13_7_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_13_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_9_LC_13_7_0  (
            .in0(_gnd_net_),
            .in1(N__9932),
            .in2(_gnd_net_),
            .in3(N__9507),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_13_7_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_10_LC_13_7_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_10_LC_13_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_10_LC_13_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_10_LC_13_7_1  (
            .in0(_gnd_net_),
            .in1(N__9503),
            .in2(_gnd_net_),
            .in3(N__9492),
            .lcout(\U409_TICK.COUNTER60Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .clk(N__10650),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_11_LC_13_7_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_11_LC_13_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_11_LC_13_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_11_LC_13_7_2  (
            .in0(_gnd_net_),
            .in1(N__9635),
            .in2(_gnd_net_),
            .in3(N__9489),
            .lcout(\U409_TICK.COUNTER60Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .clk(N__10650),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_12_LC_13_7_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_12_LC_13_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_12_LC_13_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_12_LC_13_7_3  (
            .in0(_gnd_net_),
            .in1(N__9485),
            .in2(_gnd_net_),
            .in3(N__9474),
            .lcout(\U409_TICK.COUNTER60Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .clk(N__10650),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_13_LC_13_7_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_13_LC_13_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_13_LC_13_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_13_LC_13_7_4  (
            .in0(_gnd_net_),
            .in1(N__9470),
            .in2(_gnd_net_),
            .in3(N__9459),
            .lcout(\U409_TICK.COUNTER60Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .clk(N__10650),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_13_7_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_13_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_14_LC_13_7_5  (
            .in0(_gnd_net_),
            .in1(N__9893),
            .in2(_gnd_net_),
            .in3(N__9456),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_13_7_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_13_7_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_15_LC_13_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9453),
            .in3(N__9432),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_16_LC_13_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_16_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_16_LC_13_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER60_16_LC_13_7_7  (
            .in0(_gnd_net_),
            .in1(N__9648),
            .in2(_gnd_net_),
            .in3(N__9651),
            .lcout(\U409_TICK.COUNTER60Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10650),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_13_8_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_13_8_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNI335G2_11_LC_13_8_6  (
            .in0(N__9717),
            .in1(N__9636),
            .in2(N__9624),
            .in3(N__9606),
            .lcout(\U409_TICK.TICK603_14 ),
            .ltout(\U409_TICK.TICK603_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK60_LC_13_8_7 .C_ON=1'b0;
    defparam \U409_TICK.TICK60_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK60_LC_13_8_7 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \U409_TICK.TICK60_LC_13_8_7  (
            .in0(N__9581),
            .in1(N__9802),
            .in2(N__9600),
            .in3(N__9847),
            .lcout(TICK60_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10653),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_13_10_0 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_13_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_13_10_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_0_LC_13_10_0  (
            .in0(N__10348),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10283),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_2_LC_13_10_1 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_2_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_2_LC_13_10_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_2_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(N__10344),
            .in2(_gnd_net_),
            .in3(N__10246),
            .lcout(),
            .ltout(\U409_CIA.CLK_CIA6_0_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_13_10_2 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_13_10_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_0_LC_13_10_2  (
            .in0(N__10319),
            .in1(N__10055),
            .in2(N__9570),
            .in3(N__10371),
            .lcout(),
            .ltout(\U409_CIA.CLK_CIA6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_LC_13_10_3 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_LC_13_10_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CLK_CIA_LC_13_10_3 .LUT_INIT=16'b0000111100001100;
    LogicCell40 \U409_CIA.CLK_CIA_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(N__9547),
            .in2(N__9567),
            .in3(N__10359),
            .lcout(CLK_CIA_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10283),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_2_LC_13_10_4 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_2_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_2_LC_13_10_4 .LUT_INIT=16'b0101000010100000;
    LogicCell40 \U409_CIA.VMA_RNO_2_LC_13_10_4  (
            .in0(N__10247),
            .in1(_gnd_net_),
            .in2(N__10353),
            .in3(N__10311),
            .lcout(),
            .ltout(\U409_CIA.un1_CIA_CLK_COUNT_3_0_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_1_LC_13_10_5 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_1_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_1_LC_13_10_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_CIA.VMA_RNO_1_LC_13_10_5  (
            .in0(N__10056),
            .in1(N__10269),
            .in2(N__9531),
            .in3(N__10224),
            .lcout(),
            .ltout(\U409_CIA.VMA_RNOZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_LC_13_10_6 .C_ON=1'b0;
    defparam \U409_CIA.VMA_LC_13_10_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.VMA_LC_13_10_6 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \U409_CIA.VMA_LC_13_10_6  (
            .in0(N__9711),
            .in1(N__9688),
            .in2(N__9699),
            .in3(N__10312),
            .lcout(\U409_CIA.VMAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10283),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_5_0 .C_ON=1'b1;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_5_0  (
            .in0(_gnd_net_),
            .in1(N__10123),
            .in2(N__10527),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_5_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_2_LC_14_5_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_2_LC_14_5_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_2_LC_14_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_2_LC_14_5_1  (
            .in0(_gnd_net_),
            .in1(N__10142),
            .in2(_gnd_net_),
            .in3(N__9672),
            .lcout(\U409_TICK.COUNTER50Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .clk(N__10649),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_3_LC_14_5_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_3_LC_14_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_3_LC_14_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_3_LC_14_5_2  (
            .in0(_gnd_net_),
            .in1(N__10538),
            .in2(_gnd_net_),
            .in3(N__9669),
            .lcout(\U409_TICK.COUNTER50Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .clk(N__10649),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_4_LC_14_5_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_4_LC_14_5_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_4_LC_14_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_4_LC_14_5_3  (
            .in0(_gnd_net_),
            .in1(N__10082),
            .in2(_gnd_net_),
            .in3(N__9666),
            .lcout(\U409_TICK.COUNTER50Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .clk(N__10649),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_14_5_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_14_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_5_LC_14_5_4  (
            .in0(_gnd_net_),
            .in1(N__10550),
            .in2(_gnd_net_),
            .in3(N__9663),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_14_5_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_14_5_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_14_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_6_LC_14_5_5  (
            .in0(_gnd_net_),
            .in1(N__10418),
            .in2(_gnd_net_),
            .in3(N__9660),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_7_LC_14_5_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_7_LC_14_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_7_LC_14_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_7_LC_14_5_6  (
            .in0(_gnd_net_),
            .in1(N__10097),
            .in2(_gnd_net_),
            .in3(N__9657),
            .lcout(\U409_TICK.COUNTER50Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .clk(N__10649),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_8_LC_14_5_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_8_LC_14_5_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_8_LC_14_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_8_LC_14_5_7  (
            .in0(_gnd_net_),
            .in1(N__10154),
            .in2(_gnd_net_),
            .in3(N__9654),
            .lcout(\U409_TICK.COUNTER50Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .clk(N__10649),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_14_6_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_14_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_9_LC_14_6_0  (
            .in0(_gnd_net_),
            .in1(N__10667),
            .in2(_gnd_net_),
            .in3(N__9753),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_14_6_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_10_LC_14_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_10_LC_14_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_10_LC_14_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_10_LC_14_6_1  (
            .in0(_gnd_net_),
            .in1(N__10475),
            .in2(_gnd_net_),
            .in3(N__9750),
            .lcout(\U409_TICK.COUNTER50Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .clk(N__10651),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_14_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_14_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_11_LC_14_6_2  (
            .in0(_gnd_net_),
            .in1(N__10385),
            .in2(_gnd_net_),
            .in3(N__9747),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_12_LC_14_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_12_LC_14_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_12_LC_14_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_12_LC_14_6_3  (
            .in0(_gnd_net_),
            .in1(N__10499),
            .in2(_gnd_net_),
            .in3(N__9744),
            .lcout(\U409_TICK.COUNTER50Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .clk(N__10651),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_14_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_14_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_13_LC_14_6_4  (
            .in0(_gnd_net_),
            .in1(N__10406),
            .in2(_gnd_net_),
            .in3(N__9741),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_14_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_14_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_14_LC_14_6_5  (
            .in0(_gnd_net_),
            .in1(N__10430),
            .in2(_gnd_net_),
            .in3(N__9738),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_14_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_14_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_15_LC_14_6_6  (
            .in0(_gnd_net_),
            .in1(N__10454),
            .in2(_gnd_net_),
            .in3(N__9735),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_16_LC_14_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_16_LC_14_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_16_LC_14_6_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER50_16_LC_14_6_7  (
            .in0(_gnd_net_),
            .in1(N__10110),
            .in2(_gnd_net_),
            .in3(N__9732),
            .lcout(\U409_TICK.COUNTER50Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10651),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_14_7_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_14_7_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_TICK.COUNTER60_RNIHJU51_4_LC_14_7_0  (
            .in0(N__9729),
            .in1(N__9945),
            .in2(_gnd_net_),
            .in3(N__9972),
            .lcout(\U409_TICK.TICK603_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_9_LC_14_7_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_9_LC_14_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_9_LC_14_7_1 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \U409_TICK.COUNTER60_9_LC_14_7_1  (
            .in0(N__9881),
            .in1(N__9984),
            .in2(N__9816),
            .in3(N__9846),
            .lcout(\U409_TICK.COUNTER60Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10655),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_0_LC_14_7_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_0_LC_14_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_0_LC_14_7_2 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \U409_TICK.COUNTER60_0_LC_14_7_2  (
            .in0(N__9843),
            .in1(N__9973),
            .in2(N__9882),
            .in3(N__9813),
            .lcout(\U409_TICK.COUNTER60Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10655),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_4_LC_14_7_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_4_LC_14_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_4_LC_14_7_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_4_LC_14_7_3  (
            .in0(N__9879),
            .in1(N__9844),
            .in2(N__9814),
            .in3(N__9951),
            .lcout(\U409_TICK.COUNTER60Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10655),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_14_7_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_14_7_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNICDC71_14_LC_14_7_4  (
            .in0(N__9933),
            .in1(N__9768),
            .in2(N__9921),
            .in3(N__9894),
            .lcout(\U409_TICK.TICK603_9 ),
            .ltout(\U409_TICK.TICK603_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_14_LC_14_7_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_14_LC_14_7_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_14_LC_14_7_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_14_LC_14_7_5  (
            .in0(N__9803),
            .in1(N__9873),
            .in2(N__9903),
            .in3(N__9900),
            .lcout(\U409_TICK.COUNTER60Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10655),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_8_LC_14_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_8_LC_14_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_8_LC_14_7_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_8_LC_14_7_7  (
            .in0(N__9880),
            .in1(N__9845),
            .in2(N__9815),
            .in3(N__9774),
            .lcout(\U409_TICK.COUNTER60Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10655),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_14_9_0 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_14_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_14_9_0  (
            .in0(_gnd_net_),
            .in1(N__10349),
            .in2(N__10320),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_9_0_),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_14_9_1 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_14_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_14_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_2_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(N__10223),
            .in2(_gnd_net_),
            .in3(N__9756),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .clk(N__10284),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_14_9_2 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_14_9_2 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_14_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_3_LC_14_9_2  (
            .in0(N__10043),
            .in1(N__9999),
            .in2(_gnd_net_),
            .in3(N__10071),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .clk(N__10284),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_14_9_3 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_14_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_14_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_4_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(N__10248),
            .in2(_gnd_net_),
            .in3(N__10068),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .clk(N__10284),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_14_9_4 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_14_9_4 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_14_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_5_LC_14_9_4  (
            .in0(N__10044),
            .in1(N__10268),
            .in2(_gnd_net_),
            .in3(N__10065),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .clk(N__10284),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_14_9_5 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_14_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_14_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_6_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(N__10032),
            .in2(_gnd_net_),
            .in3(N__10062),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ),
            .clk(N__10284),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_14_9_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_14_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_14_9_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_7_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(N__10016),
            .in2(_gnd_net_),
            .in3(N__10059),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10284),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIBFRM_2_LC_14_10_1 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIBFRM_2_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIBFRM_2_LC_14_10_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIBFRM_2_LC_14_10_1  (
            .in0(N__10267),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10222),
            .lcout(\U409_CIA.N_420 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIMC921_7_LC_14_10_2 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIMC921_7_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIMC921_7_LC_14_10_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIMC921_7_LC_14_10_2  (
            .in0(N__10012),
            .in1(N__10030),
            .in2(_gnd_net_),
            .in3(N__9997),
            .lcout(\U409_CIA.N_427 ),
            .ltout(\U409_CIA.N_427_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNICTDR2_0_LC_14_10_3 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNICTDR2_0_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNICTDR2_0_LC_14_10_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNICTDR2_0_LC_14_10_3  (
            .in0(N__10316),
            .in1(N__10350),
            .in2(N__10047),
            .in3(N__10203),
            .lcout(\U409_CIA.CIA_CLK_COUNT11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_3_LC_14_10_4 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_3_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_3_LC_14_10_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_3_LC_14_10_4  (
            .in0(N__10245),
            .in1(N__10031),
            .in2(N__10017),
            .in3(N__9998),
            .lcout(),
            .ltout(\U409_CIA.un1_CIA_CLK_COUNT_2_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_14_10_5 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_14_10_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_1_LC_14_10_5  (
            .in0(N__10317),
            .in1(N__10351),
            .in2(N__10374),
            .in3(N__10370),
            .lcout(\U409_CIA.CLK_CIA_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_14_10_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_14_10_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_14_10_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_1_LC_14_10_6  (
            .in0(N__10352),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10318),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10282),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_2_LC_14_10_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_2_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_2_LC_14_10_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIH7921_2_LC_14_10_7  (
            .in0(N__10266),
            .in1(N__10244),
            .in2(_gnd_net_),
            .in3(N__10221),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_0_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_5_LC_15_5_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_5_LC_15_5_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_5_LC_15_5_0 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_5_LC_15_5_0  (
            .in0(N__10746),
            .in1(N__10772),
            .in2(N__10197),
            .in3(N__10712),
            .lcout(\U409_TICK.COUNTER50Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10652),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK50_LC_15_5_1 .C_ON=1'b0;
    defparam \U409_TICK.TICK50_LC_15_5_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK50_LC_15_5_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK50_LC_15_5_1  (
            .in0(N__10774),
            .in1(N__10172),
            .in2(N__10716),
            .in3(N__10748),
            .lcout(TICK50_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10652),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_1_LC_15_5_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_1_LC_15_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_1_LC_15_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER50_1_LC_15_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10131),
            .in3(N__10525),
            .lcout(\U409_TICK.COUNTER50Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10652),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_6_LC_15_5_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_6_LC_15_5_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_6_LC_15_5_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_6_LC_15_5_3  (
            .in0(N__10773),
            .in1(N__10747),
            .in2(N__10715),
            .in3(N__10161),
            .lcout(\U409_TICK.COUNTER50Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10652),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_15_5_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_15_5_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_15_5_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER50_RNIUHF01_16_LC_15_5_4  (
            .in0(N__10155),
            .in1(N__10143),
            .in2(N__10130),
            .in3(N__10109),
            .lcout(\U409_TICK.TICK503_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_15_5_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_15_5_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_15_5_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNII24V_14_LC_15_5_6  (
            .in0(N__10431),
            .in1(N__10098),
            .in2(N__10086),
            .in3(N__10455),
            .lcout(\U409_TICK.TICK503_10 ),
            .ltout(\U409_TICK.TICK503_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_0_LC_15_5_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_0_LC_15_5_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_0_LC_15_5_7 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \U409_TICK.COUNTER50_0_LC_15_5_7  (
            .in0(N__10705),
            .in1(N__10745),
            .in2(N__10554),
            .in3(N__10526),
            .lcout(\U409_TICK.COUNTER50Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10652),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_15_6_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_15_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_15_6_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_TICK.COUNTER50_RNID6CP_3_LC_15_6_0  (
            .in0(N__10551),
            .in1(N__10539),
            .in2(_gnd_net_),
            .in3(N__10524),
            .lcout(),
            .ltout(\U409_TICK.TICK503_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_15_6_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_15_6_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_15_6_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_TICK.COUNTER50_RNITU182_10_LC_15_6_1  (
            .in0(N__10500),
            .in1(N__10488),
            .in2(N__10479),
            .in3(N__10476),
            .lcout(\U409_TICK.TICK503_14 ),
            .ltout(\U409_TICK.TICK503_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_15_LC_15_6_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_15_LC_15_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_15_LC_15_6_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_15_LC_15_6_2  (
            .in0(N__10778),
            .in1(N__10701),
            .in2(N__10464),
            .in3(N__10461),
            .lcout(\U409_TICK.COUNTER50Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10656),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_13_LC_15_6_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_13_LC_15_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_13_LC_15_6_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_13_LC_15_6_3  (
            .in0(N__10740),
            .in1(N__10776),
            .in2(N__10714),
            .in3(N__10443),
            .lcout(\U409_TICK.COUNTER50Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10656),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_14_LC_15_6_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_14_LC_15_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_14_LC_15_6_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_14_LC_15_6_4  (
            .in0(N__10777),
            .in1(N__10741),
            .in2(N__10713),
            .in3(N__10437),
            .lcout(\U409_TICK.COUNTER50Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10656),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_15_6_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_15_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_15_6_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNIH14V_11_LC_15_6_5  (
            .in0(N__10386),
            .in1(N__10419),
            .in2(N__10671),
            .in3(N__10407),
            .lcout(\U409_TICK.TICK503_9 ),
            .ltout(\U409_TICK.TICK503_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_11_LC_15_6_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_11_LC_15_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_11_LC_15_6_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_11_LC_15_6_6  (
            .in0(N__10775),
            .in1(N__10739),
            .in2(N__10395),
            .in3(N__10392),
            .lcout(\U409_TICK.COUNTER50Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10656),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_9_LC_15_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_9_LC_15_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_9_LC_15_6_7 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \U409_TICK.COUNTER50_9_LC_15_6_7  (
            .in0(N__10785),
            .in1(N__10779),
            .in2(N__10749),
            .in3(N__10700),
            .lcout(\U409_TICK.COUNTER50Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10656),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_19_8_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_19_8_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_19_8_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_19_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U409_TOP

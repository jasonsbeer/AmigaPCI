// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 14 2025 00:16:39

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U409_TOP" view "INTERFACE"

module U409_TOP (
    TM,
    TT,
    D,
    A,
    PIO_S0,
    PORTSIZE,
    TICK60,
    CIACS0n,
    CPUCONFn,
    CLK6,
    CLK_CIA,
    BUFENn,
    AUTOBOOT,
    RnW,
    PIO_P2,
    CIACS1n,
    BRIDGE_ENn,
    PIO_S1,
    PIO_P0,
    TICK50,
    TCIn,
    TBIn,
    RAMSPACEn,
    CLK40_IN,
    CLK28_IN,
    REGSPACEn,
    TSn,
    RTC_ENn,
    PIO_S2,
    ATA_ENn,
    RESETn,
    OVL,
    CONFIGENn,
    TACKn,
    ROMENn,
    PIO_P1);

    input [1:0] TM;
    input [1:0] TT;
    inout [7:4] D;
    input [31:1] A;
    output PIO_S0;
    output PORTSIZE;
    output TICK60;
    output CIACS0n;
    input CPUCONFn;
    input CLK6;
    output CLK_CIA;
    output BUFENn;
    input AUTOBOOT;
    input RnW;
    output PIO_P2;
    output CIACS1n;
    output BRIDGE_ENn;
    output PIO_S1;
    output PIO_P0;
    output TICK50;
    output TCIn;
    output TBIn;
    output RAMSPACEn;
    input CLK40_IN;
    input CLK28_IN;
    output REGSPACEn;
    input TSn;
    output RTC_ENn;
    output PIO_S2;
    output ATA_ENn;
    input RESETn;
    input OVL;
    output CONFIGENn;
    inout TACKn;
    output ROMENn;
    output PIO_P1;

    wire N__11324;
    wire N__11323;
    wire N__11322;
    wire N__11314;
    wire N__11313;
    wire N__11312;
    wire N__11304;
    wire N__11303;
    wire N__11302;
    wire N__11293;
    wire N__11292;
    wire N__11291;
    wire N__11284;
    wire N__11283;
    wire N__11282;
    wire N__11275;
    wire N__11274;
    wire N__11273;
    wire N__11266;
    wire N__11265;
    wire N__11264;
    wire N__11257;
    wire N__11256;
    wire N__11255;
    wire N__11248;
    wire N__11247;
    wire N__11246;
    wire N__11239;
    wire N__11238;
    wire N__11237;
    wire N__11230;
    wire N__11229;
    wire N__11228;
    wire N__11221;
    wire N__11220;
    wire N__11219;
    wire N__11212;
    wire N__11211;
    wire N__11210;
    wire N__11203;
    wire N__11202;
    wire N__11201;
    wire N__11194;
    wire N__11193;
    wire N__11192;
    wire N__11185;
    wire N__11184;
    wire N__11183;
    wire N__11176;
    wire N__11175;
    wire N__11174;
    wire N__11167;
    wire N__11166;
    wire N__11165;
    wire N__11158;
    wire N__11157;
    wire N__11156;
    wire N__11149;
    wire N__11148;
    wire N__11147;
    wire N__11140;
    wire N__11139;
    wire N__11138;
    wire N__11131;
    wire N__11130;
    wire N__11129;
    wire N__11122;
    wire N__11121;
    wire N__11120;
    wire N__11113;
    wire N__11112;
    wire N__11111;
    wire N__11104;
    wire N__11103;
    wire N__11102;
    wire N__11095;
    wire N__11094;
    wire N__11093;
    wire N__11086;
    wire N__11085;
    wire N__11084;
    wire N__11077;
    wire N__11076;
    wire N__11075;
    wire N__11068;
    wire N__11067;
    wire N__11066;
    wire N__11059;
    wire N__11058;
    wire N__11057;
    wire N__11050;
    wire N__11049;
    wire N__11048;
    wire N__11041;
    wire N__11040;
    wire N__11039;
    wire N__11032;
    wire N__11031;
    wire N__11030;
    wire N__11023;
    wire N__11022;
    wire N__11021;
    wire N__11014;
    wire N__11013;
    wire N__11012;
    wire N__11005;
    wire N__11004;
    wire N__11003;
    wire N__10996;
    wire N__10995;
    wire N__10994;
    wire N__10987;
    wire N__10986;
    wire N__10985;
    wire N__10978;
    wire N__10977;
    wire N__10976;
    wire N__10969;
    wire N__10968;
    wire N__10967;
    wire N__10960;
    wire N__10959;
    wire N__10958;
    wire N__10951;
    wire N__10950;
    wire N__10949;
    wire N__10942;
    wire N__10941;
    wire N__10940;
    wire N__10933;
    wire N__10932;
    wire N__10931;
    wire N__10924;
    wire N__10923;
    wire N__10922;
    wire N__10915;
    wire N__10914;
    wire N__10913;
    wire N__10906;
    wire N__10905;
    wire N__10904;
    wire N__10897;
    wire N__10896;
    wire N__10895;
    wire N__10888;
    wire N__10887;
    wire N__10886;
    wire N__10879;
    wire N__10878;
    wire N__10877;
    wire N__10870;
    wire N__10869;
    wire N__10868;
    wire N__10861;
    wire N__10860;
    wire N__10859;
    wire N__10852;
    wire N__10851;
    wire N__10850;
    wire N__10843;
    wire N__10842;
    wire N__10841;
    wire N__10834;
    wire N__10833;
    wire N__10832;
    wire N__10825;
    wire N__10824;
    wire N__10823;
    wire N__10816;
    wire N__10815;
    wire N__10814;
    wire N__10807;
    wire N__10806;
    wire N__10805;
    wire N__10798;
    wire N__10797;
    wire N__10796;
    wire N__10789;
    wire N__10788;
    wire N__10787;
    wire N__10780;
    wire N__10779;
    wire N__10778;
    wire N__10771;
    wire N__10770;
    wire N__10769;
    wire N__10762;
    wire N__10761;
    wire N__10760;
    wire N__10753;
    wire N__10752;
    wire N__10751;
    wire N__10744;
    wire N__10743;
    wire N__10742;
    wire N__10735;
    wire N__10734;
    wire N__10733;
    wire N__10716;
    wire N__10713;
    wire N__10710;
    wire N__10709;
    wire N__10706;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10691;
    wire N__10688;
    wire N__10685;
    wire N__10682;
    wire N__10679;
    wire N__10674;
    wire N__10671;
    wire N__10668;
    wire N__10665;
    wire N__10662;
    wire N__10659;
    wire N__10658;
    wire N__10653;
    wire N__10650;
    wire N__10647;
    wire N__10644;
    wire N__10641;
    wire N__10640;
    wire N__10637;
    wire N__10634;
    wire N__10631;
    wire N__10628;
    wire N__10623;
    wire N__10620;
    wire N__10617;
    wire N__10614;
    wire N__10611;
    wire N__10608;
    wire N__10605;
    wire N__10602;
    wire N__10599;
    wire N__10596;
    wire N__10593;
    wire N__10590;
    wire N__10587;
    wire N__10584;
    wire N__10583;
    wire N__10582;
    wire N__10581;
    wire N__10578;
    wire N__10575;
    wire N__10572;
    wire N__10569;
    wire N__10560;
    wire N__10557;
    wire N__10554;
    wire N__10551;
    wire N__10548;
    wire N__10547;
    wire N__10546;
    wire N__10545;
    wire N__10542;
    wire N__10539;
    wire N__10536;
    wire N__10533;
    wire N__10524;
    wire N__10521;
    wire N__10518;
    wire N__10517;
    wire N__10516;
    wire N__10515;
    wire N__10512;
    wire N__10509;
    wire N__10506;
    wire N__10503;
    wire N__10498;
    wire N__10491;
    wire N__10490;
    wire N__10489;
    wire N__10488;
    wire N__10479;
    wire N__10476;
    wire N__10473;
    wire N__10472;
    wire N__10471;
    wire N__10470;
    wire N__10469;
    wire N__10466;
    wire N__10461;
    wire N__10456;
    wire N__10449;
    wire N__10446;
    wire N__10445;
    wire N__10444;
    wire N__10443;
    wire N__10440;
    wire N__10437;
    wire N__10432;
    wire N__10425;
    wire N__10424;
    wire N__10423;
    wire N__10422;
    wire N__10419;
    wire N__10418;
    wire N__10415;
    wire N__10412;
    wire N__10407;
    wire N__10402;
    wire N__10395;
    wire N__10394;
    wire N__10393;
    wire N__10392;
    wire N__10391;
    wire N__10390;
    wire N__10387;
    wire N__10384;
    wire N__10377;
    wire N__10372;
    wire N__10365;
    wire N__10362;
    wire N__10359;
    wire N__10356;
    wire N__10355;
    wire N__10352;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10338;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10324;
    wire N__10321;
    wire N__10318;
    wire N__10315;
    wire N__10312;
    wire N__10309;
    wire N__10306;
    wire N__10299;
    wire N__10296;
    wire N__10295;
    wire N__10292;
    wire N__10289;
    wire N__10288;
    wire N__10283;
    wire N__10280;
    wire N__10279;
    wire N__10276;
    wire N__10273;
    wire N__10270;
    wire N__10269;
    wire N__10268;
    wire N__10265;
    wire N__10260;
    wire N__10255;
    wire N__10248;
    wire N__10245;
    wire N__10242;
    wire N__10239;
    wire N__10238;
    wire N__10235;
    wire N__10232;
    wire N__10231;
    wire N__10226;
    wire N__10223;
    wire N__10220;
    wire N__10217;
    wire N__10212;
    wire N__10209;
    wire N__10206;
    wire N__10203;
    wire N__10200;
    wire N__10197;
    wire N__10194;
    wire N__10191;
    wire N__10188;
    wire N__10187;
    wire N__10184;
    wire N__10181;
    wire N__10180;
    wire N__10179;
    wire N__10178;
    wire N__10177;
    wire N__10176;
    wire N__10171;
    wire N__10170;
    wire N__10169;
    wire N__10168;
    wire N__10167;
    wire N__10164;
    wire N__10161;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10153;
    wire N__10150;
    wire N__10149;
    wire N__10148;
    wire N__10147;
    wire N__10146;
    wire N__10145;
    wire N__10144;
    wire N__10141;
    wire N__10138;
    wire N__10135;
    wire N__10124;
    wire N__10121;
    wire N__10116;
    wire N__10113;
    wire N__10110;
    wire N__10107;
    wire N__10104;
    wire N__10101;
    wire N__10098;
    wire N__10095;
    wire N__10094;
    wire N__10081;
    wire N__10080;
    wire N__10073;
    wire N__10070;
    wire N__10063;
    wire N__10062;
    wire N__10061;
    wire N__10060;
    wire N__10057;
    wire N__10054;
    wire N__10051;
    wire N__10048;
    wire N__10043;
    wire N__10038;
    wire N__10035;
    wire N__10028;
    wire N__10027;
    wire N__10024;
    wire N__10017;
    wire N__10014;
    wire N__10011;
    wire N__10006;
    wire N__10005;
    wire N__10002;
    wire N__9999;
    wire N__9996;
    wire N__9993;
    wire N__9990;
    wire N__9983;
    wire N__9978;
    wire N__9975;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9965;
    wire N__9962;
    wire N__9961;
    wire N__9958;
    wire N__9955;
    wire N__9952;
    wire N__9945;
    wire N__9942;
    wire N__9939;
    wire N__9936;
    wire N__9933;
    wire N__9930;
    wire N__9927;
    wire N__9924;
    wire N__9921;
    wire N__9920;
    wire N__9919;
    wire N__9918;
    wire N__9917;
    wire N__9916;
    wire N__9911;
    wire N__9904;
    wire N__9901;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9885;
    wire N__9882;
    wire N__9879;
    wire N__9878;
    wire N__9875;
    wire N__9872;
    wire N__9867;
    wire N__9866;
    wire N__9863;
    wire N__9860;
    wire N__9855;
    wire N__9852;
    wire N__9851;
    wire N__9848;
    wire N__9845;
    wire N__9840;
    wire N__9837;
    wire N__9834;
    wire N__9833;
    wire N__9830;
    wire N__9827;
    wire N__9822;
    wire N__9819;
    wire N__9816;
    wire N__9815;
    wire N__9812;
    wire N__9809;
    wire N__9804;
    wire N__9801;
    wire N__9798;
    wire N__9797;
    wire N__9794;
    wire N__9791;
    wire N__9786;
    wire N__9785;
    wire N__9784;
    wire N__9783;
    wire N__9782;
    wire N__9781;
    wire N__9780;
    wire N__9779;
    wire N__9778;
    wire N__9773;
    wire N__9768;
    wire N__9759;
    wire N__9756;
    wire N__9753;
    wire N__9750;
    wire N__9741;
    wire N__9740;
    wire N__9737;
    wire N__9736;
    wire N__9735;
    wire N__9734;
    wire N__9733;
    wire N__9732;
    wire N__9731;
    wire N__9730;
    wire N__9727;
    wire N__9724;
    wire N__9719;
    wire N__9716;
    wire N__9707;
    wire N__9704;
    wire N__9699;
    wire N__9690;
    wire N__9687;
    wire N__9686;
    wire N__9685;
    wire N__9684;
    wire N__9683;
    wire N__9682;
    wire N__9681;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9669;
    wire N__9666;
    wire N__9663;
    wire N__9660;
    wire N__9657;
    wire N__9652;
    wire N__9649;
    wire N__9644;
    wire N__9639;
    wire N__9634;
    wire N__9627;
    wire N__9624;
    wire N__9621;
    wire N__9620;
    wire N__9617;
    wire N__9614;
    wire N__9609;
    wire N__9608;
    wire N__9607;
    wire N__9606;
    wire N__9605;
    wire N__9604;
    wire N__9603;
    wire N__9602;
    wire N__9601;
    wire N__9600;
    wire N__9599;
    wire N__9598;
    wire N__9573;
    wire N__9570;
    wire N__9567;
    wire N__9564;
    wire N__9561;
    wire N__9560;
    wire N__9557;
    wire N__9554;
    wire N__9549;
    wire N__9546;
    wire N__9543;
    wire N__9540;
    wire N__9537;
    wire N__9534;
    wire N__9533;
    wire N__9530;
    wire N__9527;
    wire N__9522;
    wire N__9519;
    wire N__9518;
    wire N__9515;
    wire N__9512;
    wire N__9507;
    wire N__9506;
    wire N__9503;
    wire N__9500;
    wire N__9497;
    wire N__9492;
    wire N__9489;
    wire N__9486;
    wire N__9483;
    wire N__9482;
    wire N__9479;
    wire N__9476;
    wire N__9471;
    wire N__9468;
    wire N__9465;
    wire N__9462;
    wire N__9459;
    wire N__9456;
    wire N__9453;
    wire N__9450;
    wire N__9447;
    wire N__9444;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9432;
    wire N__9429;
    wire N__9426;
    wire N__9423;
    wire N__9420;
    wire N__9417;
    wire N__9416;
    wire N__9413;
    wire N__9410;
    wire N__9407;
    wire N__9404;
    wire N__9399;
    wire N__9398;
    wire N__9397;
    wire N__9396;
    wire N__9395;
    wire N__9394;
    wire N__9393;
    wire N__9390;
    wire N__9383;
    wire N__9376;
    wire N__9369;
    wire N__9368;
    wire N__9367;
    wire N__9366;
    wire N__9365;
    wire N__9364;
    wire N__9363;
    wire N__9362;
    wire N__9359;
    wire N__9352;
    wire N__9343;
    wire N__9336;
    wire N__9335;
    wire N__9334;
    wire N__9333;
    wire N__9330;
    wire N__9329;
    wire N__9326;
    wire N__9325;
    wire N__9322;
    wire N__9319;
    wire N__9318;
    wire N__9315;
    wire N__9310;
    wire N__9301;
    wire N__9298;
    wire N__9291;
    wire N__9288;
    wire N__9285;
    wire N__9282;
    wire N__9279;
    wire N__9276;
    wire N__9275;
    wire N__9272;
    wire N__9269;
    wire N__9264;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9246;
    wire N__9243;
    wire N__9240;
    wire N__9237;
    wire N__9234;
    wire N__9231;
    wire N__9228;
    wire N__9227;
    wire N__9224;
    wire N__9221;
    wire N__9216;
    wire N__9213;
    wire N__9210;
    wire N__9207;
    wire N__9204;
    wire N__9201;
    wire N__9200;
    wire N__9199;
    wire N__9196;
    wire N__9193;
    wire N__9192;
    wire N__9189;
    wire N__9186;
    wire N__9183;
    wire N__9180;
    wire N__9177;
    wire N__9168;
    wire N__9165;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9147;
    wire N__9144;
    wire N__9141;
    wire N__9140;
    wire N__9137;
    wire N__9134;
    wire N__9129;
    wire N__9128;
    wire N__9125;
    wire N__9124;
    wire N__9121;
    wire N__9120;
    wire N__9117;
    wire N__9114;
    wire N__9111;
    wire N__9108;
    wire N__9105;
    wire N__9102;
    wire N__9093;
    wire N__9090;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9078;
    wire N__9075;
    wire N__9072;
    wire N__9069;
    wire N__9066;
    wire N__9063;
    wire N__9060;
    wire N__9057;
    wire N__9054;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9042;
    wire N__9039;
    wire N__9036;
    wire N__9033;
    wire N__9030;
    wire N__9029;
    wire N__9028;
    wire N__9027;
    wire N__9026;
    wire N__9025;
    wire N__9024;
    wire N__9023;
    wire N__9020;
    wire N__9019;
    wire N__9018;
    wire N__9017;
    wire N__9016;
    wire N__8991;
    wire N__8988;
    wire N__8985;
    wire N__8982;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8970;
    wire N__8967;
    wire N__8966;
    wire N__8965;
    wire N__8964;
    wire N__8959;
    wire N__8954;
    wire N__8949;
    wire N__8948;
    wire N__8947;
    wire N__8946;
    wire N__8945;
    wire N__8938;
    wire N__8933;
    wire N__8928;
    wire N__8927;
    wire N__8926;
    wire N__8925;
    wire N__8924;
    wire N__8919;
    wire N__8914;
    wire N__8911;
    wire N__8904;
    wire N__8903;
    wire N__8900;
    wire N__8899;
    wire N__8898;
    wire N__8895;
    wire N__8894;
    wire N__8893;
    wire N__8892;
    wire N__8885;
    wire N__8880;
    wire N__8875;
    wire N__8868;
    wire N__8867;
    wire N__8866;
    wire N__8865;
    wire N__8862;
    wire N__8857;
    wire N__8854;
    wire N__8847;
    wire N__8846;
    wire N__8843;
    wire N__8838;
    wire N__8835;
    wire N__8834;
    wire N__8833;
    wire N__8832;
    wire N__8831;
    wire N__8826;
    wire N__8823;
    wire N__8818;
    wire N__8815;
    wire N__8808;
    wire N__8805;
    wire N__8804;
    wire N__8803;
    wire N__8802;
    wire N__8799;
    wire N__8798;
    wire N__8797;
    wire N__8788;
    wire N__8783;
    wire N__8778;
    wire N__8777;
    wire N__8774;
    wire N__8773;
    wire N__8770;
    wire N__8767;
    wire N__8766;
    wire N__8763;
    wire N__8760;
    wire N__8757;
    wire N__8754;
    wire N__8751;
    wire N__8748;
    wire N__8743;
    wire N__8740;
    wire N__8735;
    wire N__8730;
    wire N__8729;
    wire N__8728;
    wire N__8725;
    wire N__8722;
    wire N__8719;
    wire N__8712;
    wire N__8709;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8697;
    wire N__8696;
    wire N__8693;
    wire N__8690;
    wire N__8685;
    wire N__8682;
    wire N__8681;
    wire N__8678;
    wire N__8675;
    wire N__8670;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8658;
    wire N__8655;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8643;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8628;
    wire N__8625;
    wire N__8622;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8610;
    wire N__8607;
    wire N__8604;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8592;
    wire N__8589;
    wire N__8586;
    wire N__8585;
    wire N__8584;
    wire N__8583;
    wire N__8580;
    wire N__8577;
    wire N__8572;
    wire N__8569;
    wire N__8562;
    wire N__8559;
    wire N__8558;
    wire N__8553;
    wire N__8550;
    wire N__8549;
    wire N__8548;
    wire N__8541;
    wire N__8538;
    wire N__8537;
    wire N__8536;
    wire N__8535;
    wire N__8532;
    wire N__8525;
    wire N__8520;
    wire N__8519;
    wire N__8518;
    wire N__8515;
    wire N__8510;
    wire N__8505;
    wire N__8502;
    wire N__8499;
    wire N__8496;
    wire N__8493;
    wire N__8490;
    wire N__8487;
    wire N__8484;
    wire N__8481;
    wire N__8478;
    wire N__8475;
    wire N__8472;
    wire N__8469;
    wire N__8466;
    wire N__8463;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8451;
    wire N__8448;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8436;
    wire N__8435;
    wire N__8432;
    wire N__8429;
    wire N__8426;
    wire N__8421;
    wire N__8420;
    wire N__8419;
    wire N__8416;
    wire N__8413;
    wire N__8410;
    wire N__8403;
    wire N__8400;
    wire N__8397;
    wire N__8394;
    wire N__8391;
    wire N__8388;
    wire N__8385;
    wire N__8382;
    wire N__8379;
    wire N__8376;
    wire N__8373;
    wire N__8370;
    wire N__8369;
    wire N__8368;
    wire N__8367;
    wire N__8364;
    wire N__8361;
    wire N__8358;
    wire N__8355;
    wire N__8350;
    wire N__8349;
    wire N__8348;
    wire N__8345;
    wire N__8340;
    wire N__8337;
    wire N__8334;
    wire N__8331;
    wire N__8326;
    wire N__8321;
    wire N__8318;
    wire N__8313;
    wire N__8310;
    wire N__8307;
    wire N__8306;
    wire N__8305;
    wire N__8304;
    wire N__8303;
    wire N__8302;
    wire N__8301;
    wire N__8298;
    wire N__8295;
    wire N__8292;
    wire N__8289;
    wire N__8286;
    wire N__8283;
    wire N__8280;
    wire N__8277;
    wire N__8274;
    wire N__8271;
    wire N__8270;
    wire N__8269;
    wire N__8268;
    wire N__8267;
    wire N__8266;
    wire N__8265;
    wire N__8264;
    wire N__8263;
    wire N__8262;
    wire N__8259;
    wire N__8256;
    wire N__8253;
    wire N__8250;
    wire N__8247;
    wire N__8244;
    wire N__8211;
    wire N__8208;
    wire N__8205;
    wire N__8204;
    wire N__8201;
    wire N__8198;
    wire N__8193;
    wire N__8192;
    wire N__8191;
    wire N__8190;
    wire N__8187;
    wire N__8184;
    wire N__8181;
    wire N__8174;
    wire N__8169;
    wire N__8166;
    wire N__8163;
    wire N__8160;
    wire N__8157;
    wire N__8154;
    wire N__8153;
    wire N__8150;
    wire N__8147;
    wire N__8142;
    wire N__8139;
    wire N__8136;
    wire N__8135;
    wire N__8130;
    wire N__8127;
    wire N__8124;
    wire N__8121;
    wire N__8118;
    wire N__8117;
    wire N__8114;
    wire N__8111;
    wire N__8106;
    wire N__8103;
    wire N__8102;
    wire N__8101;
    wire N__8094;
    wire N__8091;
    wire N__8088;
    wire N__8085;
    wire N__8082;
    wire N__8079;
    wire N__8076;
    wire N__8075;
    wire N__8070;
    wire N__8067;
    wire N__8066;
    wire N__8065;
    wire N__8064;
    wire N__8061;
    wire N__8058;
    wire N__8057;
    wire N__8054;
    wire N__8045;
    wire N__8040;
    wire N__8037;
    wire N__8034;
    wire N__8033;
    wire N__8032;
    wire N__8029;
    wire N__8024;
    wire N__8021;
    wire N__8016;
    wire N__8015;
    wire N__8012;
    wire N__8009;
    wire N__8004;
    wire N__8003;
    wire N__8002;
    wire N__8001;
    wire N__7998;
    wire N__7991;
    wire N__7986;
    wire N__7983;
    wire N__7982;
    wire N__7979;
    wire N__7976;
    wire N__7975;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7950;
    wire N__7947;
    wire N__7946;
    wire N__7945;
    wire N__7942;
    wire N__7937;
    wire N__7932;
    wire N__7929;
    wire N__7926;
    wire N__7925;
    wire N__7922;
    wire N__7921;
    wire N__7918;
    wire N__7915;
    wire N__7914;
    wire N__7913;
    wire N__7910;
    wire N__7909;
    wire N__7904;
    wire N__7901;
    wire N__7894;
    wire N__7887;
    wire N__7884;
    wire N__7881;
    wire N__7878;
    wire N__7877;
    wire N__7876;
    wire N__7873;
    wire N__7870;
    wire N__7869;
    wire N__7866;
    wire N__7865;
    wire N__7862;
    wire N__7859;
    wire N__7856;
    wire N__7851;
    wire N__7842;
    wire N__7841;
    wire N__7838;
    wire N__7835;
    wire N__7830;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7818;
    wire N__7817;
    wire N__7814;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7800;
    wire N__7797;
    wire N__7794;
    wire N__7793;
    wire N__7790;
    wire N__7787;
    wire N__7782;
    wire N__7779;
    wire N__7776;
    wire N__7773;
    wire N__7770;
    wire N__7767;
    wire N__7764;
    wire N__7761;
    wire N__7760;
    wire N__7757;
    wire N__7754;
    wire N__7753;
    wire N__7750;
    wire N__7747;
    wire N__7744;
    wire N__7737;
    wire N__7736;
    wire N__7733;
    wire N__7730;
    wire N__7725;
    wire N__7724;
    wire N__7721;
    wire N__7718;
    wire N__7713;
    wire N__7712;
    wire N__7707;
    wire N__7704;
    wire N__7701;
    wire N__7698;
    wire N__7695;
    wire N__7692;
    wire N__7689;
    wire N__7686;
    wire N__7683;
    wire N__7680;
    wire N__7677;
    wire N__7674;
    wire N__7671;
    wire N__7668;
    wire N__7665;
    wire N__7664;
    wire N__7661;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7637;
    wire N__7634;
    wire N__7631;
    wire N__7626;
    wire N__7625;
    wire N__7624;
    wire N__7623;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7609;
    wire N__7602;
    wire N__7601;
    wire N__7600;
    wire N__7599;
    wire N__7598;
    wire N__7593;
    wire N__7590;
    wire N__7585;
    wire N__7578;
    wire N__7575;
    wire N__7572;
    wire N__7569;
    wire N__7566;
    wire N__7563;
    wire N__7560;
    wire N__7557;
    wire N__7554;
    wire N__7551;
    wire N__7548;
    wire N__7545;
    wire N__7544;
    wire N__7541;
    wire N__7538;
    wire N__7535;
    wire N__7530;
    wire N__7527;
    wire N__7526;
    wire N__7523;
    wire N__7520;
    wire N__7515;
    wire N__7514;
    wire N__7513;
    wire N__7512;
    wire N__7509;
    wire N__7502;
    wire N__7497;
    wire N__7494;
    wire N__7491;
    wire N__7488;
    wire N__7485;
    wire N__7484;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7472;
    wire N__7467;
    wire N__7464;
    wire N__7461;
    wire N__7460;
    wire N__7457;
    wire N__7454;
    wire N__7449;
    wire N__7446;
    wire N__7443;
    wire N__7440;
    wire N__7439;
    wire N__7436;
    wire N__7433;
    wire N__7432;
    wire N__7429;
    wire N__7426;
    wire N__7423;
    wire N__7420;
    wire N__7417;
    wire N__7414;
    wire N__7411;
    wire N__7406;
    wire N__7401;
    wire N__7398;
    wire N__7397;
    wire N__7394;
    wire N__7391;
    wire N__7386;
    wire N__7385;
    wire N__7384;
    wire N__7383;
    wire N__7380;
    wire N__7373;
    wire N__7368;
    wire N__7367;
    wire N__7364;
    wire N__7361;
    wire N__7356;
    wire N__7355;
    wire N__7354;
    wire N__7353;
    wire N__7352;
    wire N__7351;
    wire N__7348;
    wire N__7347;
    wire N__7346;
    wire N__7339;
    wire N__7338;
    wire N__7327;
    wire N__7326;
    wire N__7325;
    wire N__7322;
    wire N__7319;
    wire N__7316;
    wire N__7311;
    wire N__7308;
    wire N__7305;
    wire N__7300;
    wire N__7293;
    wire N__7292;
    wire N__7291;
    wire N__7288;
    wire N__7283;
    wire N__7278;
    wire N__7277;
    wire N__7274;
    wire N__7271;
    wire N__7268;
    wire N__7265;
    wire N__7264;
    wire N__7259;
    wire N__7256;
    wire N__7253;
    wire N__7250;
    wire N__7247;
    wire N__7244;
    wire N__7239;
    wire N__7236;
    wire N__7233;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7221;
    wire N__7220;
    wire N__7217;
    wire N__7214;
    wire N__7211;
    wire N__7208;
    wire N__7203;
    wire N__7202;
    wire N__7197;
    wire N__7196;
    wire N__7193;
    wire N__7190;
    wire N__7189;
    wire N__7186;
    wire N__7183;
    wire N__7180;
    wire N__7173;
    wire N__7170;
    wire N__7169;
    wire N__7168;
    wire N__7167;
    wire N__7166;
    wire N__7163;
    wire N__7162;
    wire N__7161;
    wire N__7160;
    wire N__7159;
    wire N__7154;
    wire N__7151;
    wire N__7150;
    wire N__7147;
    wire N__7146;
    wire N__7143;
    wire N__7140;
    wire N__7137;
    wire N__7134;
    wire N__7131;
    wire N__7126;
    wire N__7123;
    wire N__7120;
    wire N__7117;
    wire N__7114;
    wire N__7105;
    wire N__7102;
    wire N__7095;
    wire N__7090;
    wire N__7085;
    wire N__7080;
    wire N__7077;
    wire N__7074;
    wire N__7073;
    wire N__7070;
    wire N__7067;
    wire N__7066;
    wire N__7061;
    wire N__7058;
    wire N__7055;
    wire N__7052;
    wire N__7049;
    wire N__7046;
    wire N__7043;
    wire N__7040;
    wire N__7037;
    wire N__7032;
    wire N__7031;
    wire N__7028;
    wire N__7027;
    wire N__7024;
    wire N__7021;
    wire N__7018;
    wire N__7015;
    wire N__7012;
    wire N__7009;
    wire N__7006;
    wire N__7001;
    wire N__6998;
    wire N__6995;
    wire N__6990;
    wire N__6987;
    wire N__6986;
    wire N__6983;
    wire N__6980;
    wire N__6977;
    wire N__6974;
    wire N__6969;
    wire N__6966;
    wire N__6963;
    wire N__6960;
    wire N__6957;
    wire N__6954;
    wire N__6951;
    wire N__6948;
    wire N__6945;
    wire N__6942;
    wire N__6939;
    wire N__6936;
    wire N__6933;
    wire N__6932;
    wire N__6929;
    wire N__6926;
    wire N__6925;
    wire N__6924;
    wire N__6923;
    wire N__6920;
    wire N__6917;
    wire N__6914;
    wire N__6911;
    wire N__6908;
    wire N__6907;
    wire N__6906;
    wire N__6903;
    wire N__6900;
    wire N__6897;
    wire N__6894;
    wire N__6893;
    wire N__6890;
    wire N__6887;
    wire N__6884;
    wire N__6875;
    wire N__6872;
    wire N__6869;
    wire N__6866;
    wire N__6859;
    wire N__6854;
    wire N__6851;
    wire N__6846;
    wire N__6843;
    wire N__6840;
    wire N__6837;
    wire N__6834;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6822;
    wire N__6819;
    wire N__6816;
    wire N__6813;
    wire N__6810;
    wire N__6807;
    wire N__6806;
    wire N__6805;
    wire N__6802;
    wire N__6799;
    wire N__6796;
    wire N__6789;
    wire N__6786;
    wire N__6783;
    wire N__6780;
    wire N__6777;
    wire N__6774;
    wire N__6771;
    wire N__6768;
    wire N__6767;
    wire N__6762;
    wire N__6759;
    wire N__6758;
    wire N__6755;
    wire N__6752;
    wire N__6747;
    wire N__6746;
    wire N__6741;
    wire N__6738;
    wire N__6735;
    wire N__6732;
    wire N__6731;
    wire N__6728;
    wire N__6725;
    wire N__6720;
    wire N__6717;
    wire N__6716;
    wire N__6711;
    wire N__6708;
    wire N__6705;
    wire N__6702;
    wire N__6699;
    wire N__6698;
    wire N__6697;
    wire N__6694;
    wire N__6691;
    wire N__6688;
    wire N__6685;
    wire N__6680;
    wire N__6677;
    wire N__6674;
    wire N__6669;
    wire N__6666;
    wire N__6663;
    wire N__6660;
    wire N__6659;
    wire N__6656;
    wire N__6653;
    wire N__6648;
    wire N__6645;
    wire N__6644;
    wire N__6641;
    wire N__6638;
    wire N__6635;
    wire N__6632;
    wire N__6627;
    wire N__6624;
    wire N__6621;
    wire N__6620;
    wire N__6617;
    wire N__6614;
    wire N__6609;
    wire N__6608;
    wire N__6607;
    wire N__6606;
    wire N__6603;
    wire N__6596;
    wire N__6591;
    wire N__6590;
    wire N__6589;
    wire N__6588;
    wire N__6585;
    wire N__6584;
    wire N__6581;
    wire N__6580;
    wire N__6577;
    wire N__6576;
    wire N__6575;
    wire N__6574;
    wire N__6573;
    wire N__6570;
    wire N__6567;
    wire N__6564;
    wire N__6561;
    wire N__6558;
    wire N__6553;
    wire N__6550;
    wire N__6547;
    wire N__6544;
    wire N__6541;
    wire N__6528;
    wire N__6523;
    wire N__6520;
    wire N__6517;
    wire N__6514;
    wire N__6507;
    wire N__6504;
    wire N__6503;
    wire N__6500;
    wire N__6497;
    wire N__6492;
    wire N__6491;
    wire N__6488;
    wire N__6487;
    wire N__6486;
    wire N__6485;
    wire N__6482;
    wire N__6481;
    wire N__6480;
    wire N__6479;
    wire N__6478;
    wire N__6475;
    wire N__6472;
    wire N__6469;
    wire N__6466;
    wire N__6463;
    wire N__6460;
    wire N__6457;
    wire N__6454;
    wire N__6451;
    wire N__6442;
    wire N__6439;
    wire N__6432;
    wire N__6429;
    wire N__6426;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6412;
    wire N__6409;
    wire N__6406;
    wire N__6403;
    wire N__6400;
    wire N__6395;
    wire N__6390;
    wire N__6387;
    wire N__6384;
    wire N__6383;
    wire N__6382;
    wire N__6381;
    wire N__6380;
    wire N__6379;
    wire N__6376;
    wire N__6373;
    wire N__6372;
    wire N__6371;
    wire N__6368;
    wire N__6363;
    wire N__6362;
    wire N__6361;
    wire N__6360;
    wire N__6359;
    wire N__6358;
    wire N__6357;
    wire N__6354;
    wire N__6353;
    wire N__6352;
    wire N__6351;
    wire N__6346;
    wire N__6343;
    wire N__6342;
    wire N__6341;
    wire N__6336;
    wire N__6333;
    wire N__6326;
    wire N__6321;
    wire N__6314;
    wire N__6311;
    wire N__6308;
    wire N__6303;
    wire N__6300;
    wire N__6297;
    wire N__6294;
    wire N__6291;
    wire N__6286;
    wire N__6279;
    wire N__6272;
    wire N__6269;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6253;
    wire N__6250;
    wire N__6245;
    wire N__6242;
    wire N__6239;
    wire N__6236;
    wire N__6231;
    wire N__6230;
    wire N__6227;
    wire N__6226;
    wire N__6223;
    wire N__6220;
    wire N__6217;
    wire N__6216;
    wire N__6215;
    wire N__6214;
    wire N__6213;
    wire N__6212;
    wire N__6211;
    wire N__6210;
    wire N__6207;
    wire N__6204;
    wire N__6201;
    wire N__6196;
    wire N__6191;
    wire N__6184;
    wire N__6171;
    wire N__6168;
    wire N__6167;
    wire N__6166;
    wire N__6165;
    wire N__6164;
    wire N__6163;
    wire N__6160;
    wire N__6155;
    wire N__6150;
    wire N__6147;
    wire N__6140;
    wire N__6135;
    wire N__6134;
    wire N__6133;
    wire N__6132;
    wire N__6131;
    wire N__6128;
    wire N__6125;
    wire N__6122;
    wire N__6119;
    wire N__6116;
    wire N__6115;
    wire N__6114;
    wire N__6111;
    wire N__6106;
    wire N__6101;
    wire N__6098;
    wire N__6095;
    wire N__6090;
    wire N__6083;
    wire N__6080;
    wire N__6077;
    wire N__6072;
    wire N__6069;
    wire N__6066;
    wire N__6063;
    wire N__6062;
    wire N__6059;
    wire N__6056;
    wire N__6051;
    wire N__6048;
    wire N__6047;
    wire N__6046;
    wire N__6045;
    wire N__6042;
    wire N__6039;
    wire N__6036;
    wire N__6033;
    wire N__6032;
    wire N__6029;
    wire N__6022;
    wire N__6019;
    wire N__6016;
    wire N__6013;
    wire N__6010;
    wire N__6003;
    wire N__6000;
    wire N__5997;
    wire N__5994;
    wire N__5991;
    wire N__5988;
    wire N__5985;
    wire N__5982;
    wire N__5981;
    wire N__5980;
    wire N__5977;
    wire N__5974;
    wire N__5971;
    wire N__5968;
    wire N__5965;
    wire N__5962;
    wire N__5959;
    wire N__5956;
    wire N__5953;
    wire N__5950;
    wire N__5947;
    wire N__5944;
    wire N__5937;
    wire N__5934;
    wire N__5931;
    wire N__5928;
    wire N__5925;
    wire N__5922;
    wire N__5919;
    wire N__5916;
    wire N__5913;
    wire N__5910;
    wire N__5907;
    wire N__5904;
    wire N__5903;
    wire N__5902;
    wire N__5899;
    wire N__5896;
    wire N__5893;
    wire N__5890;
    wire N__5887;
    wire N__5884;
    wire N__5879;
    wire N__5876;
    wire N__5873;
    wire N__5870;
    wire N__5867;
    wire N__5862;
    wire N__5859;
    wire N__5856;
    wire N__5853;
    wire N__5852;
    wire N__5849;
    wire N__5846;
    wire N__5845;
    wire N__5840;
    wire N__5837;
    wire N__5834;
    wire N__5831;
    wire N__5828;
    wire N__5823;
    wire N__5820;
    wire N__5817;
    wire N__5814;
    wire N__5811;
    wire N__5808;
    wire N__5805;
    wire N__5804;
    wire N__5801;
    wire N__5798;
    wire N__5793;
    wire N__5792;
    wire N__5791;
    wire N__5790;
    wire N__5789;
    wire N__5786;
    wire N__5777;
    wire N__5772;
    wire N__5771;
    wire N__5770;
    wire N__5769;
    wire N__5768;
    wire N__5765;
    wire N__5756;
    wire N__5751;
    wire N__5750;
    wire N__5749;
    wire N__5746;
    wire N__5741;
    wire N__5738;
    wire N__5735;
    wire N__5734;
    wire N__5729;
    wire N__5726;
    wire N__5721;
    wire N__5718;
    wire N__5715;
    wire N__5712;
    wire N__5711;
    wire N__5710;
    wire N__5707;
    wire N__5706;
    wire N__5705;
    wire N__5704;
    wire N__5703;
    wire N__5700;
    wire N__5697;
    wire N__5694;
    wire N__5689;
    wire N__5686;
    wire N__5683;
    wire N__5680;
    wire N__5667;
    wire N__5666;
    wire N__5665;
    wire N__5660;
    wire N__5657;
    wire N__5656;
    wire N__5653;
    wire N__5650;
    wire N__5647;
    wire N__5642;
    wire N__5639;
    wire N__5636;
    wire N__5631;
    wire N__5628;
    wire N__5625;
    wire N__5624;
    wire N__5621;
    wire N__5618;
    wire N__5617;
    wire N__5614;
    wire N__5611;
    wire N__5610;
    wire N__5607;
    wire N__5604;
    wire N__5601;
    wire N__5598;
    wire N__5595;
    wire N__5588;
    wire N__5585;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5571;
    wire N__5568;
    wire N__5567;
    wire N__5564;
    wire N__5561;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5549;
    wire N__5546;
    wire N__5545;
    wire N__5544;
    wire N__5543;
    wire N__5540;
    wire N__5539;
    wire N__5536;
    wire N__5531;
    wire N__5526;
    wire N__5523;
    wire N__5520;
    wire N__5517;
    wire N__5512;
    wire N__5507;
    wire N__5504;
    wire N__5499;
    wire N__5496;
    wire N__5493;
    wire N__5490;
    wire N__5487;
    wire N__5484;
    wire N__5481;
    wire N__5480;
    wire N__5479;
    wire N__5478;
    wire N__5473;
    wire N__5472;
    wire N__5471;
    wire N__5470;
    wire N__5467;
    wire N__5464;
    wire N__5461;
    wire N__5456;
    wire N__5451;
    wire N__5448;
    wire N__5445;
    wire N__5438;
    wire N__5435;
    wire N__5432;
    wire N__5427;
    wire N__5424;
    wire N__5421;
    wire N__5418;
    wire N__5415;
    wire N__5412;
    wire N__5409;
    wire N__5406;
    wire N__5403;
    wire N__5400;
    wire N__5397;
    wire N__5394;
    wire N__5391;
    wire N__5388;
    wire N__5385;
    wire N__5382;
    wire N__5379;
    wire N__5376;
    wire N__5375;
    wire N__5370;
    wire N__5367;
    wire N__5364;
    wire N__5363;
    wire N__5358;
    wire N__5355;
    wire N__5352;
    wire N__5349;
    wire N__5346;
    wire N__5345;
    wire N__5342;
    wire N__5339;
    wire N__5334;
    wire N__5333;
    wire N__5330;
    wire N__5327;
    wire N__5324;
    wire N__5321;
    wire N__5316;
    wire N__5313;
    wire N__5310;
    wire N__5307;
    wire N__5304;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5292;
    wire N__5289;
    wire N__5286;
    wire N__5285;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5268;
    wire N__5265;
    wire N__5262;
    wire N__5259;
    wire N__5256;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5235;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5223;
    wire N__5220;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5208;
    wire N__5205;
    wire N__5202;
    wire N__5199;
    wire N__5196;
    wire N__5193;
    wire N__5192;
    wire N__5189;
    wire N__5188;
    wire N__5185;
    wire N__5184;
    wire N__5175;
    wire N__5172;
    wire N__5169;
    wire N__5166;
    wire N__5163;
    wire N__5160;
    wire N__5157;
    wire N__5156;
    wire N__5155;
    wire N__5152;
    wire N__5149;
    wire N__5146;
    wire N__5139;
    wire N__5136;
    wire N__5135;
    wire N__5132;
    wire N__5129;
    wire N__5124;
    wire N__5121;
    wire N__5118;
    wire N__5115;
    wire N__5112;
    wire N__5109;
    wire N__5106;
    wire N__5103;
    wire N__5100;
    wire N__5097;
    wire N__5094;
    wire N__5091;
    wire N__5088;
    wire N__5085;
    wire N__5082;
    wire N__5079;
    wire N__5076;
    wire N__5073;
    wire N__5070;
    wire N__5067;
    wire N__5064;
    wire N__5061;
    wire N__5058;
    wire N__5055;
    wire N__5052;
    wire N__5049;
    wire N__5046;
    wire N__5043;
    wire N__5040;
    wire N__5037;
    wire N__5034;
    wire N__5031;
    wire N__5028;
    wire N__5025;
    wire N__5022;
    wire N__5019;
    wire N__5018;
    wire N__5017;
    wire N__5016;
    wire N__5011;
    wire N__5006;
    wire N__5001;
    wire N__5000;
    wire N__4997;
    wire N__4994;
    wire N__4991;
    wire N__4988;
    wire N__4985;
    wire N__4980;
    wire N__4977;
    wire N__4976;
    wire N__4975;
    wire N__4974;
    wire N__4971;
    wire N__4968;
    wire N__4965;
    wire N__4964;
    wire N__4961;
    wire N__4960;
    wire N__4959;
    wire N__4958;
    wire N__4955;
    wire N__4950;
    wire N__4949;
    wire N__4948;
    wire N__4947;
    wire N__4942;
    wire N__4939;
    wire N__4934;
    wire N__4929;
    wire N__4926;
    wire N__4921;
    wire N__4918;
    wire N__4913;
    wire N__4910;
    wire N__4905;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4893;
    wire N__4890;
    wire N__4881;
    wire N__4878;
    wire N__4875;
    wire N__4874;
    wire N__4873;
    wire N__4872;
    wire N__4871;
    wire N__4868;
    wire N__4863;
    wire N__4862;
    wire N__4859;
    wire N__4856;
    wire N__4853;
    wire N__4852;
    wire N__4851;
    wire N__4848;
    wire N__4845;
    wire N__4844;
    wire N__4843;
    wire N__4838;
    wire N__4835;
    wire N__4830;
    wire N__4827;
    wire N__4820;
    wire N__4817;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4793;
    wire N__4788;
    wire N__4785;
    wire N__4782;
    wire N__4779;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4771;
    wire N__4770;
    wire N__4769;
    wire N__4768;
    wire N__4765;
    wire N__4762;
    wire N__4757;
    wire N__4752;
    wire N__4743;
    wire N__4742;
    wire N__4741;
    wire N__4740;
    wire N__4739;
    wire N__4730;
    wire N__4727;
    wire N__4726;
    wire N__4725;
    wire N__4724;
    wire N__4723;
    wire N__4720;
    wire N__4717;
    wire N__4712;
    wire N__4709;
    wire N__4706;
    wire N__4705;
    wire N__4702;
    wire N__4695;
    wire N__4692;
    wire N__4689;
    wire N__4684;
    wire N__4679;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4667;
    wire N__4664;
    wire N__4659;
    wire N__4656;
    wire N__4653;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4641;
    wire N__4638;
    wire N__4635;
    wire N__4634;
    wire N__4631;
    wire N__4630;
    wire N__4627;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4617;
    wire N__4614;
    wire N__4611;
    wire N__4608;
    wire N__4603;
    wire N__4600;
    wire N__4597;
    wire N__4594;
    wire N__4591;
    wire N__4588;
    wire N__4585;
    wire N__4582;
    wire N__4579;
    wire N__4576;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4560;
    wire N__4557;
    wire N__4554;
    wire N__4551;
    wire N__4548;
    wire N__4545;
    wire N__4542;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4530;
    wire N__4527;
    wire N__4524;
    wire N__4521;
    wire N__4518;
    wire N__4515;
    wire N__4512;
    wire N__4509;
    wire N__4506;
    wire N__4505;
    wire N__4502;
    wire N__4497;
    wire N__4494;
    wire N__4491;
    wire N__4490;
    wire N__4487;
    wire N__4484;
    wire N__4479;
    wire N__4478;
    wire N__4477;
    wire N__4474;
    wire N__4471;
    wire N__4468;
    wire N__4461;
    wire N__4458;
    wire N__4455;
    wire N__4452;
    wire N__4449;
    wire N__4446;
    wire N__4443;
    wire N__4440;
    wire N__4437;
    wire N__4434;
    wire N__4431;
    wire N__4428;
    wire N__4425;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4407;
    wire N__4404;
    wire N__4401;
    wire N__4398;
    wire N__4397;
    wire N__4394;
    wire N__4391;
    wire N__4388;
    wire N__4385;
    wire N__4382;
    wire N__4379;
    wire N__4374;
    wire N__4371;
    wire N__4368;
    wire N__4365;
    wire N__4362;
    wire N__4359;
    wire N__4356;
    wire N__4353;
    wire N__4350;
    wire N__4347;
    wire N__4344;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4332;
    wire N__4329;
    wire N__4328;
    wire N__4323;
    wire N__4320;
    wire N__4317;
    wire N__4314;
    wire N__4311;
    wire N__4310;
    wire N__4305;
    wire N__4302;
    wire N__4299;
    wire N__4296;
    wire N__4295;
    wire N__4294;
    wire N__4293;
    wire N__4288;
    wire N__4283;
    wire N__4280;
    wire N__4279;
    wire N__4278;
    wire N__4275;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4263;
    wire N__4254;
    wire N__4251;
    wire N__4250;
    wire N__4247;
    wire N__4242;
    wire N__4241;
    wire N__4238;
    wire N__4235;
    wire N__4230;
    wire N__4227;
    wire N__4224;
    wire N__4221;
    wire N__4218;
    wire N__4215;
    wire N__4214;
    wire N__4213;
    wire N__4212;
    wire N__4209;
    wire N__4202;
    wire N__4197;
    wire N__4194;
    wire N__4193;
    wire N__4192;
    wire N__4185;
    wire N__4184;
    wire N__4181;
    wire N__4178;
    wire N__4175;
    wire N__4172;
    wire N__4167;
    wire N__4164;
    wire N__4161;
    wire N__4160;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4137;
    wire N__4136;
    wire N__4131;
    wire N__4128;
    wire N__4125;
    wire N__4122;
    wire N__4119;
    wire N__4118;
    wire N__4113;
    wire N__4110;
    wire N__4107;
    wire N__4104;
    wire N__4101;
    wire N__4098;
    wire N__4095;
    wire N__4092;
    wire N__4089;
    wire N__4086;
    wire N__4083;
    wire N__4080;
    wire N__4077;
    wire N__4074;
    wire N__4071;
    wire N__4068;
    wire N__4065;
    wire N__4062;
    wire N__4059;
    wire N__4056;
    wire N__4053;
    wire N__4050;
    wire N__4047;
    wire N__4044;
    wire N__4041;
    wire N__4038;
    wire N__4035;
    wire N__4032;
    wire N__4031;
    wire N__4030;
    wire N__4029;
    wire N__4028;
    wire N__4027;
    wire N__4026;
    wire N__4025;
    wire N__4024;
    wire N__4023;
    wire N__4022;
    wire N__4021;
    wire N__4020;
    wire N__4019;
    wire N__3990;
    wire CLK80_OUT;
    wire A_c_15;
    wire A_c_14;
    wire GNDG0;
    wire VCCG0;
    wire \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0_a3_0Z0Z_2_cascade_ ;
    wire A_c_7;
    wire A_c_6;
    wire \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4_cascade_ ;
    wire A_c_24;
    wire A_c_26;
    wire A_c_27;
    wire \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_5 ;
    wire \U409_AUTOCONFIG.N_42 ;
    wire \U409_AUTOCONFIG.N_111_cascade_ ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_1_0_cascade_ ;
    wire \U409_AUTOCONFIG.N_62 ;
    wire \U409_ADDRESS_DECODE.N_54_cascade_ ;
    wire A_c_5;
    wire \U409_AUTOCONFIG.N_92 ;
    wire \U409_AUTOCONFIG.N_86_cascade_ ;
    wire \U409_AUTOCONFIG.N_57 ;
    wire N_89_1;
    wire N_89_1_cascade_;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_3 ;
    wire A_c_25;
    wire TT_c_0;
    wire TT_c_1;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_9 ;
    wire \U409_AUTOCONFIG.N_38 ;
    wire \U409_AUTOCONFIG.N_48 ;
    wire \U409_AUTOCONFIG.N_111 ;
    wire \U409_AUTOCONFIG.N_41 ;
    wire \U409_AUTOCONFIG.N_43 ;
    wire \U409_AUTOCONFIG.N_66 ;
    wire \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_i_1_cascade_ ;
    wire \INVU409_AUTOCONFIG.LIDE_OUT_3C_net ;
    wire \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_4 ;
    wire \U409_ADDRESS_DECODE.N_112_cascade_ ;
    wire \U409_ADDRESS_DECODE.N_112 ;
    wire \U409_AUTOCONFIG.N_74_cascade_ ;
    wire \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_i_0 ;
    wire A_c_4;
    wire A_c_2;
    wire \U409_AUTOCONFIG.N_44 ;
    wire \U409_AUTOCONFIG.N_86 ;
    wire A_c_3;
    wire \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_1_85_i_i_0 ;
    wire N_121;
    wire N_121_cascade_;
    wire A_c_16;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_1 ;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_7 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_0 ;
    wire U409_AUTOCONFIG_D_OUT_0_i_0;
    wire \U409_AUTOCONFIG.N_27 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ;
    wire \U409_AUTOCONFIG.N_31 ;
    wire \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ;
    wire \U409_AUTOCONFIG.N_22 ;
    wire \U409_AUTOCONFIG.LIDE_CONF_1_sqmuxa_0_a2_0Z0Z_2 ;
    wire \U409_AUTOCONFIG.N_20 ;
    wire \INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net ;
    wire CPUCONFn_c;
    wire \U409_AUTOCONFIG.N_52 ;
    wire \U409_AUTOCONFIG.N_52_cascade_ ;
    wire \U409_AUTOCONFIG.N_56 ;
    wire \U409_AUTOCONFIG.N_67 ;
    wire \U409_AUTOCONFIG.N_56_cascade_ ;
    wire \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0Z0Z_0 ;
    wire \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa ;
    wire \U409_ADDRESS_DECODE.HIROMZ0 ;
    wire \U409_ADDRESS_DECODE.LOWROMZ0Z_2_cascade_ ;
    wire D_1_i;
    wire \U409_AUTOCONFIG.AC_STARTZ0 ;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2Z0Z_1_cascade_ ;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2Z0Z_4_cascade_ ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_10 ;
    wire N_120_cascade_;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_11 ;
    wire U409_ADDRESS_DECODE_un1_REGSPACEn_i;
    wire \U409_ADDRESS_DECODE.N_102 ;
    wire \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3Z0Z_0 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ;
    wire U409_AUTOCONFIG_D_OUT_0_i_1;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ;
    wire U409_AUTOCONFIG_D_OUT_0_i_2;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ;
    wire U409_AUTOCONFIG_D_OUT_0_i_3;
    wire \U409_AUTOCONFIG.STATEZ0Z_1 ;
    wire \U409_AUTOCONFIG.STATEZ0Z_0 ;
    wire \INVU409_AUTOCONFIG.LIDE_CONFC_net ;
    wire TM_c_0;
    wire CONFIGURED;
    wire TM_c_1;
    wire A_c_17;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1_cascade_ ;
    wire ATA_BASE_1;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_4_cascade_ ;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_ ;
    wire RnW_c;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2Z0Z_4 ;
    wire \U409_ADDRESS_DECODE.Z2_SPACE ;
    wire N_120_i;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1 ;
    wire A_c_31;
    wire N_120;
    wire \U409_ADDRESS_DECODE.PORTSIZEZ0Z_0_cascade_ ;
    wire PORTSIZE_0_i;
    wire A_c_30;
    wire A_c_29;
    wire \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_0 ;
    wire CONFIGENn_c;
    wire D_in_7;
    wire BRIDGE_BASE_3;
    wire BRIDGE_BASE_2;
    wire BRIDGE_BASE_1;
    wire \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa ;
    wire \INVU409_AUTOCONFIG.CONFIGENnC_net ;
    wire A_c_23;
    wire ATA_BASE_7;
    wire A_c_22;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3 ;
    wire A_c_1;
    wire \U409_AUTOCONFIG.LIDE_CONFZ0 ;
    wire \U409_AUTOCONFIG.N_122 ;
    wire A_c_19;
    wire ATA_BASE_3;
    wire A_c_18;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2 ;
    wire A_c_20;
    wire \U409_ADDRESS_DECODE.ATA_SPACE_1Z0Z_0 ;
    wire U409_ADDRESS_DECODE_un1_RAMSPACEn_i;
    wire U409_ADDRESS_DECODE_un1_ROMEN_0;
    wire \U409_ADDRESS_DECODE.ATA_ENZ0 ;
    wire U409_ADDRESS_DECODE_un1_ATA_ENn_i;
    wire \U409_TRANSFER_ACK.CO1 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER20 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0 ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_cascade_ ;
    wire D_in_4;
    wire ATA_BASE_4;
    wire D_in_5;
    wire ATA_BASE_5;
    wire \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42Z0Z_1 ;
    wire ATA_BASE_6;
    wire \INVU409_AUTOCONFIG.ATA_BASE_4C_net ;
    wire un1_AUTOCONFIG_SPACE;
    wire \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42Z0Z_0 ;
    wire D_in_6;
    wire ATA_BASE_2;
    wire \INVU409_AUTOCONFIG.ATA_BASE_2C_net ;
    wire \U409_ADDRESS_DECODE.LOWROMZ0Z_3 ;
    wire U409_ADDRESS_DECODE_ROMEN_1;
    wire A_c_21;
    wire OVL_c;
    wire \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ;
    wire A_c_28;
    wire BRIDGE_BASE_0;
    wire \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_3 ;
    wire U409_ADDRESS_DECODE_un1_BRIDGE_ENn_i;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ;
    wire ROMENn_c;
    wire \INVU409_TRANSFER_ACK.ROMENn_nessC_net ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_0 ;
    wire \INVU409_TRANSFER_ACK.TACK_ENC_net ;
    wire \INVU409_TRANSFER_ACK.TACK_OUTnC_net ;
    wire AC_TACK;
    wire \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_ ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER6 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ;
    wire TACK_OUTn;
    wire \U409_TRANSFER_ACK.TACK_OUTn_3_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER20_2 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ;
    wire TACKn_in;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0 ;
    wire U409_ADDRESS_DECODE_un1_REGSPACEn;
    wire U409_ADDRESS_DECODE_un1_RAMSPACEn;
    wire BUFENn_c;
    wire \U409_TRANSFER_ACK.N_119 ;
    wire GB_BUFFER_CLK40_IN_c_g_THRU_CO;
    wire CONSTANT_ONE_NET;
    wire \U409_TRANSFER_ACK.N_17_mux_cascade_ ;
    wire \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_ ;
    wire \U409_TRANSFER_ACK.N_6_0_cascade_ ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_0C_net ;
    wire \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0 ;
    wire \U409_TRANSFER_ACK.N_3_0 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ;
    wire \U409_TRANSFER_ACK.N_17_mux ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a3_3 ;
    wire \U409_TRANSFER_ACK.N_87_cascade_ ;
    wire \U409_TRANSFER_ACK.N_77 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ;
    wire TSn_c;
    wire CLK40_IN_c_g;
    wire \U409_TRANSFER_ACK.N_87 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ;
    wire RESETn_c_i;
    wire bfn_13_6_0_;
    wire \U409_TICK.un3_COUNTER60_1_cry_1 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_2 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_3 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_4 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_6 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_8 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_9 ;
    wire bfn_13_7_0_;
    wire \U409_TICK.un3_COUNTER60_1_cry_9 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_10 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_13 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_15 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_6 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_4 ;
    wire \U409_TICK.COUNTER60Z0Z_12 ;
    wire \U409_TICK.COUNTER60Z0Z_2 ;
    wire \U409_TICK.COUNTER60Z0Z_16 ;
    wire \U409_TICK.COUNTER60Z0Z_1 ;
    wire \U409_TICK.COUNTER60Z0Z_7 ;
    wire \U409_TICK.COUNTER60Z0Z_10 ;
    wire \U409_TICK.COUNTER60Z0Z_13 ;
    wire \U409_TICK.COUNTER60Z0Z_15 ;
    wire \U409_TICK.COUNTER60Z0Z_5 ;
    wire \U409_TICK.COUNTER60Z0Z_4 ;
    wire \U409_TICK.TICK603_11 ;
    wire \U409_TICK.COUNTER60Z0Z_11 ;
    wire \U409_TICK.TICK603_8_cascade_ ;
    wire \U409_TICK.COUNTER60Z0Z_3 ;
    wire \U409_TICK.TICK603_14_cascade_ ;
    wire \U409_TICK.COUNTER60Z0Z_0 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_1 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_0 ;
    wire \INVU409_TRANSFER_ACK.LASTCLK_1C_net ;
    wire RESETn_c_i_g;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ;
    wire \U409_TICK.COUNTER50Z0Z_1 ;
    wire bfn_14_5_0_;
    wire \U409_TICK.COUNTER50Z0Z_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_1 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_3 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_4 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_6 ;
    wire \U409_TICK.COUNTER50Z0Z_8 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_8 ;
    wire bfn_14_6_0_;
    wire \U409_TICK.un2_COUNTER50_1_cry_9 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_10 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_11 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_13 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_15 ;
    wire \U409_TICK.COUNTER50Z0Z_16 ;
    wire \U409_CIA.CLK_CIA_r_1_0_cascade_ ;
    wire CLK_CIA_c;
    wire \U409_TICK.COUNTER50Z0Z_5 ;
    wire \U409_TICK.COUNTER50Z0Z_3 ;
    wire \U409_TICK.COUNTER50Z0Z_0 ;
    wire \U409_TICK.COUNTER50Z0Z_10 ;
    wire \U409_TICK.TICK503_11 ;
    wire \U409_TICK.TICK503_8_cascade_ ;
    wire \U409_TICK.COUNTER50Z0Z_12 ;
    wire \U409_TICK.COUNTER60Z0Z_9 ;
    wire \U409_TICK.COUNTER60Z0Z_6 ;
    wire \U409_TICK.TICK603_9_cascade_ ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_14 ;
    wire \U409_TICK.COUNTER60Z0Z_14 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_9 ;
    wire TICK50_c;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_8 ;
    wire \U409_TICK.COUNTER60Z0Z_8 ;
    wire \U409_TICK.TICK603_14 ;
    wire \U409_TICK.TICK603_10 ;
    wire \U409_TICK.TICK603_9 ;
    wire TICK60_c;
    wire \U409_TICK.COUNTER50Z0Z_9 ;
    wire \U409_TICK.TICK503_9_cascade_ ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_6 ;
    wire \U409_TICK.COUNTER50Z0Z_6 ;
    wire \U409_TICK.COUNTER50Z0Z_7 ;
    wire \U409_TICK.COUNTER50Z0Z_4 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_13 ;
    wire \U409_TICK.COUNTER50Z0Z_13 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER50Z0Z_15 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_14 ;
    wire \U409_TICK.COUNTER50Z0Z_14 ;
    wire \U409_TICK.TICK503_10 ;
    wire \U409_TICK.TICK503_14 ;
    wire \U409_TICK.TICK503_9 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_11 ;
    wire \U409_TICK.COUNTER50Z0Z_11 ;
    wire CLK6_c_g;
    wire \U409_CIA.CLK_CIA6_3 ;
    wire \U409_CIA.CIA_CLK_COUNT11_3_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNT11_2_0 ;
    wire \U409_CIA.CIA_CLK_COUNT11_3 ;
    wire \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_ ;
    wire \U409_CIA.CLK_CIA6_4_cascade_ ;
    wire \U409_CIA.VMA_RNOZ0Z_0_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_1 ;
    wire bfn_16_7_0_;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_1 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_4 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_6 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_5 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_6 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_7 ;
    wire CLK28_IN_c_g;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_3 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_2 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_5 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_0 ;
    wire \U409_CIA.un1_CIA_CLK_COUNT_3_2 ;
    wire TACK_EN;
    wire AUTOCONFIG_SPACE;
    wire CIA_SPACE;
    wire TCIn_1_i;
    wire RESETn_c;
    wire \U409_CIA.VMAZ0 ;
    wire A_c_12;
    wire U409_ADDRESS_DECODE_un1_CIACS0n_i;
    wire CIA_ENABLE;
    wire A_c_13;
    wire U409_ADDRESS_DECODE_un1_CIACS1n_i;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="SIMPLE";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0001111;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE pll (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__7680),
            .RESETB(N__7665),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(CLK80_OUT));
    PRE_IO_GBUF CLK28_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__11322),
            .GLOBALBUFFEROUTPUT(CLK28_IN_c_g));
    IO_PAD CLK28_IN_ibuf_gb_io_iopad (
            .OE(N__11324),
            .DIN(N__11323),
            .DOUT(N__11322),
            .PACKAGEPIN(CLK28_IN));
    defparam CLK28_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK28_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK28_IN_ibuf_gb_io_preio (
            .PADOEN(N__11324),
            .PADOUT(N__11323),
            .PADIN(N__11322),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK6_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__11312),
            .GLOBALBUFFEROUTPUT(CLK6_c_g));
    IO_PAD CLK6_ibuf_gb_io_iopad (
            .OE(N__11314),
            .DIN(N__11313),
            .DOUT(N__11312),
            .PACKAGEPIN(CLK6));
    defparam CLK6_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK6_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK6_ibuf_gb_io_preio (
            .PADOEN(N__11314),
            .PADOUT(N__11313),
            .PADIN(N__11312),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK40_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__11302),
            .GLOBALBUFFEROUTPUT(CLK40_IN_c_g));
    IO_PAD CLK40_IN_ibuf_gb_io_iopad (
            .OE(N__11304),
            .DIN(N__11303),
            .DOUT(N__11302),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_gb_io_preio (
            .PADOEN(N__11304),
            .PADOUT(N__11303),
            .PADIN(N__11302),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__11293),
            .DIN(N__11292),
            .DOUT(N__11291),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__11293),
            .PADOUT(N__11292),
            .PADIN(N__11291),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_0_iopad (
            .OE(N__11284),
            .DIN(N__11283),
            .DOUT(N__11282),
            .PACKAGEPIN(TT[0]));
    defparam TT_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_0_preio (
            .PADOEN(N__11284),
            .PADOUT(N__11283),
            .PADIN(N__11282),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_P1_obuf_iopad (
            .OE(N__11275),
            .DIN(N__11274),
            .DOUT(N__11273),
            .PACKAGEPIN(PIO_P1));
    defparam PIO_P1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_P1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_P1_obuf_preio (
            .PADOEN(N__11275),
            .PADOUT(N__11274),
            .PADIN(N__11273),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10647),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_7_iopad (
            .OE(N__11266),
            .DIN(N__11265),
            .DOUT(N__11264),
            .PACKAGEPIN(D[7]));
    defparam D_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_7_preio (
            .PADOEN(N__11266),
            .PADOUT(N__11265),
            .PADIN(N__11264),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5160),
            .DIN0(D_in_7),
            .DOUT0(N__5223),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__11257),
            .DIN(N__11256),
            .DOUT(N__11255),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__11257),
            .PADOUT(N__11256),
            .PADIN(N__11255),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CPUCONFn_ibuf_iopad (
            .OE(N__11248),
            .DIN(N__11247),
            .DOUT(N__11246),
            .PACKAGEPIN(CPUCONFn));
    defparam CPUCONFn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CPUCONFn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CPUCONFn_ibuf_preio (
            .PADOEN(N__11248),
            .PADOUT(N__11247),
            .PADIN(N__11246),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CPUCONFn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RTC_ENn_obuf_iopad (
            .OE(N__11239),
            .DIN(N__11238),
            .DOUT(N__11237),
            .PACKAGEPIN(RTC_ENn));
    defparam RTC_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RTC_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RTC_ENn_obuf_preio (
            .PADOEN(N__11239),
            .PADOUT(N__11238),
            .PADIN(N__11237),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5427),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_24_iopad (
            .OE(N__11230),
            .DIN(N__11229),
            .DOUT(N__11228),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__11230),
            .PADOUT(N__11229),
            .PADIN(N__11228),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_4_iopad (
            .OE(N__11221),
            .DIN(N__11220),
            .DOUT(N__11219),
            .PACKAGEPIN(D[4]));
    defparam D_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_4_preio (
            .PADOEN(N__11221),
            .PADOUT(N__11220),
            .PADIN(N__11219),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5135),
            .DIN0(D_in_4),
            .DOUT0(N__4530),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__11212),
            .DIN(N__11211),
            .DOUT(N__11210),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__11212),
            .PADOUT(N__11211),
            .PADIN(N__11210),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TM_ibuf_1_iopad (
            .OE(N__11203),
            .DIN(N__11202),
            .DOUT(N__11201),
            .PACKAGEPIN(TM[1]));
    defparam TM_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TM_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TM_ibuf_1_preio (
            .PADOEN(N__11203),
            .PADOUT(N__11202),
            .PADIN(N__11201),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TM_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_21_iopad (
            .OE(N__11194),
            .DIN(N__11193),
            .DOUT(N__11192),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__11194),
            .PADOUT(N__11193),
            .PADIN(N__11192),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_obuf_iopad (
            .OE(N__11185),
            .DIN(N__11184),
            .DOUT(N__11183),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMSPACEn_obuf_preio (
            .PADOEN(N__11185),
            .PADOUT(N__11184),
            .PADIN(N__11183),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6840),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__11176),
            .DIN(N__11175),
            .DOUT(N__11174),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__11176),
            .PADOUT(N__11175),
            .PADIN(N__11174),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ROMENn_obuf_iopad (
            .OE(N__11167),
            .DIN(N__11166),
            .DOUT(N__11165),
            .PACKAGEPIN(ROMENn));
    defparam ROMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ROMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ROMENn_obuf_preio (
            .PADOEN(N__11167),
            .PADOUT(N__11166),
            .PADIN(N__11165),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7578),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuft_iopad (
            .OE(N__11158),
            .DIN(N__11157),
            .DOUT(N__11156),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TBIn_obuft_preio (
            .PADOEN(N__11158),
            .PADOUT(N__11157),
            .PADIN(N__11156),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10359),
            .DIN0(),
            .DOUT0(N__7982),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__11149),
            .DIN(N__11148),
            .DOUT(N__11147),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__11149),
            .PADOUT(N__11148),
            .PADIN(N__11147),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORTSIZE_obuf_iopad (
            .OE(N__11140),
            .DIN(N__11139),
            .DOUT(N__11138),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PORTSIZE_obuf_preio (
            .PADOEN(N__11140),
            .PADOUT(N__11139),
            .PADIN(N__11138),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5928),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_P2_obuf_iopad (
            .OE(N__11131),
            .DIN(N__11130),
            .DOUT(N__11129),
            .PACKAGEPIN(PIO_P2));
    defparam PIO_P2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_P2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_P2_obuf_preio (
            .PADOEN(N__11131),
            .PADOUT(N__11130),
            .PADIN(N__11129),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4056),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__11122),
            .DIN(N__11121),
            .DOUT(N__11120),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__11122),
            .PADOUT(N__11121),
            .PADIN(N__11120),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BRIDGE_ENn_obuf_iopad (
            .OE(N__11113),
            .DIN(N__11112),
            .DOUT(N__11111),
            .PACKAGEPIN(BRIDGE_ENn));
    defparam BRIDGE_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BRIDGE_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BRIDGE_ENn_obuf_preio (
            .PADOEN(N__11113),
            .PADOUT(N__11112),
            .PADIN(N__11111),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6957),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_22_iopad (
            .OE(N__11104),
            .DIN(N__11103),
            .DOUT(N__11102),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__11104),
            .PADOUT(N__11103),
            .PADIN(N__11102),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__11095),
            .DIN(N__11094),
            .DOUT(N__11093),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__11095),
            .PADOUT(N__11094),
            .PADIN(N__11093),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__11086),
            .DIN(N__11085),
            .DOUT(N__11084),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__11086),
            .PADOUT(N__11085),
            .PADIN(N__11084),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__11077),
            .DIN(N__11076),
            .DOUT(N__11075),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__11077),
            .PADOUT(N__11076),
            .PADIN(N__11075),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__11068),
            .DIN(N__11067),
            .DOUT(N__11066),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__11068),
            .PADOUT(N__11067),
            .PADIN(N__11066),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_25_iopad (
            .OE(N__11059),
            .DIN(N__11058),
            .DOUT(N__11057),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__11059),
            .PADOUT(N__11058),
            .PADIN(N__11057),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS0n_obuf_iopad (
            .OE(N__11050),
            .DIN(N__11049),
            .DOUT(N__11048),
            .PACKAGEPIN(CIACS0n));
    defparam CIACS0n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS0n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS0n_obuf_preio (
            .PADOEN(N__11050),
            .PADOUT(N__11049),
            .PADIN(N__11048),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10674),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK50_obuf_iopad (
            .OE(N__11041),
            .DIN(N__11040),
            .DOUT(N__11039),
            .PACKAGEPIN(TICK50));
    defparam TICK50_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK50_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK50_obuf_preio (
            .PADOEN(N__11041),
            .PADOUT(N__11040),
            .PADIN(N__11039),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9459),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__11032),
            .DIN(N__11031),
            .DOUT(N__11030),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__11032),
            .PADOUT(N__11031),
            .PADIN(N__11030),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_28_iopad (
            .OE(N__11023),
            .DIN(N__11022),
            .DOUT(N__11021),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__11023),
            .PADOUT(N__11022),
            .PADIN(N__11021),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_30_iopad (
            .OE(N__11014),
            .DIN(N__11013),
            .DOUT(N__11012),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__11014),
            .PADOUT(N__11013),
            .PADIN(N__11012),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD OVL_ibuf_iopad (
            .OE(N__11005),
            .DIN(N__11004),
            .DOUT(N__11003),
            .PACKAGEPIN(OVL));
    defparam OVL_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam OVL_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO OVL_ibuf_preio (
            .PADOEN(N__11005),
            .PADOUT(N__11004),
            .PADIN(N__11003),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(OVL_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuft_iopad (
            .OE(N__10996),
            .DIN(N__10995),
            .DOUT(N__10994),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TCIn_obuft_preio (
            .PADOEN(N__10996),
            .PADOUT(N__10995),
            .PADIN(N__10994),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10212),
            .DIN0(),
            .DOUT0(N__7983),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_5_iopad (
            .OE(N__10987),
            .DIN(N__10986),
            .DOUT(N__10985),
            .PACKAGEPIN(D[5]));
    defparam D_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_5_preio (
            .PADOEN(N__10987),
            .PADOUT(N__10986),
            .PADIN(N__10985),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5155),
            .DIN0(D_in_5),
            .DOUT0(N__5316),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__10978),
            .DIN(N__10977),
            .DOUT(N__10976),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__10978),
            .PADOUT(N__10977),
            .PADIN(N__10976),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__10969),
            .DIN(N__10968),
            .DOUT(N__10967),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__10969),
            .PADOUT(N__10968),
            .PADIN(N__10967),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__10960),
            .DIN(N__10959),
            .DOUT(N__10958),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__10960),
            .PADOUT(N__10959),
            .PADIN(N__10958),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CONFIGENn_obuf_iopad (
            .OE(N__10951),
            .DIN(N__10950),
            .DOUT(N__10949),
            .PACKAGEPIN(CONFIGENn));
    defparam CONFIGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CONFIGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CONFIGENn_obuf_preio (
            .PADOEN(N__10951),
            .PADOUT(N__10950),
            .PADIN(N__10949),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5814),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK60_obuf_iopad (
            .OE(N__10942),
            .DIN(N__10941),
            .DOUT(N__10940),
            .PACKAGEPIN(TICK60));
    defparam TICK60_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK60_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK60_obuf_preio (
            .PADOEN(N__10942),
            .PADOUT(N__10941),
            .PADIN(N__10940),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9291),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_26_iopad (
            .OE(N__10933),
            .DIN(N__10932),
            .DOUT(N__10931),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__10933),
            .PADOUT(N__10932),
            .PADIN(N__10931),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_P0_obuf_iopad (
            .OE(N__10924),
            .DIN(N__10923),
            .DOUT(N__10922),
            .PACKAGEPIN(PIO_P0));
    defparam PIO_P0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_P0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_P0_obuf_preio (
            .PADOEN(N__10924),
            .PADOUT(N__10923),
            .PADIN(N__10922),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10716),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_23_iopad (
            .OE(N__10915),
            .DIN(N__10914),
            .DOUT(N__10913),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__10915),
            .PADOUT(N__10914),
            .PADIN(N__10913),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__10906),
            .DIN(N__10905),
            .DOUT(N__10904),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__10906),
            .PADOUT(N__10905),
            .PADIN(N__10904),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ATA_ENn_obuf_iopad (
            .OE(N__10897),
            .DIN(N__10896),
            .DOUT(N__10895),
            .PACKAGEPIN(ATA_ENn));
    defparam ATA_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ATA_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ATA_ENn_obuf_preio (
            .PADOEN(N__10897),
            .PADOUT(N__10896),
            .PADIN(N__10895),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6789),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_31_iopad (
            .OE(N__10888),
            .DIN(N__10887),
            .DOUT(N__10886),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__10888),
            .PADOUT(N__10887),
            .PADIN(N__10886),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS1n_obuf_iopad (
            .OE(N__10879),
            .DIN(N__10878),
            .DOUT(N__10877),
            .PACKAGEPIN(CIACS1n));
    defparam CIACS1n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS1n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS1n_obuf_preio (
            .PADOEN(N__10879),
            .PADOUT(N__10878),
            .PADIN(N__10877),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10611),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_obuf_iopad (
            .OE(N__10870),
            .DIN(N__10869),
            .DOUT(N__10868),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGSPACEn_obuf_preio (
            .PADOEN(N__10870),
            .PADOUT(N__10869),
            .PADIN(N__10868),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5400),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__10861),
            .DIN(N__10860),
            .DOUT(N__10859),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__10861),
            .PADOUT(N__10860),
            .PADIN(N__10859),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_CIA_obuf_iopad (
            .OE(N__10852),
            .DIN(N__10851),
            .DOUT(N__10850),
            .PACKAGEPIN(CLK_CIA));
    defparam CLK_CIA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_CIA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_CIA_obuf_preio (
            .PADOEN(N__10852),
            .PADOUT(N__10851),
            .PADIN(N__10850),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9213),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__10843),
            .DIN(N__10842),
            .DOUT(N__10841),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__10843),
            .PADOUT(N__10842),
            .PADIN(N__10841),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__10834),
            .DIN(N__10833),
            .DOUT(N__10832),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__10834),
            .PADOUT(N__10833),
            .PADIN(N__10832),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10355),
            .DIN0(TACKn_in),
            .DOUT0(N__7975),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_1_iopad (
            .OE(N__10825),
            .DIN(N__10824),
            .DOUT(N__10823),
            .PACKAGEPIN(TT[1]));
    defparam TT_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_1_preio (
            .PADOEN(N__10825),
            .PADOUT(N__10824),
            .PADIN(N__10823),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__10816),
            .DIN(N__10815),
            .DOUT(N__10814),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__10816),
            .PADOUT(N__10815),
            .PADIN(N__10814),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7704),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_S0_obuf_iopad (
            .OE(N__10807),
            .DIN(N__10806),
            .DOUT(N__10805),
            .PACKAGEPIN(PIO_S0));
    defparam PIO_S0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_S0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_S0_obuf_preio (
            .PADOEN(N__10807),
            .PADOUT(N__10806),
            .PADIN(N__10805),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4080),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_29_iopad (
            .OE(N__10798),
            .DIN(N__10797),
            .DOUT(N__10796),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__10798),
            .PADOUT(N__10797),
            .PADIN(N__10796),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_S2_obuf_iopad (
            .OE(N__10789),
            .DIN(N__10788),
            .DOUT(N__10787),
            .PACKAGEPIN(PIO_S2));
    defparam PIO_S2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_S2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_S2_obuf_preio (
            .PADOEN(N__10789),
            .PADOUT(N__10788),
            .PADIN(N__10787),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7664),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_6_iopad (
            .OE(N__10780),
            .DIN(N__10779),
            .DOUT(N__10778),
            .PACKAGEPIN(D[6]));
    defparam D_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_6_preio (
            .PADOEN(N__10780),
            .PADOUT(N__10779),
            .PADIN(N__10778),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5156),
            .DIN0(D_in_6),
            .DOUT0(N__5268),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__10771),
            .DIN(N__10770),
            .DOUT(N__10769),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__10771),
            .PADOUT(N__10770),
            .PADIN(N__10769),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_27_iopad (
            .OE(N__10762),
            .DIN(N__10761),
            .DOUT(N__10760),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__10762),
            .PADOUT(N__10761),
            .PADIN(N__10760),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_S1_obuf_iopad (
            .OE(N__10753),
            .DIN(N__10752),
            .DOUT(N__10751),
            .PACKAGEPIN(PIO_S1));
    defparam PIO_S1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_S1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_S1_obuf_preio (
            .PADOEN(N__10753),
            .PADOUT(N__10752),
            .PADIN(N__10751),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4638),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TM_ibuf_0_iopad (
            .OE(N__10744),
            .DIN(N__10743),
            .DOUT(N__10742),
            .PACKAGEPIN(TM[0]));
    defparam TM_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TM_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TM_ibuf_0_preio (
            .PADOEN(N__10744),
            .PADOUT(N__10743),
            .PADIN(N__10742),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TM_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__10735),
            .DIN(N__10734),
            .DOUT(N__10733),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__10735),
            .PADOUT(N__10734),
            .PADIN(N__10733),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IoInMux I__2593 (
            .O(N__10716),
            .I(N__10713));
    LocalMux I__2592 (
            .O(N__10713),
            .I(N__10710));
    Span4Mux_s0_h I__2591 (
            .O(N__10710),
            .I(N__10706));
    InMux I__2590 (
            .O(N__10709),
            .I(N__10703));
    Sp12to4 I__2589 (
            .O(N__10706),
            .I(N__10700));
    LocalMux I__2588 (
            .O(N__10703),
            .I(N__10697));
    Span12Mux_s10_v I__2587 (
            .O(N__10700),
            .I(N__10694));
    Span12Mux_s10_v I__2586 (
            .O(N__10697),
            .I(N__10691));
    Span12Mux_h I__2585 (
            .O(N__10694),
            .I(N__10688));
    Span12Mux_h I__2584 (
            .O(N__10691),
            .I(N__10685));
    Span12Mux_h I__2583 (
            .O(N__10688),
            .I(N__10682));
    Span12Mux_h I__2582 (
            .O(N__10685),
            .I(N__10679));
    Odrv12 I__2581 (
            .O(N__10682),
            .I(A_c_12));
    Odrv12 I__2580 (
            .O(N__10679),
            .I(A_c_12));
    IoInMux I__2579 (
            .O(N__10674),
            .I(N__10671));
    LocalMux I__2578 (
            .O(N__10671),
            .I(N__10668));
    Span4Mux_s3_h I__2577 (
            .O(N__10668),
            .I(N__10665));
    Span4Mux_v I__2576 (
            .O(N__10665),
            .I(N__10662));
    Odrv4 I__2575 (
            .O(N__10662),
            .I(U409_ADDRESS_DECODE_un1_CIACS0n_i));
    InMux I__2574 (
            .O(N__10659),
            .I(N__10653));
    InMux I__2573 (
            .O(N__10658),
            .I(N__10653));
    LocalMux I__2572 (
            .O(N__10653),
            .I(N__10650));
    Odrv12 I__2571 (
            .O(N__10650),
            .I(CIA_ENABLE));
    IoInMux I__2570 (
            .O(N__10647),
            .I(N__10644));
    LocalMux I__2569 (
            .O(N__10644),
            .I(N__10641));
    IoSpan4Mux I__2568 (
            .O(N__10641),
            .I(N__10637));
    InMux I__2567 (
            .O(N__10640),
            .I(N__10634));
    IoSpan4Mux I__2566 (
            .O(N__10637),
            .I(N__10631));
    LocalMux I__2565 (
            .O(N__10634),
            .I(N__10628));
    Span4Mux_s3_h I__2564 (
            .O(N__10631),
            .I(N__10623));
    Span4Mux_v I__2563 (
            .O(N__10628),
            .I(N__10623));
    Sp12to4 I__2562 (
            .O(N__10623),
            .I(N__10620));
    Span12Mux_h I__2561 (
            .O(N__10620),
            .I(N__10617));
    Span12Mux_h I__2560 (
            .O(N__10617),
            .I(N__10614));
    Odrv12 I__2559 (
            .O(N__10614),
            .I(A_c_13));
    IoInMux I__2558 (
            .O(N__10611),
            .I(N__10608));
    LocalMux I__2557 (
            .O(N__10608),
            .I(N__10605));
    Span4Mux_s3_h I__2556 (
            .O(N__10605),
            .I(N__10602));
    Span4Mux_v I__2555 (
            .O(N__10602),
            .I(N__10599));
    Odrv4 I__2554 (
            .O(N__10599),
            .I(U409_ADDRESS_DECODE_un1_CIACS1n_i));
    InMux I__2553 (
            .O(N__10596),
            .I(N__10593));
    LocalMux I__2552 (
            .O(N__10593),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ));
    InMux I__2551 (
            .O(N__10590),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ));
    InMux I__2550 (
            .O(N__10587),
            .I(N__10584));
    LocalMux I__2549 (
            .O(N__10584),
            .I(N__10578));
    InMux I__2548 (
            .O(N__10583),
            .I(N__10575));
    InMux I__2547 (
            .O(N__10582),
            .I(N__10572));
    InMux I__2546 (
            .O(N__10581),
            .I(N__10569));
    Odrv4 I__2545 (
            .O(N__10578),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__2544 (
            .O(N__10575),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__2543 (
            .O(N__10572),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__2542 (
            .O(N__10569),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    InMux I__2541 (
            .O(N__10560),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ));
    InMux I__2540 (
            .O(N__10557),
            .I(N__10554));
    LocalMux I__2539 (
            .O(N__10554),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO ));
    InMux I__2538 (
            .O(N__10551),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ));
    InMux I__2537 (
            .O(N__10548),
            .I(N__10542));
    InMux I__2536 (
            .O(N__10547),
            .I(N__10539));
    InMux I__2535 (
            .O(N__10546),
            .I(N__10536));
    InMux I__2534 (
            .O(N__10545),
            .I(N__10533));
    LocalMux I__2533 (
            .O(N__10542),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__2532 (
            .O(N__10539),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__2531 (
            .O(N__10536),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__2530 (
            .O(N__10533),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    InMux I__2529 (
            .O(N__10524),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ));
    InMux I__2528 (
            .O(N__10521),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ));
    CascadeMux I__2527 (
            .O(N__10518),
            .I(N__10512));
    CascadeMux I__2526 (
            .O(N__10517),
            .I(N__10509));
    InMux I__2525 (
            .O(N__10516),
            .I(N__10506));
    InMux I__2524 (
            .O(N__10515),
            .I(N__10503));
    InMux I__2523 (
            .O(N__10512),
            .I(N__10498));
    InMux I__2522 (
            .O(N__10509),
            .I(N__10498));
    LocalMux I__2521 (
            .O(N__10506),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    LocalMux I__2520 (
            .O(N__10503),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    LocalMux I__2519 (
            .O(N__10498),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    ClkMux I__2518 (
            .O(N__10491),
            .I(N__10479));
    ClkMux I__2517 (
            .O(N__10490),
            .I(N__10479));
    ClkMux I__2516 (
            .O(N__10489),
            .I(N__10479));
    ClkMux I__2515 (
            .O(N__10488),
            .I(N__10479));
    GlobalMux I__2514 (
            .O(N__10479),
            .I(N__10476));
    gio2CtrlBuf I__2513 (
            .O(N__10476),
            .I(CLK28_IN_c_g));
    InMux I__2512 (
            .O(N__10473),
            .I(N__10466));
    InMux I__2511 (
            .O(N__10472),
            .I(N__10461));
    InMux I__2510 (
            .O(N__10471),
            .I(N__10461));
    InMux I__2509 (
            .O(N__10470),
            .I(N__10456));
    InMux I__2508 (
            .O(N__10469),
            .I(N__10456));
    LocalMux I__2507 (
            .O(N__10466),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__2506 (
            .O(N__10461),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__2505 (
            .O(N__10456),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    InMux I__2504 (
            .O(N__10449),
            .I(N__10446));
    LocalMux I__2503 (
            .O(N__10446),
            .I(N__10440));
    InMux I__2502 (
            .O(N__10445),
            .I(N__10437));
    InMux I__2501 (
            .O(N__10444),
            .I(N__10432));
    InMux I__2500 (
            .O(N__10443),
            .I(N__10432));
    Odrv4 I__2499 (
            .O(N__10440),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__2498 (
            .O(N__10437),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__2497 (
            .O(N__10432),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    CascadeMux I__2496 (
            .O(N__10425),
            .I(N__10419));
    CascadeMux I__2495 (
            .O(N__10424),
            .I(N__10415));
    InMux I__2494 (
            .O(N__10423),
            .I(N__10412));
    InMux I__2493 (
            .O(N__10422),
            .I(N__10407));
    InMux I__2492 (
            .O(N__10419),
            .I(N__10407));
    InMux I__2491 (
            .O(N__10418),
            .I(N__10402));
    InMux I__2490 (
            .O(N__10415),
            .I(N__10402));
    LocalMux I__2489 (
            .O(N__10412),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__2488 (
            .O(N__10407),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__2487 (
            .O(N__10402),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    CascadeMux I__2486 (
            .O(N__10395),
            .I(N__10387));
    InMux I__2485 (
            .O(N__10394),
            .I(N__10384));
    InMux I__2484 (
            .O(N__10393),
            .I(N__10377));
    InMux I__2483 (
            .O(N__10392),
            .I(N__10377));
    InMux I__2482 (
            .O(N__10391),
            .I(N__10377));
    InMux I__2481 (
            .O(N__10390),
            .I(N__10372));
    InMux I__2480 (
            .O(N__10387),
            .I(N__10372));
    LocalMux I__2479 (
            .O(N__10384),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__2478 (
            .O(N__10377),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__2477 (
            .O(N__10372),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    InMux I__2476 (
            .O(N__10365),
            .I(N__10362));
    LocalMux I__2475 (
            .O(N__10362),
            .I(\U409_CIA.un1_CIA_CLK_COUNT_3_2 ));
    IoInMux I__2474 (
            .O(N__10359),
            .I(N__10356));
    LocalMux I__2473 (
            .O(N__10356),
            .I(N__10352));
    IoInMux I__2472 (
            .O(N__10355),
            .I(N__10349));
    IoSpan4Mux I__2471 (
            .O(N__10352),
            .I(N__10346));
    LocalMux I__2470 (
            .O(N__10349),
            .I(N__10343));
    Span4Mux_s0_v I__2469 (
            .O(N__10346),
            .I(N__10338));
    Span4Mux_s0_v I__2468 (
            .O(N__10343),
            .I(N__10338));
    Span4Mux_v I__2467 (
            .O(N__10338),
            .I(N__10334));
    InMux I__2466 (
            .O(N__10337),
            .I(N__10331));
    Sp12to4 I__2465 (
            .O(N__10334),
            .I(N__10328));
    LocalMux I__2464 (
            .O(N__10331),
            .I(N__10325));
    Span12Mux_s9_h I__2463 (
            .O(N__10328),
            .I(N__10321));
    Span4Mux_v I__2462 (
            .O(N__10325),
            .I(N__10318));
    CascadeMux I__2461 (
            .O(N__10324),
            .I(N__10315));
    Span12Mux_v I__2460 (
            .O(N__10321),
            .I(N__10312));
    Span4Mux_h I__2459 (
            .O(N__10318),
            .I(N__10309));
    InMux I__2458 (
            .O(N__10315),
            .I(N__10306));
    Odrv12 I__2457 (
            .O(N__10312),
            .I(TACK_EN));
    Odrv4 I__2456 (
            .O(N__10309),
            .I(TACK_EN));
    LocalMux I__2455 (
            .O(N__10306),
            .I(TACK_EN));
    InMux I__2454 (
            .O(N__10299),
            .I(N__10296));
    LocalMux I__2453 (
            .O(N__10296),
            .I(N__10292));
    InMux I__2452 (
            .O(N__10295),
            .I(N__10289));
    Span4Mux_h I__2451 (
            .O(N__10292),
            .I(N__10283));
    LocalMux I__2450 (
            .O(N__10289),
            .I(N__10283));
    InMux I__2449 (
            .O(N__10288),
            .I(N__10280));
    Span4Mux_h I__2448 (
            .O(N__10283),
            .I(N__10276));
    LocalMux I__2447 (
            .O(N__10280),
            .I(N__10273));
    InMux I__2446 (
            .O(N__10279),
            .I(N__10270));
    Span4Mux_h I__2445 (
            .O(N__10276),
            .I(N__10265));
    Span4Mux_v I__2444 (
            .O(N__10273),
            .I(N__10260));
    LocalMux I__2443 (
            .O(N__10270),
            .I(N__10260));
    InMux I__2442 (
            .O(N__10269),
            .I(N__10255));
    InMux I__2441 (
            .O(N__10268),
            .I(N__10255));
    Odrv4 I__2440 (
            .O(N__10265),
            .I(AUTOCONFIG_SPACE));
    Odrv4 I__2439 (
            .O(N__10260),
            .I(AUTOCONFIG_SPACE));
    LocalMux I__2438 (
            .O(N__10255),
            .I(AUTOCONFIG_SPACE));
    InMux I__2437 (
            .O(N__10248),
            .I(N__10245));
    LocalMux I__2436 (
            .O(N__10245),
            .I(N__10242));
    Span4Mux_v I__2435 (
            .O(N__10242),
            .I(N__10239));
    Span4Mux_v I__2434 (
            .O(N__10239),
            .I(N__10235));
    InMux I__2433 (
            .O(N__10238),
            .I(N__10232));
    Sp12to4 I__2432 (
            .O(N__10235),
            .I(N__10226));
    LocalMux I__2431 (
            .O(N__10232),
            .I(N__10226));
    InMux I__2430 (
            .O(N__10231),
            .I(N__10223));
    Span12Mux_h I__2429 (
            .O(N__10226),
            .I(N__10220));
    LocalMux I__2428 (
            .O(N__10223),
            .I(N__10217));
    Odrv12 I__2427 (
            .O(N__10220),
            .I(CIA_SPACE));
    Odrv4 I__2426 (
            .O(N__10217),
            .I(CIA_SPACE));
    IoInMux I__2425 (
            .O(N__10212),
            .I(N__10209));
    LocalMux I__2424 (
            .O(N__10209),
            .I(N__10206));
    Span4Mux_s1_v I__2423 (
            .O(N__10206),
            .I(N__10203));
    Sp12to4 I__2422 (
            .O(N__10203),
            .I(N__10200));
    Span12Mux_h I__2421 (
            .O(N__10200),
            .I(N__10197));
    Span12Mux_v I__2420 (
            .O(N__10197),
            .I(N__10194));
    Odrv12 I__2419 (
            .O(N__10194),
            .I(TCIn_1_i));
    InMux I__2418 (
            .O(N__10191),
            .I(N__10188));
    LocalMux I__2417 (
            .O(N__10188),
            .I(N__10184));
    InMux I__2416 (
            .O(N__10187),
            .I(N__10181));
    Span4Mux_v I__2415 (
            .O(N__10184),
            .I(N__10171));
    LocalMux I__2414 (
            .O(N__10181),
            .I(N__10171));
    CascadeMux I__2413 (
            .O(N__10180),
            .I(N__10164));
    CascadeMux I__2412 (
            .O(N__10179),
            .I(N__10161));
    InMux I__2411 (
            .O(N__10178),
            .I(N__10157));
    CascadeMux I__2410 (
            .O(N__10177),
            .I(N__10154));
    InMux I__2409 (
            .O(N__10176),
            .I(N__10150));
    Span4Mux_v I__2408 (
            .O(N__10171),
            .I(N__10141));
    InMux I__2407 (
            .O(N__10170),
            .I(N__10138));
    InMux I__2406 (
            .O(N__10169),
            .I(N__10135));
    InMux I__2405 (
            .O(N__10168),
            .I(N__10124));
    InMux I__2404 (
            .O(N__10167),
            .I(N__10124));
    InMux I__2403 (
            .O(N__10164),
            .I(N__10124));
    InMux I__2402 (
            .O(N__10161),
            .I(N__10124));
    InMux I__2401 (
            .O(N__10160),
            .I(N__10124));
    LocalMux I__2400 (
            .O(N__10157),
            .I(N__10121));
    InMux I__2399 (
            .O(N__10154),
            .I(N__10116));
    InMux I__2398 (
            .O(N__10153),
            .I(N__10116));
    LocalMux I__2397 (
            .O(N__10150),
            .I(N__10113));
    InMux I__2396 (
            .O(N__10149),
            .I(N__10110));
    InMux I__2395 (
            .O(N__10148),
            .I(N__10107));
    InMux I__2394 (
            .O(N__10147),
            .I(N__10104));
    CascadeMux I__2393 (
            .O(N__10146),
            .I(N__10101));
    CascadeMux I__2392 (
            .O(N__10145),
            .I(N__10098));
    CascadeMux I__2391 (
            .O(N__10144),
            .I(N__10095));
    Span4Mux_h I__2390 (
            .O(N__10141),
            .I(N__10081));
    LocalMux I__2389 (
            .O(N__10138),
            .I(N__10081));
    LocalMux I__2388 (
            .O(N__10135),
            .I(N__10081));
    LocalMux I__2387 (
            .O(N__10124),
            .I(N__10081));
    Span4Mux_h I__2386 (
            .O(N__10121),
            .I(N__10081));
    LocalMux I__2385 (
            .O(N__10116),
            .I(N__10081));
    Span4Mux_v I__2384 (
            .O(N__10113),
            .I(N__10073));
    LocalMux I__2383 (
            .O(N__10110),
            .I(N__10073));
    LocalMux I__2382 (
            .O(N__10107),
            .I(N__10073));
    LocalMux I__2381 (
            .O(N__10104),
            .I(N__10070));
    InMux I__2380 (
            .O(N__10101),
            .I(N__10063));
    InMux I__2379 (
            .O(N__10098),
            .I(N__10063));
    InMux I__2378 (
            .O(N__10095),
            .I(N__10063));
    InMux I__2377 (
            .O(N__10094),
            .I(N__10057));
    Span4Mux_v I__2376 (
            .O(N__10081),
            .I(N__10054));
    InMux I__2375 (
            .O(N__10080),
            .I(N__10051));
    Span4Mux_v I__2374 (
            .O(N__10073),
            .I(N__10048));
    Span4Mux_h I__2373 (
            .O(N__10070),
            .I(N__10043));
    LocalMux I__2372 (
            .O(N__10063),
            .I(N__10043));
    InMux I__2371 (
            .O(N__10062),
            .I(N__10038));
    InMux I__2370 (
            .O(N__10061),
            .I(N__10038));
    InMux I__2369 (
            .O(N__10060),
            .I(N__10035));
    LocalMux I__2368 (
            .O(N__10057),
            .I(N__10028));
    Span4Mux_h I__2367 (
            .O(N__10054),
            .I(N__10028));
    LocalMux I__2366 (
            .O(N__10051),
            .I(N__10028));
    Span4Mux_h I__2365 (
            .O(N__10048),
            .I(N__10024));
    Span4Mux_h I__2364 (
            .O(N__10043),
            .I(N__10017));
    LocalMux I__2363 (
            .O(N__10038),
            .I(N__10017));
    LocalMux I__2362 (
            .O(N__10035),
            .I(N__10017));
    Span4Mux_v I__2361 (
            .O(N__10028),
            .I(N__10014));
    InMux I__2360 (
            .O(N__10027),
            .I(N__10011));
    Span4Mux_h I__2359 (
            .O(N__10024),
            .I(N__10006));
    Span4Mux_v I__2358 (
            .O(N__10017),
            .I(N__10006));
    Sp12to4 I__2357 (
            .O(N__10014),
            .I(N__10002));
    LocalMux I__2356 (
            .O(N__10011),
            .I(N__9999));
    Span4Mux_v I__2355 (
            .O(N__10006),
            .I(N__9996));
    InMux I__2354 (
            .O(N__10005),
            .I(N__9993));
    Span12Mux_h I__2353 (
            .O(N__10002),
            .I(N__9990));
    Span12Mux_v I__2352 (
            .O(N__9999),
            .I(N__9983));
    Sp12to4 I__2351 (
            .O(N__9996),
            .I(N__9983));
    LocalMux I__2350 (
            .O(N__9993),
            .I(N__9983));
    Span12Mux_v I__2349 (
            .O(N__9990),
            .I(N__9978));
    Span12Mux_h I__2348 (
            .O(N__9983),
            .I(N__9978));
    Odrv12 I__2347 (
            .O(N__9978),
            .I(RESETn_c));
    InMux I__2346 (
            .O(N__9975),
            .I(N__9971));
    InMux I__2345 (
            .O(N__9974),
            .I(N__9968));
    LocalMux I__2344 (
            .O(N__9971),
            .I(N__9965));
    LocalMux I__2343 (
            .O(N__9968),
            .I(N__9962));
    Span12Mux_s11_v I__2342 (
            .O(N__9965),
            .I(N__9958));
    Span4Mux_h I__2341 (
            .O(N__9962),
            .I(N__9955));
    InMux I__2340 (
            .O(N__9961),
            .I(N__9952));
    Odrv12 I__2339 (
            .O(N__9958),
            .I(\U409_CIA.VMAZ0 ));
    Odrv4 I__2338 (
            .O(N__9955),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__2337 (
            .O(N__9952),
            .I(\U409_CIA.VMAZ0 ));
    CascadeMux I__2336 (
            .O(N__9945),
            .I(\U409_CIA.CIA_CLK_COUNT11_3_cascade_ ));
    InMux I__2335 (
            .O(N__9942),
            .I(N__9939));
    LocalMux I__2334 (
            .O(N__9939),
            .I(\U409_CIA.CIA_CLK_COUNT11_2_0 ));
    InMux I__2333 (
            .O(N__9936),
            .I(N__9933));
    LocalMux I__2332 (
            .O(N__9933),
            .I(\U409_CIA.CIA_CLK_COUNT11_3 ));
    CascadeMux I__2331 (
            .O(N__9930),
            .I(\U409_CIA.CIA_CLK_COUNT11_2_0_cascade_ ));
    CascadeMux I__2330 (
            .O(N__9927),
            .I(\U409_CIA.CLK_CIA6_4_cascade_ ));
    CascadeMux I__2329 (
            .O(N__9924),
            .I(\U409_CIA.VMA_RNOZ0Z_0_cascade_ ));
    InMux I__2328 (
            .O(N__9921),
            .I(N__9911));
    InMux I__2327 (
            .O(N__9920),
            .I(N__9911));
    InMux I__2326 (
            .O(N__9919),
            .I(N__9904));
    InMux I__2325 (
            .O(N__9918),
            .I(N__9904));
    InMux I__2324 (
            .O(N__9917),
            .I(N__9904));
    InMux I__2323 (
            .O(N__9916),
            .I(N__9901));
    LocalMux I__2322 (
            .O(N__9911),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__2321 (
            .O(N__9904),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__2320 (
            .O(N__9901),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    InMux I__2319 (
            .O(N__9894),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ));
    CascadeMux I__2318 (
            .O(N__9891),
            .I(\U409_TICK.TICK503_9_cascade_ ));
    InMux I__2317 (
            .O(N__9888),
            .I(N__9885));
    LocalMux I__2316 (
            .O(N__9885),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ));
    CascadeMux I__2315 (
            .O(N__9882),
            .I(N__9879));
    InMux I__2314 (
            .O(N__9879),
            .I(N__9875));
    InMux I__2313 (
            .O(N__9878),
            .I(N__9872));
    LocalMux I__2312 (
            .O(N__9875),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    LocalMux I__2311 (
            .O(N__9872),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    InMux I__2310 (
            .O(N__9867),
            .I(N__9863));
    InMux I__2309 (
            .O(N__9866),
            .I(N__9860));
    LocalMux I__2308 (
            .O(N__9863),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    LocalMux I__2307 (
            .O(N__9860),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    CascadeMux I__2306 (
            .O(N__9855),
            .I(N__9852));
    InMux I__2305 (
            .O(N__9852),
            .I(N__9848));
    InMux I__2304 (
            .O(N__9851),
            .I(N__9845));
    LocalMux I__2303 (
            .O(N__9848),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    LocalMux I__2302 (
            .O(N__9845),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    InMux I__2301 (
            .O(N__9840),
            .I(N__9837));
    LocalMux I__2300 (
            .O(N__9837),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ));
    InMux I__2299 (
            .O(N__9834),
            .I(N__9830));
    InMux I__2298 (
            .O(N__9833),
            .I(N__9827));
    LocalMux I__2297 (
            .O(N__9830),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    LocalMux I__2296 (
            .O(N__9827),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    InMux I__2295 (
            .O(N__9822),
            .I(N__9819));
    LocalMux I__2294 (
            .O(N__9819),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ));
    InMux I__2293 (
            .O(N__9816),
            .I(N__9812));
    InMux I__2292 (
            .O(N__9815),
            .I(N__9809));
    LocalMux I__2291 (
            .O(N__9812),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    LocalMux I__2290 (
            .O(N__9809),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    InMux I__2289 (
            .O(N__9804),
            .I(N__9801));
    LocalMux I__2288 (
            .O(N__9801),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ));
    InMux I__2287 (
            .O(N__9798),
            .I(N__9794));
    InMux I__2286 (
            .O(N__9797),
            .I(N__9791));
    LocalMux I__2285 (
            .O(N__9794),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    LocalMux I__2284 (
            .O(N__9791),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    InMux I__2283 (
            .O(N__9786),
            .I(N__9773));
    InMux I__2282 (
            .O(N__9785),
            .I(N__9773));
    InMux I__2281 (
            .O(N__9784),
            .I(N__9768));
    InMux I__2280 (
            .O(N__9783),
            .I(N__9768));
    InMux I__2279 (
            .O(N__9782),
            .I(N__9759));
    InMux I__2278 (
            .O(N__9781),
            .I(N__9759));
    InMux I__2277 (
            .O(N__9780),
            .I(N__9759));
    InMux I__2276 (
            .O(N__9779),
            .I(N__9759));
    InMux I__2275 (
            .O(N__9778),
            .I(N__9756));
    LocalMux I__2274 (
            .O(N__9773),
            .I(N__9753));
    LocalMux I__2273 (
            .O(N__9768),
            .I(N__9750));
    LocalMux I__2272 (
            .O(N__9759),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__2271 (
            .O(N__9756),
            .I(\U409_TICK.TICK503_10 ));
    Odrv4 I__2270 (
            .O(N__9753),
            .I(\U409_TICK.TICK503_10 ));
    Odrv4 I__2269 (
            .O(N__9750),
            .I(\U409_TICK.TICK503_10 ));
    CascadeMux I__2268 (
            .O(N__9741),
            .I(N__9737));
    InMux I__2267 (
            .O(N__9740),
            .I(N__9727));
    InMux I__2266 (
            .O(N__9737),
            .I(N__9724));
    InMux I__2265 (
            .O(N__9736),
            .I(N__9719));
    InMux I__2264 (
            .O(N__9735),
            .I(N__9719));
    InMux I__2263 (
            .O(N__9734),
            .I(N__9716));
    InMux I__2262 (
            .O(N__9733),
            .I(N__9707));
    InMux I__2261 (
            .O(N__9732),
            .I(N__9707));
    InMux I__2260 (
            .O(N__9731),
            .I(N__9707));
    InMux I__2259 (
            .O(N__9730),
            .I(N__9707));
    LocalMux I__2258 (
            .O(N__9727),
            .I(N__9704));
    LocalMux I__2257 (
            .O(N__9724),
            .I(N__9699));
    LocalMux I__2256 (
            .O(N__9719),
            .I(N__9699));
    LocalMux I__2255 (
            .O(N__9716),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__2254 (
            .O(N__9707),
            .I(\U409_TICK.TICK503_14 ));
    Odrv4 I__2253 (
            .O(N__9704),
            .I(\U409_TICK.TICK503_14 ));
    Odrv4 I__2252 (
            .O(N__9699),
            .I(\U409_TICK.TICK503_14 ));
    CascadeMux I__2251 (
            .O(N__9690),
            .I(N__9687));
    InMux I__2250 (
            .O(N__9687),
            .I(N__9677));
    InMux I__2249 (
            .O(N__9686),
            .I(N__9674));
    InMux I__2248 (
            .O(N__9685),
            .I(N__9669));
    InMux I__2247 (
            .O(N__9684),
            .I(N__9669));
    CascadeMux I__2246 (
            .O(N__9683),
            .I(N__9666));
    CascadeMux I__2245 (
            .O(N__9682),
            .I(N__9663));
    CascadeMux I__2244 (
            .O(N__9681),
            .I(N__9660));
    CascadeMux I__2243 (
            .O(N__9680),
            .I(N__9657));
    LocalMux I__2242 (
            .O(N__9677),
            .I(N__9652));
    LocalMux I__2241 (
            .O(N__9674),
            .I(N__9652));
    LocalMux I__2240 (
            .O(N__9669),
            .I(N__9649));
    InMux I__2239 (
            .O(N__9666),
            .I(N__9644));
    InMux I__2238 (
            .O(N__9663),
            .I(N__9644));
    InMux I__2237 (
            .O(N__9660),
            .I(N__9639));
    InMux I__2236 (
            .O(N__9657),
            .I(N__9639));
    Span4Mux_h I__2235 (
            .O(N__9652),
            .I(N__9634));
    Span4Mux_v I__2234 (
            .O(N__9649),
            .I(N__9634));
    LocalMux I__2233 (
            .O(N__9644),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__2232 (
            .O(N__9639),
            .I(\U409_TICK.TICK503_9 ));
    Odrv4 I__2231 (
            .O(N__9634),
            .I(\U409_TICK.TICK503_9 ));
    InMux I__2230 (
            .O(N__9627),
            .I(N__9624));
    LocalMux I__2229 (
            .O(N__9624),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ));
    InMux I__2228 (
            .O(N__9621),
            .I(N__9617));
    InMux I__2227 (
            .O(N__9620),
            .I(N__9614));
    LocalMux I__2226 (
            .O(N__9617),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    LocalMux I__2225 (
            .O(N__9614),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    ClkMux I__2224 (
            .O(N__9609),
            .I(N__9573));
    ClkMux I__2223 (
            .O(N__9608),
            .I(N__9573));
    ClkMux I__2222 (
            .O(N__9607),
            .I(N__9573));
    ClkMux I__2221 (
            .O(N__9606),
            .I(N__9573));
    ClkMux I__2220 (
            .O(N__9605),
            .I(N__9573));
    ClkMux I__2219 (
            .O(N__9604),
            .I(N__9573));
    ClkMux I__2218 (
            .O(N__9603),
            .I(N__9573));
    ClkMux I__2217 (
            .O(N__9602),
            .I(N__9573));
    ClkMux I__2216 (
            .O(N__9601),
            .I(N__9573));
    ClkMux I__2215 (
            .O(N__9600),
            .I(N__9573));
    ClkMux I__2214 (
            .O(N__9599),
            .I(N__9573));
    ClkMux I__2213 (
            .O(N__9598),
            .I(N__9573));
    GlobalMux I__2212 (
            .O(N__9573),
            .I(N__9570));
    gio2CtrlBuf I__2211 (
            .O(N__9570),
            .I(CLK6_c_g));
    InMux I__2210 (
            .O(N__9567),
            .I(N__9564));
    LocalMux I__2209 (
            .O(N__9564),
            .I(\U409_CIA.CLK_CIA6_3 ));
    InMux I__2208 (
            .O(N__9561),
            .I(N__9557));
    InMux I__2207 (
            .O(N__9560),
            .I(N__9554));
    LocalMux I__2206 (
            .O(N__9557),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    LocalMux I__2205 (
            .O(N__9554),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    InMux I__2204 (
            .O(N__9549),
            .I(N__9546));
    LocalMux I__2203 (
            .O(N__9546),
            .I(N__9543));
    Span4Mux_h I__2202 (
            .O(N__9543),
            .I(N__9540));
    Odrv4 I__2201 (
            .O(N__9540),
            .I(\U409_TICK.TICK503_11 ));
    CascadeMux I__2200 (
            .O(N__9537),
            .I(\U409_TICK.TICK503_8_cascade_ ));
    InMux I__2199 (
            .O(N__9534),
            .I(N__9530));
    InMux I__2198 (
            .O(N__9533),
            .I(N__9527));
    LocalMux I__2197 (
            .O(N__9530),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    LocalMux I__2196 (
            .O(N__9527),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    InMux I__2195 (
            .O(N__9522),
            .I(N__9519));
    LocalMux I__2194 (
            .O(N__9519),
            .I(N__9515));
    InMux I__2193 (
            .O(N__9518),
            .I(N__9512));
    Odrv4 I__2192 (
            .O(N__9515),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    LocalMux I__2191 (
            .O(N__9512),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    InMux I__2190 (
            .O(N__9507),
            .I(N__9503));
    InMux I__2189 (
            .O(N__9506),
            .I(N__9500));
    LocalMux I__2188 (
            .O(N__9503),
            .I(N__9497));
    LocalMux I__2187 (
            .O(N__9500),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    Odrv4 I__2186 (
            .O(N__9497),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    CascadeMux I__2185 (
            .O(N__9492),
            .I(\U409_TICK.TICK603_9_cascade_ ));
    InMux I__2184 (
            .O(N__9489),
            .I(N__9486));
    LocalMux I__2183 (
            .O(N__9486),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ));
    InMux I__2182 (
            .O(N__9483),
            .I(N__9479));
    InMux I__2181 (
            .O(N__9482),
            .I(N__9476));
    LocalMux I__2180 (
            .O(N__9479),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    LocalMux I__2179 (
            .O(N__9476),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    CascadeMux I__2178 (
            .O(N__9471),
            .I(N__9468));
    InMux I__2177 (
            .O(N__9468),
            .I(N__9465));
    LocalMux I__2176 (
            .O(N__9465),
            .I(N__9462));
    Odrv4 I__2175 (
            .O(N__9462),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ));
    IoInMux I__2174 (
            .O(N__9459),
            .I(N__9456));
    LocalMux I__2173 (
            .O(N__9456),
            .I(N__9453));
    Span4Mux_s2_v I__2172 (
            .O(N__9453),
            .I(N__9450));
    Span4Mux_v I__2171 (
            .O(N__9450),
            .I(N__9447));
    Sp12to4 I__2170 (
            .O(N__9447),
            .I(N__9444));
    Span12Mux_h I__2169 (
            .O(N__9444),
            .I(N__9440));
    InMux I__2168 (
            .O(N__9443),
            .I(N__9437));
    Odrv12 I__2167 (
            .O(N__9440),
            .I(TICK50_c));
    LocalMux I__2166 (
            .O(N__9437),
            .I(TICK50_c));
    CascadeMux I__2165 (
            .O(N__9432),
            .I(N__9429));
    InMux I__2164 (
            .O(N__9429),
            .I(N__9426));
    LocalMux I__2163 (
            .O(N__9426),
            .I(N__9423));
    Span4Mux_h I__2162 (
            .O(N__9423),
            .I(N__9420));
    Odrv4 I__2161 (
            .O(N__9420),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ));
    CascadeMux I__2160 (
            .O(N__9417),
            .I(N__9413));
    InMux I__2159 (
            .O(N__9416),
            .I(N__9410));
    InMux I__2158 (
            .O(N__9413),
            .I(N__9407));
    LocalMux I__2157 (
            .O(N__9410),
            .I(N__9404));
    LocalMux I__2156 (
            .O(N__9407),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    Odrv4 I__2155 (
            .O(N__9404),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    InMux I__2154 (
            .O(N__9399),
            .I(N__9390));
    InMux I__2153 (
            .O(N__9398),
            .I(N__9383));
    InMux I__2152 (
            .O(N__9397),
            .I(N__9383));
    InMux I__2151 (
            .O(N__9396),
            .I(N__9383));
    InMux I__2150 (
            .O(N__9395),
            .I(N__9376));
    InMux I__2149 (
            .O(N__9394),
            .I(N__9376));
    InMux I__2148 (
            .O(N__9393),
            .I(N__9376));
    LocalMux I__2147 (
            .O(N__9390),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__2146 (
            .O(N__9383),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__2145 (
            .O(N__9376),
            .I(\U409_TICK.TICK603_14 ));
    InMux I__2144 (
            .O(N__9369),
            .I(N__9359));
    InMux I__2143 (
            .O(N__9368),
            .I(N__9352));
    InMux I__2142 (
            .O(N__9367),
            .I(N__9352));
    InMux I__2141 (
            .O(N__9366),
            .I(N__9352));
    InMux I__2140 (
            .O(N__9365),
            .I(N__9343));
    InMux I__2139 (
            .O(N__9364),
            .I(N__9343));
    InMux I__2138 (
            .O(N__9363),
            .I(N__9343));
    InMux I__2137 (
            .O(N__9362),
            .I(N__9343));
    LocalMux I__2136 (
            .O(N__9359),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__2135 (
            .O(N__9352),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__2134 (
            .O(N__9343),
            .I(\U409_TICK.TICK603_10 ));
    CascadeMux I__2133 (
            .O(N__9336),
            .I(N__9330));
    CascadeMux I__2132 (
            .O(N__9335),
            .I(N__9326));
    CascadeMux I__2131 (
            .O(N__9334),
            .I(N__9322));
    CascadeMux I__2130 (
            .O(N__9333),
            .I(N__9319));
    InMux I__2129 (
            .O(N__9330),
            .I(N__9315));
    InMux I__2128 (
            .O(N__9329),
            .I(N__9310));
    InMux I__2127 (
            .O(N__9326),
            .I(N__9310));
    InMux I__2126 (
            .O(N__9325),
            .I(N__9301));
    InMux I__2125 (
            .O(N__9322),
            .I(N__9301));
    InMux I__2124 (
            .O(N__9319),
            .I(N__9301));
    InMux I__2123 (
            .O(N__9318),
            .I(N__9301));
    LocalMux I__2122 (
            .O(N__9315),
            .I(N__9298));
    LocalMux I__2121 (
            .O(N__9310),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__2120 (
            .O(N__9301),
            .I(\U409_TICK.TICK603_9 ));
    Odrv4 I__2119 (
            .O(N__9298),
            .I(\U409_TICK.TICK603_9 ));
    IoInMux I__2118 (
            .O(N__9291),
            .I(N__9288));
    LocalMux I__2117 (
            .O(N__9288),
            .I(N__9285));
    Span4Mux_s3_v I__2116 (
            .O(N__9285),
            .I(N__9282));
    Span4Mux_v I__2115 (
            .O(N__9282),
            .I(N__9279));
    Span4Mux_v I__2114 (
            .O(N__9279),
            .I(N__9276));
    Span4Mux_h I__2113 (
            .O(N__9276),
            .I(N__9272));
    InMux I__2112 (
            .O(N__9275),
            .I(N__9269));
    Odrv4 I__2111 (
            .O(N__9272),
            .I(TICK60_c));
    LocalMux I__2110 (
            .O(N__9269),
            .I(TICK60_c));
    InMux I__2109 (
            .O(N__9264),
            .I(N__9260));
    InMux I__2108 (
            .O(N__9263),
            .I(N__9257));
    LocalMux I__2107 (
            .O(N__9260),
            .I(N__9254));
    LocalMux I__2106 (
            .O(N__9257),
            .I(N__9251));
    Odrv4 I__2105 (
            .O(N__9254),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    Odrv4 I__2104 (
            .O(N__9251),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    InMux I__2103 (
            .O(N__9246),
            .I(\U409_TICK.un2_COUNTER50_1_cry_10 ));
    InMux I__2102 (
            .O(N__9243),
            .I(\U409_TICK.un2_COUNTER50_1_cry_11 ));
    InMux I__2101 (
            .O(N__9240),
            .I(\U409_TICK.un2_COUNTER50_1_cry_12 ));
    InMux I__2100 (
            .O(N__9237),
            .I(\U409_TICK.un2_COUNTER50_1_cry_13 ));
    InMux I__2099 (
            .O(N__9234),
            .I(\U409_TICK.un2_COUNTER50_1_cry_14 ));
    InMux I__2098 (
            .O(N__9231),
            .I(\U409_TICK.un2_COUNTER50_1_cry_15 ));
    InMux I__2097 (
            .O(N__9228),
            .I(N__9224));
    InMux I__2096 (
            .O(N__9227),
            .I(N__9221));
    LocalMux I__2095 (
            .O(N__9224),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    LocalMux I__2094 (
            .O(N__9221),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    CascadeMux I__2093 (
            .O(N__9216),
            .I(\U409_CIA.CLK_CIA_r_1_0_cascade_ ));
    IoInMux I__2092 (
            .O(N__9213),
            .I(N__9210));
    LocalMux I__2091 (
            .O(N__9210),
            .I(N__9207));
    IoSpan4Mux I__2090 (
            .O(N__9207),
            .I(N__9204));
    Span4Mux_s3_v I__2089 (
            .O(N__9204),
            .I(N__9201));
    Sp12to4 I__2088 (
            .O(N__9201),
            .I(N__9196));
    InMux I__2087 (
            .O(N__9200),
            .I(N__9193));
    CascadeMux I__2086 (
            .O(N__9199),
            .I(N__9189));
    Span12Mux_s10_v I__2085 (
            .O(N__9196),
            .I(N__9186));
    LocalMux I__2084 (
            .O(N__9193),
            .I(N__9183));
    InMux I__2083 (
            .O(N__9192),
            .I(N__9180));
    InMux I__2082 (
            .O(N__9189),
            .I(N__9177));
    Odrv12 I__2081 (
            .O(N__9186),
            .I(CLK_CIA_c));
    Odrv4 I__2080 (
            .O(N__9183),
            .I(CLK_CIA_c));
    LocalMux I__2079 (
            .O(N__9180),
            .I(CLK_CIA_c));
    LocalMux I__2078 (
            .O(N__9177),
            .I(CLK_CIA_c));
    InMux I__2077 (
            .O(N__9168),
            .I(N__9165));
    LocalMux I__2076 (
            .O(N__9165),
            .I(N__9161));
    CascadeMux I__2075 (
            .O(N__9164),
            .I(N__9158));
    Span4Mux_h I__2074 (
            .O(N__9161),
            .I(N__9155));
    InMux I__2073 (
            .O(N__9158),
            .I(N__9152));
    Odrv4 I__2072 (
            .O(N__9155),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    LocalMux I__2071 (
            .O(N__9152),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    CascadeMux I__2070 (
            .O(N__9147),
            .I(N__9144));
    InMux I__2069 (
            .O(N__9144),
            .I(N__9141));
    LocalMux I__2068 (
            .O(N__9141),
            .I(N__9137));
    InMux I__2067 (
            .O(N__9140),
            .I(N__9134));
    Odrv12 I__2066 (
            .O(N__9137),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    LocalMux I__2065 (
            .O(N__9134),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    InMux I__2064 (
            .O(N__9129),
            .I(N__9125));
    CascadeMux I__2063 (
            .O(N__9128),
            .I(N__9121));
    LocalMux I__2062 (
            .O(N__9125),
            .I(N__9117));
    CascadeMux I__2061 (
            .O(N__9124),
            .I(N__9114));
    InMux I__2060 (
            .O(N__9121),
            .I(N__9111));
    InMux I__2059 (
            .O(N__9120),
            .I(N__9108));
    Span4Mux_h I__2058 (
            .O(N__9117),
            .I(N__9105));
    InMux I__2057 (
            .O(N__9114),
            .I(N__9102));
    LocalMux I__2056 (
            .O(N__9111),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__2055 (
            .O(N__9108),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    Odrv4 I__2054 (
            .O(N__9105),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__2053 (
            .O(N__9102),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    CascadeMux I__2052 (
            .O(N__9093),
            .I(N__9090));
    InMux I__2051 (
            .O(N__9090),
            .I(N__9086));
    InMux I__2050 (
            .O(N__9089),
            .I(N__9083));
    LocalMux I__2049 (
            .O(N__9086),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    LocalMux I__2048 (
            .O(N__9083),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    InMux I__2047 (
            .O(N__9078),
            .I(\U409_TICK.un2_COUNTER50_1_cry_1 ));
    InMux I__2046 (
            .O(N__9075),
            .I(\U409_TICK.un2_COUNTER50_1_cry_2 ));
    InMux I__2045 (
            .O(N__9072),
            .I(\U409_TICK.un2_COUNTER50_1_cry_3 ));
    InMux I__2044 (
            .O(N__9069),
            .I(N__9066));
    LocalMux I__2043 (
            .O(N__9066),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ));
    InMux I__2042 (
            .O(N__9063),
            .I(\U409_TICK.un2_COUNTER50_1_cry_4 ));
    InMux I__2041 (
            .O(N__9060),
            .I(\U409_TICK.un2_COUNTER50_1_cry_5 ));
    InMux I__2040 (
            .O(N__9057),
            .I(\U409_TICK.un2_COUNTER50_1_cry_6 ));
    InMux I__2039 (
            .O(N__9054),
            .I(N__9050));
    InMux I__2038 (
            .O(N__9053),
            .I(N__9047));
    LocalMux I__2037 (
            .O(N__9050),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    LocalMux I__2036 (
            .O(N__9047),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    InMux I__2035 (
            .O(N__9042),
            .I(\U409_TICK.un2_COUNTER50_1_cry_7 ));
    InMux I__2034 (
            .O(N__9039),
            .I(bfn_14_6_0_));
    InMux I__2033 (
            .O(N__9036),
            .I(\U409_TICK.un2_COUNTER50_1_cry_9 ));
    InMux I__2032 (
            .O(N__9033),
            .I(N__9030));
    LocalMux I__2031 (
            .O(N__9030),
            .I(N__9020));
    SRMux I__2030 (
            .O(N__9029),
            .I(N__8991));
    SRMux I__2029 (
            .O(N__9028),
            .I(N__8991));
    SRMux I__2028 (
            .O(N__9027),
            .I(N__8991));
    SRMux I__2027 (
            .O(N__9026),
            .I(N__8991));
    SRMux I__2026 (
            .O(N__9025),
            .I(N__8991));
    SRMux I__2025 (
            .O(N__9024),
            .I(N__8991));
    SRMux I__2024 (
            .O(N__9023),
            .I(N__8991));
    Glb2LocalMux I__2023 (
            .O(N__9020),
            .I(N__8991));
    SRMux I__2022 (
            .O(N__9019),
            .I(N__8991));
    SRMux I__2021 (
            .O(N__9018),
            .I(N__8991));
    SRMux I__2020 (
            .O(N__9017),
            .I(N__8991));
    SRMux I__2019 (
            .O(N__9016),
            .I(N__8991));
    GlobalMux I__2018 (
            .O(N__8991),
            .I(N__8988));
    gio2CtrlBuf I__2017 (
            .O(N__8988),
            .I(RESETn_c_i_g));
    CascadeMux I__2016 (
            .O(N__8985),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1_cascade_ ));
    InMux I__2015 (
            .O(N__8982),
            .I(N__8978));
    InMux I__2014 (
            .O(N__8981),
            .I(N__8975));
    LocalMux I__2013 (
            .O(N__8978),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ));
    LocalMux I__2012 (
            .O(N__8975),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ));
    CascadeMux I__2011 (
            .O(N__8970),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out_cascade_ ));
    InMux I__2010 (
            .O(N__8967),
            .I(N__8959));
    InMux I__2009 (
            .O(N__8966),
            .I(N__8959));
    InMux I__2008 (
            .O(N__8965),
            .I(N__8954));
    InMux I__2007 (
            .O(N__8964),
            .I(N__8954));
    LocalMux I__2006 (
            .O(N__8959),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__2005 (
            .O(N__8954),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    InMux I__2004 (
            .O(N__8949),
            .I(N__8938));
    InMux I__2003 (
            .O(N__8948),
            .I(N__8938));
    InMux I__2002 (
            .O(N__8947),
            .I(N__8938));
    InMux I__2001 (
            .O(N__8946),
            .I(N__8933));
    InMux I__2000 (
            .O(N__8945),
            .I(N__8933));
    LocalMux I__1999 (
            .O(N__8938),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__1998 (
            .O(N__8933),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    InMux I__1997 (
            .O(N__8928),
            .I(N__8919));
    InMux I__1996 (
            .O(N__8927),
            .I(N__8919));
    InMux I__1995 (
            .O(N__8926),
            .I(N__8914));
    InMux I__1994 (
            .O(N__8925),
            .I(N__8914));
    InMux I__1993 (
            .O(N__8924),
            .I(N__8911));
    LocalMux I__1992 (
            .O(N__8919),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1991 (
            .O(N__8914),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1990 (
            .O(N__8911),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    CascadeMux I__1989 (
            .O(N__8904),
            .I(N__8900));
    CascadeMux I__1988 (
            .O(N__8903),
            .I(N__8895));
    InMux I__1987 (
            .O(N__8900),
            .I(N__8885));
    InMux I__1986 (
            .O(N__8899),
            .I(N__8885));
    InMux I__1985 (
            .O(N__8898),
            .I(N__8885));
    InMux I__1984 (
            .O(N__8895),
            .I(N__8880));
    InMux I__1983 (
            .O(N__8894),
            .I(N__8880));
    InMux I__1982 (
            .O(N__8893),
            .I(N__8875));
    InMux I__1981 (
            .O(N__8892),
            .I(N__8875));
    LocalMux I__1980 (
            .O(N__8885),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1979 (
            .O(N__8880),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1978 (
            .O(N__8875),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    InMux I__1977 (
            .O(N__8868),
            .I(N__8862));
    InMux I__1976 (
            .O(N__8867),
            .I(N__8857));
    InMux I__1975 (
            .O(N__8866),
            .I(N__8857));
    InMux I__1974 (
            .O(N__8865),
            .I(N__8854));
    LocalMux I__1973 (
            .O(N__8862),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1972 (
            .O(N__8857),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1971 (
            .O(N__8854),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    CascadeMux I__1970 (
            .O(N__8847),
            .I(N__8843));
    InMux I__1969 (
            .O(N__8846),
            .I(N__8838));
    InMux I__1968 (
            .O(N__8843),
            .I(N__8838));
    LocalMux I__1967 (
            .O(N__8838),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ));
    InMux I__1966 (
            .O(N__8835),
            .I(N__8826));
    InMux I__1965 (
            .O(N__8834),
            .I(N__8826));
    InMux I__1964 (
            .O(N__8833),
            .I(N__8823));
    InMux I__1963 (
            .O(N__8832),
            .I(N__8818));
    InMux I__1962 (
            .O(N__8831),
            .I(N__8818));
    LocalMux I__1961 (
            .O(N__8826),
            .I(N__8815));
    LocalMux I__1960 (
            .O(N__8823),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__1959 (
            .O(N__8818),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    Odrv4 I__1958 (
            .O(N__8815),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    CascadeMux I__1957 (
            .O(N__8808),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ));
    CascadeMux I__1956 (
            .O(N__8805),
            .I(N__8799));
    InMux I__1955 (
            .O(N__8804),
            .I(N__8788));
    InMux I__1954 (
            .O(N__8803),
            .I(N__8788));
    InMux I__1953 (
            .O(N__8802),
            .I(N__8788));
    InMux I__1952 (
            .O(N__8799),
            .I(N__8788));
    InMux I__1951 (
            .O(N__8798),
            .I(N__8783));
    InMux I__1950 (
            .O(N__8797),
            .I(N__8783));
    LocalMux I__1949 (
            .O(N__8788),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1948 (
            .O(N__8783),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    SRMux I__1947 (
            .O(N__8778),
            .I(N__8774));
    SRMux I__1946 (
            .O(N__8777),
            .I(N__8770));
    LocalMux I__1945 (
            .O(N__8774),
            .I(N__8767));
    SRMux I__1944 (
            .O(N__8773),
            .I(N__8763));
    LocalMux I__1943 (
            .O(N__8770),
            .I(N__8760));
    Span4Mux_h I__1942 (
            .O(N__8767),
            .I(N__8757));
    SRMux I__1941 (
            .O(N__8766),
            .I(N__8754));
    LocalMux I__1940 (
            .O(N__8763),
            .I(N__8751));
    Span4Mux_v I__1939 (
            .O(N__8760),
            .I(N__8748));
    Span4Mux_v I__1938 (
            .O(N__8757),
            .I(N__8743));
    LocalMux I__1937 (
            .O(N__8754),
            .I(N__8743));
    Span4Mux_v I__1936 (
            .O(N__8751),
            .I(N__8740));
    Sp12to4 I__1935 (
            .O(N__8748),
            .I(N__8735));
    Sp12to4 I__1934 (
            .O(N__8743),
            .I(N__8735));
    Odrv4 I__1933 (
            .O(N__8740),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    Odrv12 I__1932 (
            .O(N__8735),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    InMux I__1931 (
            .O(N__8730),
            .I(N__8725));
    InMux I__1930 (
            .O(N__8729),
            .I(N__8722));
    InMux I__1929 (
            .O(N__8728),
            .I(N__8719));
    LocalMux I__1928 (
            .O(N__8725),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__1927 (
            .O(N__8722),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__1926 (
            .O(N__8719),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    InMux I__1925 (
            .O(N__8712),
            .I(N__8709));
    LocalMux I__1924 (
            .O(N__8709),
            .I(N__8705));
    InMux I__1923 (
            .O(N__8708),
            .I(N__8702));
    Odrv4 I__1922 (
            .O(N__8705),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    LocalMux I__1921 (
            .O(N__8702),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    InMux I__1920 (
            .O(N__8697),
            .I(N__8693));
    InMux I__1919 (
            .O(N__8696),
            .I(N__8690));
    LocalMux I__1918 (
            .O(N__8693),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    LocalMux I__1917 (
            .O(N__8690),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    CascadeMux I__1916 (
            .O(N__8685),
            .I(N__8682));
    InMux I__1915 (
            .O(N__8682),
            .I(N__8678));
    InMux I__1914 (
            .O(N__8681),
            .I(N__8675));
    LocalMux I__1913 (
            .O(N__8678),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    LocalMux I__1912 (
            .O(N__8675),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    InMux I__1911 (
            .O(N__8670),
            .I(N__8666));
    InMux I__1910 (
            .O(N__8669),
            .I(N__8663));
    LocalMux I__1909 (
            .O(N__8666),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    LocalMux I__1908 (
            .O(N__8663),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    InMux I__1907 (
            .O(N__8658),
            .I(N__8655));
    LocalMux I__1906 (
            .O(N__8655),
            .I(N__8651));
    InMux I__1905 (
            .O(N__8654),
            .I(N__8648));
    Odrv4 I__1904 (
            .O(N__8651),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    LocalMux I__1903 (
            .O(N__8648),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    InMux I__1902 (
            .O(N__8643),
            .I(N__8639));
    InMux I__1901 (
            .O(N__8642),
            .I(N__8636));
    LocalMux I__1900 (
            .O(N__8639),
            .I(N__8633));
    LocalMux I__1899 (
            .O(N__8636),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    Odrv4 I__1898 (
            .O(N__8633),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    InMux I__1897 (
            .O(N__8628),
            .I(N__8625));
    LocalMux I__1896 (
            .O(N__8625),
            .I(\U409_TICK.TICK603_11 ));
    InMux I__1895 (
            .O(N__8622),
            .I(N__8618));
    InMux I__1894 (
            .O(N__8621),
            .I(N__8615));
    LocalMux I__1893 (
            .O(N__8618),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    LocalMux I__1892 (
            .O(N__8615),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    CascadeMux I__1891 (
            .O(N__8610),
            .I(\U409_TICK.TICK603_8_cascade_ ));
    InMux I__1890 (
            .O(N__8607),
            .I(N__8604));
    LocalMux I__1889 (
            .O(N__8604),
            .I(N__8600));
    InMux I__1888 (
            .O(N__8603),
            .I(N__8597));
    Odrv4 I__1887 (
            .O(N__8600),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    LocalMux I__1886 (
            .O(N__8597),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    CascadeMux I__1885 (
            .O(N__8592),
            .I(\U409_TICK.TICK603_14_cascade_ ));
    CascadeMux I__1884 (
            .O(N__8589),
            .I(N__8586));
    InMux I__1883 (
            .O(N__8586),
            .I(N__8580));
    InMux I__1882 (
            .O(N__8585),
            .I(N__8577));
    InMux I__1881 (
            .O(N__8584),
            .I(N__8572));
    InMux I__1880 (
            .O(N__8583),
            .I(N__8572));
    LocalMux I__1879 (
            .O(N__8580),
            .I(N__8569));
    LocalMux I__1878 (
            .O(N__8577),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__1877 (
            .O(N__8572),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    Odrv4 I__1876 (
            .O(N__8569),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    CascadeMux I__1875 (
            .O(N__8562),
            .I(N__8559));
    InMux I__1874 (
            .O(N__8559),
            .I(N__8553));
    InMux I__1873 (
            .O(N__8558),
            .I(N__8553));
    LocalMux I__1872 (
            .O(N__8553),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    InMux I__1871 (
            .O(N__8550),
            .I(N__8541));
    InMux I__1870 (
            .O(N__8549),
            .I(N__8541));
    InMux I__1869 (
            .O(N__8548),
            .I(N__8541));
    LocalMux I__1868 (
            .O(N__8541),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    InMux I__1867 (
            .O(N__8538),
            .I(N__8532));
    InMux I__1866 (
            .O(N__8537),
            .I(N__8525));
    InMux I__1865 (
            .O(N__8536),
            .I(N__8525));
    InMux I__1864 (
            .O(N__8535),
            .I(N__8525));
    LocalMux I__1863 (
            .O(N__8532),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__1862 (
            .O(N__8525),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    InMux I__1861 (
            .O(N__8520),
            .I(N__8515));
    InMux I__1860 (
            .O(N__8519),
            .I(N__8510));
    InMux I__1859 (
            .O(N__8518),
            .I(N__8510));
    LocalMux I__1858 (
            .O(N__8515),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__1857 (
            .O(N__8510),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    InMux I__1856 (
            .O(N__8505),
            .I(\U409_TICK.un3_COUNTER60_1_cry_11 ));
    InMux I__1855 (
            .O(N__8502),
            .I(\U409_TICK.un3_COUNTER60_1_cry_12 ));
    InMux I__1854 (
            .O(N__8499),
            .I(\U409_TICK.un3_COUNTER60_1_cry_13 ));
    InMux I__1853 (
            .O(N__8496),
            .I(\U409_TICK.un3_COUNTER60_1_cry_14 ));
    InMux I__1852 (
            .O(N__8493),
            .I(\U409_TICK.un3_COUNTER60_1_cry_15 ));
    InMux I__1851 (
            .O(N__8490),
            .I(N__8487));
    LocalMux I__1850 (
            .O(N__8487),
            .I(N__8484));
    Odrv12 I__1849 (
            .O(N__8484),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ));
    CascadeMux I__1848 (
            .O(N__8481),
            .I(N__8478));
    InMux I__1847 (
            .O(N__8478),
            .I(N__8475));
    LocalMux I__1846 (
            .O(N__8475),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ));
    InMux I__1845 (
            .O(N__8472),
            .I(N__8469));
    LocalMux I__1844 (
            .O(N__8469),
            .I(N__8466));
    Odrv4 I__1843 (
            .O(N__8466),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ));
    InMux I__1842 (
            .O(N__8463),
            .I(N__8459));
    InMux I__1841 (
            .O(N__8462),
            .I(N__8456));
    LocalMux I__1840 (
            .O(N__8459),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    LocalMux I__1839 (
            .O(N__8456),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    InMux I__1838 (
            .O(N__8451),
            .I(N__8448));
    LocalMux I__1837 (
            .O(N__8448),
            .I(N__8444));
    InMux I__1836 (
            .O(N__8447),
            .I(N__8441));
    Odrv4 I__1835 (
            .O(N__8444),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    LocalMux I__1834 (
            .O(N__8441),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    CascadeMux I__1833 (
            .O(N__8436),
            .I(N__8432));
    InMux I__1832 (
            .O(N__8435),
            .I(N__8429));
    InMux I__1831 (
            .O(N__8432),
            .I(N__8426));
    LocalMux I__1830 (
            .O(N__8429),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    LocalMux I__1829 (
            .O(N__8426),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    InMux I__1828 (
            .O(N__8421),
            .I(N__8416));
    InMux I__1827 (
            .O(N__8420),
            .I(N__8413));
    InMux I__1826 (
            .O(N__8419),
            .I(N__8410));
    LocalMux I__1825 (
            .O(N__8416),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__1824 (
            .O(N__8413),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__1823 (
            .O(N__8410),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    InMux I__1822 (
            .O(N__8403),
            .I(\U409_TICK.un3_COUNTER60_1_cry_2 ));
    InMux I__1821 (
            .O(N__8400),
            .I(\U409_TICK.un3_COUNTER60_1_cry_3 ));
    InMux I__1820 (
            .O(N__8397),
            .I(\U409_TICK.un3_COUNTER60_1_cry_4 ));
    InMux I__1819 (
            .O(N__8394),
            .I(\U409_TICK.un3_COUNTER60_1_cry_5 ));
    InMux I__1818 (
            .O(N__8391),
            .I(\U409_TICK.un3_COUNTER60_1_cry_6 ));
    InMux I__1817 (
            .O(N__8388),
            .I(\U409_TICK.un3_COUNTER60_1_cry_7 ));
    InMux I__1816 (
            .O(N__8385),
            .I(N__8382));
    LocalMux I__1815 (
            .O(N__8382),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ));
    InMux I__1814 (
            .O(N__8379),
            .I(bfn_13_7_0_));
    InMux I__1813 (
            .O(N__8376),
            .I(\U409_TICK.un3_COUNTER60_1_cry_9 ));
    InMux I__1812 (
            .O(N__8373),
            .I(\U409_TICK.un3_COUNTER60_1_cry_10 ));
    InMux I__1811 (
            .O(N__8370),
            .I(N__8364));
    InMux I__1810 (
            .O(N__8369),
            .I(N__8361));
    InMux I__1809 (
            .O(N__8368),
            .I(N__8358));
    InMux I__1808 (
            .O(N__8367),
            .I(N__8355));
    LocalMux I__1807 (
            .O(N__8364),
            .I(N__8350));
    LocalMux I__1806 (
            .O(N__8361),
            .I(N__8350));
    LocalMux I__1805 (
            .O(N__8358),
            .I(N__8345));
    LocalMux I__1804 (
            .O(N__8355),
            .I(N__8340));
    Span4Mux_v I__1803 (
            .O(N__8350),
            .I(N__8340));
    InMux I__1802 (
            .O(N__8349),
            .I(N__8337));
    InMux I__1801 (
            .O(N__8348),
            .I(N__8334));
    Span4Mux_v I__1800 (
            .O(N__8345),
            .I(N__8331));
    Span4Mux_h I__1799 (
            .O(N__8340),
            .I(N__8326));
    LocalMux I__1798 (
            .O(N__8337),
            .I(N__8326));
    LocalMux I__1797 (
            .O(N__8334),
            .I(N__8321));
    Sp12to4 I__1796 (
            .O(N__8331),
            .I(N__8321));
    Span4Mux_h I__1795 (
            .O(N__8326),
            .I(N__8318));
    Span12Mux_h I__1794 (
            .O(N__8321),
            .I(N__8313));
    Sp12to4 I__1793 (
            .O(N__8318),
            .I(N__8313));
    Span12Mux_v I__1792 (
            .O(N__8313),
            .I(N__8310));
    Odrv12 I__1791 (
            .O(N__8310),
            .I(TSn_c));
    CascadeMux I__1790 (
            .O(N__8307),
            .I(N__8298));
    CascadeMux I__1789 (
            .O(N__8306),
            .I(N__8295));
    InMux I__1788 (
            .O(N__8305),
            .I(N__8292));
    InMux I__1787 (
            .O(N__8304),
            .I(N__8289));
    InMux I__1786 (
            .O(N__8303),
            .I(N__8286));
    InMux I__1785 (
            .O(N__8302),
            .I(N__8283));
    InMux I__1784 (
            .O(N__8301),
            .I(N__8280));
    InMux I__1783 (
            .O(N__8298),
            .I(N__8277));
    InMux I__1782 (
            .O(N__8295),
            .I(N__8274));
    LocalMux I__1781 (
            .O(N__8292),
            .I(N__8271));
    LocalMux I__1780 (
            .O(N__8289),
            .I(N__8259));
    LocalMux I__1779 (
            .O(N__8286),
            .I(N__8256));
    LocalMux I__1778 (
            .O(N__8283),
            .I(N__8253));
    LocalMux I__1777 (
            .O(N__8280),
            .I(N__8250));
    LocalMux I__1776 (
            .O(N__8277),
            .I(N__8247));
    LocalMux I__1775 (
            .O(N__8274),
            .I(N__8244));
    Glb2LocalMux I__1774 (
            .O(N__8271),
            .I(N__8211));
    ClkMux I__1773 (
            .O(N__8270),
            .I(N__8211));
    ClkMux I__1772 (
            .O(N__8269),
            .I(N__8211));
    ClkMux I__1771 (
            .O(N__8268),
            .I(N__8211));
    ClkMux I__1770 (
            .O(N__8267),
            .I(N__8211));
    ClkMux I__1769 (
            .O(N__8266),
            .I(N__8211));
    ClkMux I__1768 (
            .O(N__8265),
            .I(N__8211));
    ClkMux I__1767 (
            .O(N__8264),
            .I(N__8211));
    ClkMux I__1766 (
            .O(N__8263),
            .I(N__8211));
    ClkMux I__1765 (
            .O(N__8262),
            .I(N__8211));
    Glb2LocalMux I__1764 (
            .O(N__8259),
            .I(N__8211));
    Glb2LocalMux I__1763 (
            .O(N__8256),
            .I(N__8211));
    Glb2LocalMux I__1762 (
            .O(N__8253),
            .I(N__8211));
    Glb2LocalMux I__1761 (
            .O(N__8250),
            .I(N__8211));
    Glb2LocalMux I__1760 (
            .O(N__8247),
            .I(N__8211));
    Glb2LocalMux I__1759 (
            .O(N__8244),
            .I(N__8211));
    GlobalMux I__1758 (
            .O(N__8211),
            .I(N__8208));
    gio2CtrlBuf I__1757 (
            .O(N__8208),
            .I(CLK40_IN_c_g));
    InMux I__1756 (
            .O(N__8205),
            .I(N__8201));
    InMux I__1755 (
            .O(N__8204),
            .I(N__8198));
    LocalMux I__1754 (
            .O(N__8201),
            .I(\U409_TRANSFER_ACK.N_87 ));
    LocalMux I__1753 (
            .O(N__8198),
            .I(\U409_TRANSFER_ACK.N_87 ));
    CascadeMux I__1752 (
            .O(N__8193),
            .I(N__8187));
    CascadeMux I__1751 (
            .O(N__8192),
            .I(N__8184));
    InMux I__1750 (
            .O(N__8191),
            .I(N__8181));
    InMux I__1749 (
            .O(N__8190),
            .I(N__8174));
    InMux I__1748 (
            .O(N__8187),
            .I(N__8174));
    InMux I__1747 (
            .O(N__8184),
            .I(N__8174));
    LocalMux I__1746 (
            .O(N__8181),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__1745 (
            .O(N__8174),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    IoInMux I__1744 (
            .O(N__8169),
            .I(N__8166));
    LocalMux I__1743 (
            .O(N__8166),
            .I(N__8163));
    Span12Mux_s1_v I__1742 (
            .O(N__8163),
            .I(N__8160));
    Odrv12 I__1741 (
            .O(N__8160),
            .I(RESETn_c_i));
    InMux I__1740 (
            .O(N__8157),
            .I(\U409_TICK.un3_COUNTER60_1_cry_1 ));
    InMux I__1739 (
            .O(N__8154),
            .I(N__8150));
    InMux I__1738 (
            .O(N__8153),
            .I(N__8147));
    LocalMux I__1737 (
            .O(N__8150),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    LocalMux I__1736 (
            .O(N__8147),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    CascadeMux I__1735 (
            .O(N__8142),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3_cascade_ ));
    CascadeMux I__1734 (
            .O(N__8139),
            .I(N__8136));
    InMux I__1733 (
            .O(N__8136),
            .I(N__8130));
    InMux I__1732 (
            .O(N__8135),
            .I(N__8130));
    LocalMux I__1731 (
            .O(N__8130),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ));
    InMux I__1730 (
            .O(N__8127),
            .I(N__8124));
    LocalMux I__1729 (
            .O(N__8124),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a3_3 ));
    CascadeMux I__1728 (
            .O(N__8121),
            .I(\U409_TRANSFER_ACK.N_87_cascade_ ));
    InMux I__1727 (
            .O(N__8118),
            .I(N__8114));
    InMux I__1726 (
            .O(N__8117),
            .I(N__8111));
    LocalMux I__1725 (
            .O(N__8114),
            .I(\U409_TRANSFER_ACK.N_77 ));
    LocalMux I__1724 (
            .O(N__8111),
            .I(\U409_TRANSFER_ACK.N_77 ));
    CascadeMux I__1723 (
            .O(N__8106),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ));
    InMux I__1722 (
            .O(N__8103),
            .I(N__8094));
    InMux I__1721 (
            .O(N__8102),
            .I(N__8094));
    InMux I__1720 (
            .O(N__8101),
            .I(N__8094));
    LocalMux I__1719 (
            .O(N__8094),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    CascadeMux I__1718 (
            .O(N__8091),
            .I(\U409_TRANSFER_ACK.N_17_mux_cascade_ ));
    CascadeMux I__1717 (
            .O(N__8088),
            .I(\U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_ ));
    CascadeMux I__1716 (
            .O(N__8085),
            .I(\U409_TRANSFER_ACK.N_6_0_cascade_ ));
    InMux I__1715 (
            .O(N__8082),
            .I(N__8079));
    LocalMux I__1714 (
            .O(N__8079),
            .I(\U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0 ));
    InMux I__1713 (
            .O(N__8076),
            .I(N__8070));
    InMux I__1712 (
            .O(N__8075),
            .I(N__8070));
    LocalMux I__1711 (
            .O(N__8070),
            .I(\U409_TRANSFER_ACK.N_3_0 ));
    CascadeMux I__1710 (
            .O(N__8067),
            .I(N__8061));
    CascadeMux I__1709 (
            .O(N__8066),
            .I(N__8058));
    InMux I__1708 (
            .O(N__8065),
            .I(N__8054));
    InMux I__1707 (
            .O(N__8064),
            .I(N__8045));
    InMux I__1706 (
            .O(N__8061),
            .I(N__8045));
    InMux I__1705 (
            .O(N__8058),
            .I(N__8045));
    InMux I__1704 (
            .O(N__8057),
            .I(N__8045));
    LocalMux I__1703 (
            .O(N__8054),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__1702 (
            .O(N__8045),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    InMux I__1701 (
            .O(N__8040),
            .I(N__8037));
    LocalMux I__1700 (
            .O(N__8037),
            .I(\U409_TRANSFER_ACK.N_17_mux ));
    CascadeMux I__1699 (
            .O(N__8034),
            .I(N__8029));
    InMux I__1698 (
            .O(N__8033),
            .I(N__8024));
    InMux I__1697 (
            .O(N__8032),
            .I(N__8024));
    InMux I__1696 (
            .O(N__8029),
            .I(N__8021));
    LocalMux I__1695 (
            .O(N__8024),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__1694 (
            .O(N__8021),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    InMux I__1693 (
            .O(N__8016),
            .I(N__8012));
    InMux I__1692 (
            .O(N__8015),
            .I(N__8009));
    LocalMux I__1691 (
            .O(N__8012),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    LocalMux I__1690 (
            .O(N__8009),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    InMux I__1689 (
            .O(N__8004),
            .I(N__7998));
    InMux I__1688 (
            .O(N__8003),
            .I(N__7991));
    InMux I__1687 (
            .O(N__8002),
            .I(N__7991));
    InMux I__1686 (
            .O(N__8001),
            .I(N__7991));
    LocalMux I__1685 (
            .O(N__7998),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    LocalMux I__1684 (
            .O(N__7991),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    CascadeMux I__1683 (
            .O(N__7986),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ));
    IoInMux I__1682 (
            .O(N__7983),
            .I(N__7979));
    IoInMux I__1681 (
            .O(N__7982),
            .I(N__7976));
    LocalMux I__1680 (
            .O(N__7979),
            .I(N__7970));
    LocalMux I__1679 (
            .O(N__7976),
            .I(N__7970));
    IoInMux I__1678 (
            .O(N__7975),
            .I(N__7967));
    IoSpan4Mux I__1677 (
            .O(N__7970),
            .I(N__7964));
    LocalMux I__1676 (
            .O(N__7967),
            .I(N__7961));
    Span4Mux_s3_v I__1675 (
            .O(N__7964),
            .I(N__7958));
    Span4Mux_s3_v I__1674 (
            .O(N__7961),
            .I(N__7955));
    Sp12to4 I__1673 (
            .O(N__7958),
            .I(N__7950));
    Sp12to4 I__1672 (
            .O(N__7955),
            .I(N__7950));
    Span12Mux_s9_h I__1671 (
            .O(N__7950),
            .I(N__7947));
    Span12Mux_v I__1670 (
            .O(N__7947),
            .I(N__7942));
    InMux I__1669 (
            .O(N__7946),
            .I(N__7937));
    InMux I__1668 (
            .O(N__7945),
            .I(N__7937));
    Odrv12 I__1667 (
            .O(N__7942),
            .I(TACK_OUTn));
    LocalMux I__1666 (
            .O(N__7937),
            .I(TACK_OUTn));
    InMux I__1665 (
            .O(N__7932),
            .I(N__7929));
    LocalMux I__1664 (
            .O(N__7929),
            .I(\U409_TRANSFER_ACK.TACK_OUTn_3_0 ));
    InMux I__1663 (
            .O(N__7926),
            .I(N__7922));
    InMux I__1662 (
            .O(N__7925),
            .I(N__7918));
    LocalMux I__1661 (
            .O(N__7922),
            .I(N__7915));
    CascadeMux I__1660 (
            .O(N__7921),
            .I(N__7910));
    LocalMux I__1659 (
            .O(N__7918),
            .I(N__7904));
    Span4Mux_v I__1658 (
            .O(N__7915),
            .I(N__7904));
    InMux I__1657 (
            .O(N__7914),
            .I(N__7901));
    InMux I__1656 (
            .O(N__7913),
            .I(N__7894));
    InMux I__1655 (
            .O(N__7910),
            .I(N__7894));
    InMux I__1654 (
            .O(N__7909),
            .I(N__7894));
    Odrv4 I__1653 (
            .O(N__7904),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1652 (
            .O(N__7901),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1651 (
            .O(N__7894),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    CascadeMux I__1650 (
            .O(N__7887),
            .I(N__7884));
    InMux I__1649 (
            .O(N__7884),
            .I(N__7881));
    LocalMux I__1648 (
            .O(N__7881),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20_2 ));
    InMux I__1647 (
            .O(N__7878),
            .I(N__7873));
    InMux I__1646 (
            .O(N__7877),
            .I(N__7870));
    CascadeMux I__1645 (
            .O(N__7876),
            .I(N__7866));
    LocalMux I__1644 (
            .O(N__7873),
            .I(N__7862));
    LocalMux I__1643 (
            .O(N__7870),
            .I(N__7859));
    InMux I__1642 (
            .O(N__7869),
            .I(N__7856));
    InMux I__1641 (
            .O(N__7866),
            .I(N__7851));
    InMux I__1640 (
            .O(N__7865),
            .I(N__7851));
    Odrv4 I__1639 (
            .O(N__7862),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    Odrv4 I__1638 (
            .O(N__7859),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1637 (
            .O(N__7856),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1636 (
            .O(N__7851),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    InMux I__1635 (
            .O(N__7842),
            .I(N__7838));
    InMux I__1634 (
            .O(N__7841),
            .I(N__7835));
    LocalMux I__1633 (
            .O(N__7838),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    LocalMux I__1632 (
            .O(N__7835),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    InMux I__1631 (
            .O(N__7830),
            .I(N__7826));
    InMux I__1630 (
            .O(N__7829),
            .I(N__7823));
    LocalMux I__1629 (
            .O(N__7826),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    LocalMux I__1628 (
            .O(N__7823),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    CascadeMux I__1627 (
            .O(N__7818),
            .I(N__7814));
    CascadeMux I__1626 (
            .O(N__7817),
            .I(N__7811));
    InMux I__1625 (
            .O(N__7814),
            .I(N__7808));
    InMux I__1624 (
            .O(N__7811),
            .I(N__7805));
    LocalMux I__1623 (
            .O(N__7808),
            .I(N__7800));
    LocalMux I__1622 (
            .O(N__7805),
            .I(N__7800));
    Span4Mux_h I__1621 (
            .O(N__7800),
            .I(N__7797));
    Odrv4 I__1620 (
            .O(N__7797),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz ));
    InMux I__1619 (
            .O(N__7794),
            .I(N__7790));
    InMux I__1618 (
            .O(N__7793),
            .I(N__7787));
    LocalMux I__1617 (
            .O(N__7790),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    LocalMux I__1616 (
            .O(N__7787),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    InMux I__1615 (
            .O(N__7782),
            .I(N__7779));
    LocalMux I__1614 (
            .O(N__7779),
            .I(N__7776));
    Sp12to4 I__1613 (
            .O(N__7776),
            .I(N__7773));
    Span12Mux_h I__1612 (
            .O(N__7773),
            .I(N__7770));
    Span12Mux_v I__1611 (
            .O(N__7770),
            .I(N__7767));
    Odrv12 I__1610 (
            .O(N__7767),
            .I(TACKn_in));
    InMux I__1609 (
            .O(N__7764),
            .I(N__7761));
    LocalMux I__1608 (
            .O(N__7761),
            .I(N__7757));
    InMux I__1607 (
            .O(N__7760),
            .I(N__7754));
    Span4Mux_v I__1606 (
            .O(N__7757),
            .I(N__7750));
    LocalMux I__1605 (
            .O(N__7754),
            .I(N__7747));
    InMux I__1604 (
            .O(N__7753),
            .I(N__7744));
    Odrv4 I__1603 (
            .O(N__7750),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0 ));
    Odrv4 I__1602 (
            .O(N__7747),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0 ));
    LocalMux I__1601 (
            .O(N__7744),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0 ));
    CascadeMux I__1600 (
            .O(N__7737),
            .I(N__7733));
    CascadeMux I__1599 (
            .O(N__7736),
            .I(N__7730));
    InMux I__1598 (
            .O(N__7733),
            .I(N__7725));
    InMux I__1597 (
            .O(N__7730),
            .I(N__7725));
    LocalMux I__1596 (
            .O(N__7725),
            .I(N__7721));
    InMux I__1595 (
            .O(N__7724),
            .I(N__7718));
    Odrv12 I__1594 (
            .O(N__7721),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn));
    LocalMux I__1593 (
            .O(N__7718),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn));
    InMux I__1592 (
            .O(N__7713),
            .I(N__7707));
    InMux I__1591 (
            .O(N__7712),
            .I(N__7707));
    LocalMux I__1590 (
            .O(N__7707),
            .I(U409_ADDRESS_DECODE_un1_RAMSPACEn));
    IoInMux I__1589 (
            .O(N__7704),
            .I(N__7701));
    LocalMux I__1588 (
            .O(N__7701),
            .I(N__7698));
    Span12Mux_s1_v I__1587 (
            .O(N__7698),
            .I(N__7695));
    Span12Mux_v I__1586 (
            .O(N__7695),
            .I(N__7692));
    Odrv12 I__1585 (
            .O(N__7692),
            .I(BUFENn_c));
    InMux I__1584 (
            .O(N__7689),
            .I(N__7686));
    LocalMux I__1583 (
            .O(N__7686),
            .I(N__7683));
    Odrv4 I__1582 (
            .O(N__7683),
            .I(\U409_TRANSFER_ACK.N_119 ));
    IoInMux I__1581 (
            .O(N__7680),
            .I(N__7677));
    LocalMux I__1580 (
            .O(N__7677),
            .I(N__7674));
    Span4Mux_s3_v I__1579 (
            .O(N__7674),
            .I(N__7671));
    Span4Mux_h I__1578 (
            .O(N__7671),
            .I(N__7668));
    Odrv4 I__1577 (
            .O(N__7668),
            .I(GB_BUFFER_CLK40_IN_c_g_THRU_CO));
    IoInMux I__1576 (
            .O(N__7665),
            .I(N__7661));
    IoInMux I__1575 (
            .O(N__7664),
            .I(N__7658));
    LocalMux I__1574 (
            .O(N__7661),
            .I(N__7655));
    LocalMux I__1573 (
            .O(N__7658),
            .I(N__7652));
    Span4Mux_s0_v I__1572 (
            .O(N__7655),
            .I(N__7649));
    IoSpan4Mux I__1571 (
            .O(N__7652),
            .I(N__7646));
    Span4Mux_v I__1570 (
            .O(N__7649),
            .I(N__7643));
    Span4Mux_s3_h I__1569 (
            .O(N__7646),
            .I(N__7640));
    Span4Mux_v I__1568 (
            .O(N__7643),
            .I(N__7637));
    Sp12to4 I__1567 (
            .O(N__7640),
            .I(N__7634));
    Span4Mux_v I__1566 (
            .O(N__7637),
            .I(N__7631));
    Odrv12 I__1565 (
            .O(N__7634),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1564 (
            .O(N__7631),
            .I(CONSTANT_ONE_NET));
    InMux I__1563 (
            .O(N__7626),
            .I(N__7619));
    InMux I__1562 (
            .O(N__7625),
            .I(N__7616));
    InMux I__1561 (
            .O(N__7624),
            .I(N__7609));
    InMux I__1560 (
            .O(N__7623),
            .I(N__7609));
    InMux I__1559 (
            .O(N__7622),
            .I(N__7609));
    LocalMux I__1558 (
            .O(N__7619),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1557 (
            .O(N__7616),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1556 (
            .O(N__7609),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    InMux I__1555 (
            .O(N__7602),
            .I(N__7593));
    InMux I__1554 (
            .O(N__7601),
            .I(N__7593));
    InMux I__1553 (
            .O(N__7600),
            .I(N__7590));
    InMux I__1552 (
            .O(N__7599),
            .I(N__7585));
    InMux I__1551 (
            .O(N__7598),
            .I(N__7585));
    LocalMux I__1550 (
            .O(N__7593),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1549 (
            .O(N__7590),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1548 (
            .O(N__7585),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    IoInMux I__1547 (
            .O(N__7578),
            .I(N__7575));
    LocalMux I__1546 (
            .O(N__7575),
            .I(N__7572));
    Span4Mux_s3_v I__1545 (
            .O(N__7572),
            .I(N__7569));
    Sp12to4 I__1544 (
            .O(N__7569),
            .I(N__7566));
    Span12Mux_h I__1543 (
            .O(N__7566),
            .I(N__7563));
    Odrv12 I__1542 (
            .O(N__7563),
            .I(ROMENn_c));
    CEMux I__1541 (
            .O(N__7560),
            .I(N__7557));
    LocalMux I__1540 (
            .O(N__7557),
            .I(N__7554));
    Span4Mux_h I__1539 (
            .O(N__7554),
            .I(N__7551));
    Odrv4 I__1538 (
            .O(N__7551),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_0 ));
    InMux I__1537 (
            .O(N__7548),
            .I(N__7545));
    LocalMux I__1536 (
            .O(N__7545),
            .I(N__7541));
    InMux I__1535 (
            .O(N__7544),
            .I(N__7538));
    Span4Mux_h I__1534 (
            .O(N__7541),
            .I(N__7535));
    LocalMux I__1533 (
            .O(N__7538),
            .I(AC_TACK));
    Odrv4 I__1532 (
            .O(N__7535),
            .I(AC_TACK));
    CascadeMux I__1531 (
            .O(N__7530),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_ ));
    InMux I__1530 (
            .O(N__7527),
            .I(N__7523));
    InMux I__1529 (
            .O(N__7526),
            .I(N__7520));
    LocalMux I__1528 (
            .O(N__7523),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    LocalMux I__1527 (
            .O(N__7520),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    InMux I__1526 (
            .O(N__7515),
            .I(N__7509));
    InMux I__1525 (
            .O(N__7514),
            .I(N__7502));
    InMux I__1524 (
            .O(N__7513),
            .I(N__7502));
    InMux I__1523 (
            .O(N__7512),
            .I(N__7502));
    LocalMux I__1522 (
            .O(N__7509),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    LocalMux I__1521 (
            .O(N__7502),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    CascadeMux I__1520 (
            .O(N__7497),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_cascade_ ));
    CascadeMux I__1519 (
            .O(N__7494),
            .I(N__7491));
    InMux I__1518 (
            .O(N__7491),
            .I(N__7488));
    LocalMux I__1517 (
            .O(N__7488),
            .I(N__7485));
    Span4Mux_v I__1516 (
            .O(N__7485),
            .I(N__7481));
    InMux I__1515 (
            .O(N__7484),
            .I(N__7478));
    Span4Mux_h I__1514 (
            .O(N__7481),
            .I(N__7475));
    LocalMux I__1513 (
            .O(N__7478),
            .I(N__7472));
    Sp12to4 I__1512 (
            .O(N__7475),
            .I(N__7467));
    Span12Mux_h I__1511 (
            .O(N__7472),
            .I(N__7467));
    Span12Mux_v I__1510 (
            .O(N__7467),
            .I(N__7464));
    Odrv12 I__1509 (
            .O(N__7464),
            .I(D_in_4));
    InMux I__1508 (
            .O(N__7461),
            .I(N__7457));
    InMux I__1507 (
            .O(N__7460),
            .I(N__7454));
    LocalMux I__1506 (
            .O(N__7457),
            .I(ATA_BASE_4));
    LocalMux I__1505 (
            .O(N__7454),
            .I(ATA_BASE_4));
    CascadeMux I__1504 (
            .O(N__7449),
            .I(N__7446));
    InMux I__1503 (
            .O(N__7446),
            .I(N__7443));
    LocalMux I__1502 (
            .O(N__7443),
            .I(N__7440));
    Span4Mux_v I__1501 (
            .O(N__7440),
            .I(N__7436));
    InMux I__1500 (
            .O(N__7439),
            .I(N__7433));
    Span4Mux_v I__1499 (
            .O(N__7436),
            .I(N__7429));
    LocalMux I__1498 (
            .O(N__7433),
            .I(N__7426));
    CascadeMux I__1497 (
            .O(N__7432),
            .I(N__7423));
    Span4Mux_v I__1496 (
            .O(N__7429),
            .I(N__7420));
    Span4Mux_h I__1495 (
            .O(N__7426),
            .I(N__7417));
    InMux I__1494 (
            .O(N__7423),
            .I(N__7414));
    Sp12to4 I__1493 (
            .O(N__7420),
            .I(N__7411));
    Sp12to4 I__1492 (
            .O(N__7417),
            .I(N__7406));
    LocalMux I__1491 (
            .O(N__7414),
            .I(N__7406));
    Span12Mux_h I__1490 (
            .O(N__7411),
            .I(N__7401));
    Span12Mux_v I__1489 (
            .O(N__7406),
            .I(N__7401));
    Odrv12 I__1488 (
            .O(N__7401),
            .I(D_in_5));
    InMux I__1487 (
            .O(N__7398),
            .I(N__7394));
    InMux I__1486 (
            .O(N__7397),
            .I(N__7391));
    LocalMux I__1485 (
            .O(N__7394),
            .I(ATA_BASE_5));
    LocalMux I__1484 (
            .O(N__7391),
            .I(ATA_BASE_5));
    InMux I__1483 (
            .O(N__7386),
            .I(N__7380));
    InMux I__1482 (
            .O(N__7385),
            .I(N__7373));
    InMux I__1481 (
            .O(N__7384),
            .I(N__7373));
    InMux I__1480 (
            .O(N__7383),
            .I(N__7373));
    LocalMux I__1479 (
            .O(N__7380),
            .I(\U409_AUTOCONFIG.LIDE_CONF_RNIUPP42Z0Z_1 ));
    LocalMux I__1478 (
            .O(N__7373),
            .I(\U409_AUTOCONFIG.LIDE_CONF_RNIUPP42Z0Z_1 ));
    InMux I__1477 (
            .O(N__7368),
            .I(N__7364));
    InMux I__1476 (
            .O(N__7367),
            .I(N__7361));
    LocalMux I__1475 (
            .O(N__7364),
            .I(ATA_BASE_6));
    LocalMux I__1474 (
            .O(N__7361),
            .I(ATA_BASE_6));
    CascadeMux I__1473 (
            .O(N__7356),
            .I(N__7348));
    InMux I__1472 (
            .O(N__7355),
            .I(N__7339));
    InMux I__1471 (
            .O(N__7354),
            .I(N__7339));
    InMux I__1470 (
            .O(N__7353),
            .I(N__7339));
    InMux I__1469 (
            .O(N__7352),
            .I(N__7327));
    InMux I__1468 (
            .O(N__7351),
            .I(N__7327));
    InMux I__1467 (
            .O(N__7348),
            .I(N__7327));
    InMux I__1466 (
            .O(N__7347),
            .I(N__7327));
    InMux I__1465 (
            .O(N__7346),
            .I(N__7327));
    LocalMux I__1464 (
            .O(N__7339),
            .I(N__7322));
    InMux I__1463 (
            .O(N__7338),
            .I(N__7319));
    LocalMux I__1462 (
            .O(N__7327),
            .I(N__7316));
    InMux I__1461 (
            .O(N__7326),
            .I(N__7311));
    InMux I__1460 (
            .O(N__7325),
            .I(N__7311));
    Span4Mux_h I__1459 (
            .O(N__7322),
            .I(N__7308));
    LocalMux I__1458 (
            .O(N__7319),
            .I(N__7305));
    Span4Mux_h I__1457 (
            .O(N__7316),
            .I(N__7300));
    LocalMux I__1456 (
            .O(N__7311),
            .I(N__7300));
    Odrv4 I__1455 (
            .O(N__7308),
            .I(un1_AUTOCONFIG_SPACE));
    Odrv4 I__1454 (
            .O(N__7305),
            .I(un1_AUTOCONFIG_SPACE));
    Odrv4 I__1453 (
            .O(N__7300),
            .I(un1_AUTOCONFIG_SPACE));
    InMux I__1452 (
            .O(N__7293),
            .I(N__7288));
    InMux I__1451 (
            .O(N__7292),
            .I(N__7283));
    InMux I__1450 (
            .O(N__7291),
            .I(N__7283));
    LocalMux I__1449 (
            .O(N__7288),
            .I(\U409_AUTOCONFIG.LIDE_CONF_RNIUPP42Z0Z_0 ));
    LocalMux I__1448 (
            .O(N__7283),
            .I(\U409_AUTOCONFIG.LIDE_CONF_RNIUPP42Z0Z_0 ));
    CascadeMux I__1447 (
            .O(N__7278),
            .I(N__7274));
    CascadeMux I__1446 (
            .O(N__7277),
            .I(N__7271));
    InMux I__1445 (
            .O(N__7274),
            .I(N__7268));
    InMux I__1444 (
            .O(N__7271),
            .I(N__7265));
    LocalMux I__1443 (
            .O(N__7268),
            .I(N__7259));
    LocalMux I__1442 (
            .O(N__7265),
            .I(N__7259));
    InMux I__1441 (
            .O(N__7264),
            .I(N__7256));
    Span4Mux_v I__1440 (
            .O(N__7259),
            .I(N__7253));
    LocalMux I__1439 (
            .O(N__7256),
            .I(N__7250));
    Sp12to4 I__1438 (
            .O(N__7253),
            .I(N__7247));
    Span4Mux_h I__1437 (
            .O(N__7250),
            .I(N__7244));
    Span12Mux_h I__1436 (
            .O(N__7247),
            .I(N__7239));
    Sp12to4 I__1435 (
            .O(N__7244),
            .I(N__7239));
    Span12Mux_v I__1434 (
            .O(N__7239),
            .I(N__7236));
    Odrv12 I__1433 (
            .O(N__7236),
            .I(D_in_6));
    InMux I__1432 (
            .O(N__7233),
            .I(N__7229));
    InMux I__1431 (
            .O(N__7232),
            .I(N__7226));
    LocalMux I__1430 (
            .O(N__7229),
            .I(ATA_BASE_2));
    LocalMux I__1429 (
            .O(N__7226),
            .I(ATA_BASE_2));
    CascadeMux I__1428 (
            .O(N__7221),
            .I(N__7217));
    InMux I__1427 (
            .O(N__7220),
            .I(N__7214));
    InMux I__1426 (
            .O(N__7217),
            .I(N__7211));
    LocalMux I__1425 (
            .O(N__7214),
            .I(N__7208));
    LocalMux I__1424 (
            .O(N__7211),
            .I(\U409_ADDRESS_DECODE.LOWROMZ0Z_3 ));
    Odrv4 I__1423 (
            .O(N__7208),
            .I(\U409_ADDRESS_DECODE.LOWROMZ0Z_3 ));
    InMux I__1422 (
            .O(N__7203),
            .I(N__7197));
    InMux I__1421 (
            .O(N__7202),
            .I(N__7197));
    LocalMux I__1420 (
            .O(N__7197),
            .I(N__7193));
    InMux I__1419 (
            .O(N__7196),
            .I(N__7190));
    Span4Mux_v I__1418 (
            .O(N__7193),
            .I(N__7186));
    LocalMux I__1417 (
            .O(N__7190),
            .I(N__7183));
    InMux I__1416 (
            .O(N__7189),
            .I(N__7180));
    Odrv4 I__1415 (
            .O(N__7186),
            .I(U409_ADDRESS_DECODE_ROMEN_1));
    Odrv12 I__1414 (
            .O(N__7183),
            .I(U409_ADDRESS_DECODE_ROMEN_1));
    LocalMux I__1413 (
            .O(N__7180),
            .I(U409_ADDRESS_DECODE_ROMEN_1));
    CascadeMux I__1412 (
            .O(N__7173),
            .I(N__7170));
    InMux I__1411 (
            .O(N__7170),
            .I(N__7163));
    InMux I__1410 (
            .O(N__7169),
            .I(N__7154));
    InMux I__1409 (
            .O(N__7168),
            .I(N__7154));
    InMux I__1408 (
            .O(N__7167),
            .I(N__7151));
    CascadeMux I__1407 (
            .O(N__7166),
            .I(N__7147));
    LocalMux I__1406 (
            .O(N__7163),
            .I(N__7143));
    InMux I__1405 (
            .O(N__7162),
            .I(N__7140));
    InMux I__1404 (
            .O(N__7161),
            .I(N__7137));
    InMux I__1403 (
            .O(N__7160),
            .I(N__7134));
    InMux I__1402 (
            .O(N__7159),
            .I(N__7131));
    LocalMux I__1401 (
            .O(N__7154),
            .I(N__7126));
    LocalMux I__1400 (
            .O(N__7151),
            .I(N__7126));
    InMux I__1399 (
            .O(N__7150),
            .I(N__7123));
    InMux I__1398 (
            .O(N__7147),
            .I(N__7120));
    InMux I__1397 (
            .O(N__7146),
            .I(N__7117));
    Span4Mux_v I__1396 (
            .O(N__7143),
            .I(N__7114));
    LocalMux I__1395 (
            .O(N__7140),
            .I(N__7105));
    LocalMux I__1394 (
            .O(N__7137),
            .I(N__7105));
    LocalMux I__1393 (
            .O(N__7134),
            .I(N__7105));
    LocalMux I__1392 (
            .O(N__7131),
            .I(N__7105));
    Span4Mux_v I__1391 (
            .O(N__7126),
            .I(N__7102));
    LocalMux I__1390 (
            .O(N__7123),
            .I(N__7095));
    LocalMux I__1389 (
            .O(N__7120),
            .I(N__7095));
    LocalMux I__1388 (
            .O(N__7117),
            .I(N__7095));
    Span4Mux_h I__1387 (
            .O(N__7114),
            .I(N__7090));
    Span4Mux_v I__1386 (
            .O(N__7105),
            .I(N__7090));
    Span4Mux_h I__1385 (
            .O(N__7102),
            .I(N__7085));
    Span4Mux_v I__1384 (
            .O(N__7095),
            .I(N__7085));
    Sp12to4 I__1383 (
            .O(N__7090),
            .I(N__7080));
    Sp12to4 I__1382 (
            .O(N__7085),
            .I(N__7080));
    Odrv12 I__1381 (
            .O(N__7080),
            .I(A_c_21));
    InMux I__1380 (
            .O(N__7077),
            .I(N__7074));
    LocalMux I__1379 (
            .O(N__7074),
            .I(N__7070));
    InMux I__1378 (
            .O(N__7073),
            .I(N__7067));
    Span4Mux_h I__1377 (
            .O(N__7070),
            .I(N__7061));
    LocalMux I__1376 (
            .O(N__7067),
            .I(N__7061));
    InMux I__1375 (
            .O(N__7066),
            .I(N__7058));
    Span4Mux_v I__1374 (
            .O(N__7061),
            .I(N__7055));
    LocalMux I__1373 (
            .O(N__7058),
            .I(N__7052));
    Sp12to4 I__1372 (
            .O(N__7055),
            .I(N__7049));
    Span12Mux_h I__1371 (
            .O(N__7052),
            .I(N__7046));
    Span12Mux_h I__1370 (
            .O(N__7049),
            .I(N__7043));
    Span12Mux_v I__1369 (
            .O(N__7046),
            .I(N__7040));
    Span12Mux_v I__1368 (
            .O(N__7043),
            .I(N__7037));
    Odrv12 I__1367 (
            .O(N__7040),
            .I(OVL_c));
    Odrv12 I__1366 (
            .O(N__7037),
            .I(OVL_c));
    InMux I__1365 (
            .O(N__7032),
            .I(N__7028));
    InMux I__1364 (
            .O(N__7031),
            .I(N__7024));
    LocalMux I__1363 (
            .O(N__7028),
            .I(N__7021));
    InMux I__1362 (
            .O(N__7027),
            .I(N__7018));
    LocalMux I__1361 (
            .O(N__7024),
            .I(N__7015));
    Span4Mux_h I__1360 (
            .O(N__7021),
            .I(N__7012));
    LocalMux I__1359 (
            .O(N__7018),
            .I(N__7009));
    Span12Mux_h I__1358 (
            .O(N__7015),
            .I(N__7006));
    Sp12to4 I__1357 (
            .O(N__7012),
            .I(N__7001));
    Sp12to4 I__1356 (
            .O(N__7009),
            .I(N__7001));
    Span12Mux_v I__1355 (
            .O(N__7006),
            .I(N__6998));
    Span12Mux_v I__1354 (
            .O(N__7001),
            .I(N__6995));
    Odrv12 I__1353 (
            .O(N__6998),
            .I(A_c_28));
    Odrv12 I__1352 (
            .O(N__6995),
            .I(A_c_28));
    CascadeMux I__1351 (
            .O(N__6990),
            .I(N__6987));
    InMux I__1350 (
            .O(N__6987),
            .I(N__6983));
    CascadeMux I__1349 (
            .O(N__6986),
            .I(N__6980));
    LocalMux I__1348 (
            .O(N__6983),
            .I(N__6977));
    InMux I__1347 (
            .O(N__6980),
            .I(N__6974));
    Odrv4 I__1346 (
            .O(N__6977),
            .I(BRIDGE_BASE_0));
    LocalMux I__1345 (
            .O(N__6974),
            .I(BRIDGE_BASE_0));
    InMux I__1344 (
            .O(N__6969),
            .I(N__6966));
    LocalMux I__1343 (
            .O(N__6966),
            .I(N__6963));
    Span4Mux_v I__1342 (
            .O(N__6963),
            .I(N__6960));
    Odrv4 I__1341 (
            .O(N__6960),
            .I(\U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_3 ));
    IoInMux I__1340 (
            .O(N__6957),
            .I(N__6954));
    LocalMux I__1339 (
            .O(N__6954),
            .I(N__6951));
    IoSpan4Mux I__1338 (
            .O(N__6951),
            .I(N__6948));
    Span4Mux_s3_h I__1337 (
            .O(N__6948),
            .I(N__6945));
    Sp12to4 I__1336 (
            .O(N__6945),
            .I(N__6942));
    Span12Mux_h I__1335 (
            .O(N__6942),
            .I(N__6939));
    Odrv12 I__1334 (
            .O(N__6939),
            .I(U409_ADDRESS_DECODE_un1_BRIDGE_ENn_i));
    CascadeMux I__1333 (
            .O(N__6936),
            .I(N__6933));
    InMux I__1332 (
            .O(N__6933),
            .I(N__6929));
    InMux I__1331 (
            .O(N__6932),
            .I(N__6926));
    LocalMux I__1330 (
            .O(N__6929),
            .I(N__6920));
    LocalMux I__1329 (
            .O(N__6926),
            .I(N__6917));
    InMux I__1328 (
            .O(N__6925),
            .I(N__6914));
    InMux I__1327 (
            .O(N__6924),
            .I(N__6911));
    InMux I__1326 (
            .O(N__6923),
            .I(N__6908));
    Span4Mux_v I__1325 (
            .O(N__6920),
            .I(N__6903));
    Span4Mux_v I__1324 (
            .O(N__6917),
            .I(N__6900));
    LocalMux I__1323 (
            .O(N__6914),
            .I(N__6897));
    LocalMux I__1322 (
            .O(N__6911),
            .I(N__6894));
    LocalMux I__1321 (
            .O(N__6908),
            .I(N__6890));
    InMux I__1320 (
            .O(N__6907),
            .I(N__6887));
    InMux I__1319 (
            .O(N__6906),
            .I(N__6884));
    Span4Mux_h I__1318 (
            .O(N__6903),
            .I(N__6875));
    Span4Mux_h I__1317 (
            .O(N__6900),
            .I(N__6875));
    Span4Mux_v I__1316 (
            .O(N__6897),
            .I(N__6875));
    Span4Mux_v I__1315 (
            .O(N__6894),
            .I(N__6875));
    InMux I__1314 (
            .O(N__6893),
            .I(N__6872));
    Span4Mux_v I__1313 (
            .O(N__6890),
            .I(N__6869));
    LocalMux I__1312 (
            .O(N__6887),
            .I(N__6866));
    LocalMux I__1311 (
            .O(N__6884),
            .I(N__6859));
    Sp12to4 I__1310 (
            .O(N__6875),
            .I(N__6859));
    LocalMux I__1309 (
            .O(N__6872),
            .I(N__6859));
    Sp12to4 I__1308 (
            .O(N__6869),
            .I(N__6854));
    Span12Mux_v I__1307 (
            .O(N__6866),
            .I(N__6854));
    Span12Mux_h I__1306 (
            .O(N__6859),
            .I(N__6851));
    Odrv12 I__1305 (
            .O(N__6854),
            .I(A_c_20));
    Odrv12 I__1304 (
            .O(N__6851),
            .I(A_c_20));
    InMux I__1303 (
            .O(N__6846),
            .I(N__6843));
    LocalMux I__1302 (
            .O(N__6843),
            .I(\U409_ADDRESS_DECODE.ATA_SPACE_1Z0Z_0 ));
    IoInMux I__1301 (
            .O(N__6840),
            .I(N__6837));
    LocalMux I__1300 (
            .O(N__6837),
            .I(N__6834));
    IoSpan4Mux I__1299 (
            .O(N__6834),
            .I(N__6831));
    Span4Mux_s2_v I__1298 (
            .O(N__6831),
            .I(N__6828));
    Sp12to4 I__1297 (
            .O(N__6828),
            .I(N__6825));
    Span12Mux_v I__1296 (
            .O(N__6825),
            .I(N__6822));
    Odrv12 I__1295 (
            .O(N__6822),
            .I(U409_ADDRESS_DECODE_un1_RAMSPACEn_i));
    InMux I__1294 (
            .O(N__6819),
            .I(N__6816));
    LocalMux I__1293 (
            .O(N__6816),
            .I(N__6813));
    Odrv12 I__1292 (
            .O(N__6813),
            .I(U409_ADDRESS_DECODE_un1_ROMEN_0));
    InMux I__1291 (
            .O(N__6810),
            .I(N__6807));
    LocalMux I__1290 (
            .O(N__6807),
            .I(N__6802));
    InMux I__1289 (
            .O(N__6806),
            .I(N__6799));
    InMux I__1288 (
            .O(N__6805),
            .I(N__6796));
    Odrv12 I__1287 (
            .O(N__6802),
            .I(\U409_ADDRESS_DECODE.ATA_ENZ0 ));
    LocalMux I__1286 (
            .O(N__6799),
            .I(\U409_ADDRESS_DECODE.ATA_ENZ0 ));
    LocalMux I__1285 (
            .O(N__6796),
            .I(\U409_ADDRESS_DECODE.ATA_ENZ0 ));
    IoInMux I__1284 (
            .O(N__6789),
            .I(N__6786));
    LocalMux I__1283 (
            .O(N__6786),
            .I(N__6783));
    IoSpan4Mux I__1282 (
            .O(N__6783),
            .I(N__6780));
    Sp12to4 I__1281 (
            .O(N__6780),
            .I(N__6777));
    Span12Mux_s7_h I__1280 (
            .O(N__6777),
            .I(N__6774));
    Span12Mux_h I__1279 (
            .O(N__6774),
            .I(N__6771));
    Odrv12 I__1278 (
            .O(N__6771),
            .I(U409_ADDRESS_DECODE_un1_ATA_ENn_i));
    InMux I__1277 (
            .O(N__6768),
            .I(N__6762));
    InMux I__1276 (
            .O(N__6767),
            .I(N__6762));
    LocalMux I__1275 (
            .O(N__6762),
            .I(\U409_TRANSFER_ACK.CO1 ));
    InMux I__1274 (
            .O(N__6759),
            .I(N__6755));
    InMux I__1273 (
            .O(N__6758),
            .I(N__6752));
    LocalMux I__1272 (
            .O(N__6755),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20 ));
    LocalMux I__1271 (
            .O(N__6752),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20 ));
    InMux I__1270 (
            .O(N__6747),
            .I(N__6741));
    InMux I__1269 (
            .O(N__6746),
            .I(N__6741));
    LocalMux I__1268 (
            .O(N__6741),
            .I(N__6738));
    Odrv4 I__1267 (
            .O(N__6738),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15 ));
    CascadeMux I__1266 (
            .O(N__6735),
            .I(N__6732));
    InMux I__1265 (
            .O(N__6732),
            .I(N__6728));
    InMux I__1264 (
            .O(N__6731),
            .I(N__6725));
    LocalMux I__1263 (
            .O(N__6728),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ));
    LocalMux I__1262 (
            .O(N__6725),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ));
    CascadeMux I__1261 (
            .O(N__6720),
            .I(N__6717));
    InMux I__1260 (
            .O(N__6717),
            .I(N__6711));
    InMux I__1259 (
            .O(N__6716),
            .I(N__6711));
    LocalMux I__1258 (
            .O(N__6711),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0 ));
    CascadeMux I__1257 (
            .O(N__6708),
            .I(N__6705));
    InMux I__1256 (
            .O(N__6705),
            .I(N__6702));
    LocalMux I__1255 (
            .O(N__6702),
            .I(N__6699));
    Span4Mux_v I__1254 (
            .O(N__6699),
            .I(N__6694));
    CascadeMux I__1253 (
            .O(N__6698),
            .I(N__6691));
    CascadeMux I__1252 (
            .O(N__6697),
            .I(N__6688));
    Span4Mux_h I__1251 (
            .O(N__6694),
            .I(N__6685));
    InMux I__1250 (
            .O(N__6691),
            .I(N__6680));
    InMux I__1249 (
            .O(N__6688),
            .I(N__6680));
    Sp12to4 I__1248 (
            .O(N__6685),
            .I(N__6677));
    LocalMux I__1247 (
            .O(N__6680),
            .I(N__6674));
    Span12Mux_h I__1246 (
            .O(N__6677),
            .I(N__6669));
    Span12Mux_h I__1245 (
            .O(N__6674),
            .I(N__6669));
    Span12Mux_v I__1244 (
            .O(N__6669),
            .I(N__6666));
    Odrv12 I__1243 (
            .O(N__6666),
            .I(D_in_7));
    InMux I__1242 (
            .O(N__6663),
            .I(N__6660));
    LocalMux I__1241 (
            .O(N__6660),
            .I(N__6656));
    InMux I__1240 (
            .O(N__6659),
            .I(N__6653));
    Odrv4 I__1239 (
            .O(N__6656),
            .I(BRIDGE_BASE_3));
    LocalMux I__1238 (
            .O(N__6653),
            .I(BRIDGE_BASE_3));
    InMux I__1237 (
            .O(N__6648),
            .I(N__6645));
    LocalMux I__1236 (
            .O(N__6645),
            .I(N__6641));
    CascadeMux I__1235 (
            .O(N__6644),
            .I(N__6638));
    Span4Mux_v I__1234 (
            .O(N__6641),
            .I(N__6635));
    InMux I__1233 (
            .O(N__6638),
            .I(N__6632));
    Odrv4 I__1232 (
            .O(N__6635),
            .I(BRIDGE_BASE_2));
    LocalMux I__1231 (
            .O(N__6632),
            .I(BRIDGE_BASE_2));
    InMux I__1230 (
            .O(N__6627),
            .I(N__6624));
    LocalMux I__1229 (
            .O(N__6624),
            .I(N__6621));
    Span12Mux_v I__1228 (
            .O(N__6621),
            .I(N__6617));
    InMux I__1227 (
            .O(N__6620),
            .I(N__6614));
    Odrv12 I__1226 (
            .O(N__6617),
            .I(BRIDGE_BASE_1));
    LocalMux I__1225 (
            .O(N__6614),
            .I(BRIDGE_BASE_1));
    InMux I__1224 (
            .O(N__6609),
            .I(N__6603));
    InMux I__1223 (
            .O(N__6608),
            .I(N__6596));
    InMux I__1222 (
            .O(N__6607),
            .I(N__6596));
    InMux I__1221 (
            .O(N__6606),
            .I(N__6596));
    LocalMux I__1220 (
            .O(N__6603),
            .I(\U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa ));
    LocalMux I__1219 (
            .O(N__6596),
            .I(\U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa ));
    InMux I__1218 (
            .O(N__6591),
            .I(N__6585));
    CascadeMux I__1217 (
            .O(N__6590),
            .I(N__6581));
    CascadeMux I__1216 (
            .O(N__6589),
            .I(N__6577));
    InMux I__1215 (
            .O(N__6588),
            .I(N__6570));
    LocalMux I__1214 (
            .O(N__6585),
            .I(N__6567));
    InMux I__1213 (
            .O(N__6584),
            .I(N__6564));
    InMux I__1212 (
            .O(N__6581),
            .I(N__6561));
    InMux I__1211 (
            .O(N__6580),
            .I(N__6558));
    InMux I__1210 (
            .O(N__6577),
            .I(N__6553));
    InMux I__1209 (
            .O(N__6576),
            .I(N__6553));
    InMux I__1208 (
            .O(N__6575),
            .I(N__6550));
    InMux I__1207 (
            .O(N__6574),
            .I(N__6547));
    InMux I__1206 (
            .O(N__6573),
            .I(N__6544));
    LocalMux I__1205 (
            .O(N__6570),
            .I(N__6541));
    Span4Mux_h I__1204 (
            .O(N__6567),
            .I(N__6528));
    LocalMux I__1203 (
            .O(N__6564),
            .I(N__6528));
    LocalMux I__1202 (
            .O(N__6561),
            .I(N__6528));
    LocalMux I__1201 (
            .O(N__6558),
            .I(N__6528));
    LocalMux I__1200 (
            .O(N__6553),
            .I(N__6528));
    LocalMux I__1199 (
            .O(N__6550),
            .I(N__6528));
    LocalMux I__1198 (
            .O(N__6547),
            .I(N__6523));
    LocalMux I__1197 (
            .O(N__6544),
            .I(N__6523));
    Span4Mux_v I__1196 (
            .O(N__6541),
            .I(N__6520));
    Span4Mux_v I__1195 (
            .O(N__6528),
            .I(N__6517));
    Span4Mux_v I__1194 (
            .O(N__6523),
            .I(N__6514));
    Sp12to4 I__1193 (
            .O(N__6520),
            .I(N__6507));
    Sp12to4 I__1192 (
            .O(N__6517),
            .I(N__6507));
    Sp12to4 I__1191 (
            .O(N__6514),
            .I(N__6507));
    Odrv12 I__1190 (
            .O(N__6507),
            .I(A_c_23));
    InMux I__1189 (
            .O(N__6504),
            .I(N__6500));
    InMux I__1188 (
            .O(N__6503),
            .I(N__6497));
    LocalMux I__1187 (
            .O(N__6500),
            .I(ATA_BASE_7));
    LocalMux I__1186 (
            .O(N__6497),
            .I(ATA_BASE_7));
    CascadeMux I__1185 (
            .O(N__6492),
            .I(N__6488));
    InMux I__1184 (
            .O(N__6491),
            .I(N__6482));
    InMux I__1183 (
            .O(N__6488),
            .I(N__6475));
    InMux I__1182 (
            .O(N__6487),
            .I(N__6472));
    InMux I__1181 (
            .O(N__6486),
            .I(N__6469));
    InMux I__1180 (
            .O(N__6485),
            .I(N__6466));
    LocalMux I__1179 (
            .O(N__6482),
            .I(N__6463));
    InMux I__1178 (
            .O(N__6481),
            .I(N__6460));
    InMux I__1177 (
            .O(N__6480),
            .I(N__6457));
    InMux I__1176 (
            .O(N__6479),
            .I(N__6454));
    CascadeMux I__1175 (
            .O(N__6478),
            .I(N__6451));
    LocalMux I__1174 (
            .O(N__6475),
            .I(N__6442));
    LocalMux I__1173 (
            .O(N__6472),
            .I(N__6442));
    LocalMux I__1172 (
            .O(N__6469),
            .I(N__6442));
    LocalMux I__1171 (
            .O(N__6466),
            .I(N__6442));
    Span4Mux_v I__1170 (
            .O(N__6463),
            .I(N__6439));
    LocalMux I__1169 (
            .O(N__6460),
            .I(N__6432));
    LocalMux I__1168 (
            .O(N__6457),
            .I(N__6432));
    LocalMux I__1167 (
            .O(N__6454),
            .I(N__6432));
    InMux I__1166 (
            .O(N__6451),
            .I(N__6429));
    Span4Mux_v I__1165 (
            .O(N__6442),
            .I(N__6426));
    Span4Mux_h I__1164 (
            .O(N__6439),
            .I(N__6421));
    Span4Mux_v I__1163 (
            .O(N__6432),
            .I(N__6421));
    LocalMux I__1162 (
            .O(N__6429),
            .I(N__6418));
    Span4Mux_v I__1161 (
            .O(N__6426),
            .I(N__6415));
    Span4Mux_v I__1160 (
            .O(N__6421),
            .I(N__6412));
    Span12Mux_h I__1159 (
            .O(N__6418),
            .I(N__6409));
    Span4Mux_v I__1158 (
            .O(N__6415),
            .I(N__6406));
    Span4Mux_v I__1157 (
            .O(N__6412),
            .I(N__6403));
    Span12Mux_v I__1156 (
            .O(N__6409),
            .I(N__6400));
    Sp12to4 I__1155 (
            .O(N__6406),
            .I(N__6395));
    Sp12to4 I__1154 (
            .O(N__6403),
            .I(N__6395));
    Odrv12 I__1153 (
            .O(N__6400),
            .I(A_c_22));
    Odrv12 I__1152 (
            .O(N__6395),
            .I(A_c_22));
    InMux I__1151 (
            .O(N__6390),
            .I(N__6387));
    LocalMux I__1150 (
            .O(N__6387),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3 ));
    InMux I__1149 (
            .O(N__6384),
            .I(N__6376));
    InMux I__1148 (
            .O(N__6383),
            .I(N__6373));
    CascadeMux I__1147 (
            .O(N__6382),
            .I(N__6368));
    InMux I__1146 (
            .O(N__6381),
            .I(N__6363));
    InMux I__1145 (
            .O(N__6380),
            .I(N__6363));
    CascadeMux I__1144 (
            .O(N__6379),
            .I(N__6354));
    LocalMux I__1143 (
            .O(N__6376),
            .I(N__6346));
    LocalMux I__1142 (
            .O(N__6373),
            .I(N__6346));
    InMux I__1141 (
            .O(N__6372),
            .I(N__6343));
    InMux I__1140 (
            .O(N__6371),
            .I(N__6336));
    InMux I__1139 (
            .O(N__6368),
            .I(N__6336));
    LocalMux I__1138 (
            .O(N__6363),
            .I(N__6333));
    InMux I__1137 (
            .O(N__6362),
            .I(N__6326));
    InMux I__1136 (
            .O(N__6361),
            .I(N__6326));
    InMux I__1135 (
            .O(N__6360),
            .I(N__6326));
    InMux I__1134 (
            .O(N__6359),
            .I(N__6321));
    InMux I__1133 (
            .O(N__6358),
            .I(N__6321));
    InMux I__1132 (
            .O(N__6357),
            .I(N__6314));
    InMux I__1131 (
            .O(N__6354),
            .I(N__6314));
    InMux I__1130 (
            .O(N__6353),
            .I(N__6314));
    InMux I__1129 (
            .O(N__6352),
            .I(N__6311));
    InMux I__1128 (
            .O(N__6351),
            .I(N__6308));
    Span4Mux_h I__1127 (
            .O(N__6346),
            .I(N__6303));
    LocalMux I__1126 (
            .O(N__6343),
            .I(N__6303));
    InMux I__1125 (
            .O(N__6342),
            .I(N__6300));
    InMux I__1124 (
            .O(N__6341),
            .I(N__6297));
    LocalMux I__1123 (
            .O(N__6336),
            .I(N__6294));
    Span4Mux_v I__1122 (
            .O(N__6333),
            .I(N__6291));
    LocalMux I__1121 (
            .O(N__6326),
            .I(N__6286));
    LocalMux I__1120 (
            .O(N__6321),
            .I(N__6286));
    LocalMux I__1119 (
            .O(N__6314),
            .I(N__6279));
    LocalMux I__1118 (
            .O(N__6311),
            .I(N__6279));
    LocalMux I__1117 (
            .O(N__6308),
            .I(N__6279));
    Span4Mux_h I__1116 (
            .O(N__6303),
            .I(N__6272));
    LocalMux I__1115 (
            .O(N__6300),
            .I(N__6272));
    LocalMux I__1114 (
            .O(N__6297),
            .I(N__6272));
    Span4Mux_v I__1113 (
            .O(N__6294),
            .I(N__6269));
    Span4Mux_h I__1112 (
            .O(N__6291),
            .I(N__6262));
    Span4Mux_v I__1111 (
            .O(N__6286),
            .I(N__6262));
    Span4Mux_v I__1110 (
            .O(N__6279),
            .I(N__6262));
    Span4Mux_v I__1109 (
            .O(N__6272),
            .I(N__6259));
    Span4Mux_v I__1108 (
            .O(N__6269),
            .I(N__6256));
    Span4Mux_v I__1107 (
            .O(N__6262),
            .I(N__6253));
    Span4Mux_h I__1106 (
            .O(N__6259),
            .I(N__6250));
    Sp12to4 I__1105 (
            .O(N__6256),
            .I(N__6245));
    Sp12to4 I__1104 (
            .O(N__6253),
            .I(N__6245));
    Sp12to4 I__1103 (
            .O(N__6250),
            .I(N__6242));
    Span12Mux_h I__1102 (
            .O(N__6245),
            .I(N__6239));
    Span12Mux_v I__1101 (
            .O(N__6242),
            .I(N__6236));
    Odrv12 I__1100 (
            .O(N__6239),
            .I(A_c_1));
    Odrv12 I__1099 (
            .O(N__6236),
            .I(A_c_1));
    CascadeMux I__1098 (
            .O(N__6231),
            .I(N__6227));
    CascadeMux I__1097 (
            .O(N__6230),
            .I(N__6223));
    InMux I__1096 (
            .O(N__6227),
            .I(N__6220));
    CascadeMux I__1095 (
            .O(N__6226),
            .I(N__6217));
    InMux I__1094 (
            .O(N__6223),
            .I(N__6207));
    LocalMux I__1093 (
            .O(N__6220),
            .I(N__6204));
    InMux I__1092 (
            .O(N__6217),
            .I(N__6201));
    InMux I__1091 (
            .O(N__6216),
            .I(N__6196));
    InMux I__1090 (
            .O(N__6215),
            .I(N__6196));
    InMux I__1089 (
            .O(N__6214),
            .I(N__6191));
    InMux I__1088 (
            .O(N__6213),
            .I(N__6191));
    InMux I__1087 (
            .O(N__6212),
            .I(N__6184));
    InMux I__1086 (
            .O(N__6211),
            .I(N__6184));
    InMux I__1085 (
            .O(N__6210),
            .I(N__6184));
    LocalMux I__1084 (
            .O(N__6207),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    Odrv4 I__1083 (
            .O(N__6204),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    LocalMux I__1082 (
            .O(N__6201),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    LocalMux I__1081 (
            .O(N__6196),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    LocalMux I__1080 (
            .O(N__6191),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    LocalMux I__1079 (
            .O(N__6184),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    InMux I__1078 (
            .O(N__6171),
            .I(N__6168));
    LocalMux I__1077 (
            .O(N__6168),
            .I(N__6160));
    InMux I__1076 (
            .O(N__6167),
            .I(N__6155));
    InMux I__1075 (
            .O(N__6166),
            .I(N__6155));
    InMux I__1074 (
            .O(N__6165),
            .I(N__6150));
    InMux I__1073 (
            .O(N__6164),
            .I(N__6150));
    InMux I__1072 (
            .O(N__6163),
            .I(N__6147));
    Span4Mux_v I__1071 (
            .O(N__6160),
            .I(N__6140));
    LocalMux I__1070 (
            .O(N__6155),
            .I(N__6140));
    LocalMux I__1069 (
            .O(N__6150),
            .I(N__6140));
    LocalMux I__1068 (
            .O(N__6147),
            .I(\U409_AUTOCONFIG.N_122 ));
    Odrv4 I__1067 (
            .O(N__6140),
            .I(\U409_AUTOCONFIG.N_122 ));
    InMux I__1066 (
            .O(N__6135),
            .I(N__6128));
    InMux I__1065 (
            .O(N__6134),
            .I(N__6125));
    InMux I__1064 (
            .O(N__6133),
            .I(N__6122));
    InMux I__1063 (
            .O(N__6132),
            .I(N__6119));
    InMux I__1062 (
            .O(N__6131),
            .I(N__6116));
    LocalMux I__1061 (
            .O(N__6128),
            .I(N__6111));
    LocalMux I__1060 (
            .O(N__6125),
            .I(N__6106));
    LocalMux I__1059 (
            .O(N__6122),
            .I(N__6106));
    LocalMux I__1058 (
            .O(N__6119),
            .I(N__6101));
    LocalMux I__1057 (
            .O(N__6116),
            .I(N__6101));
    InMux I__1056 (
            .O(N__6115),
            .I(N__6098));
    InMux I__1055 (
            .O(N__6114),
            .I(N__6095));
    Span4Mux_h I__1054 (
            .O(N__6111),
            .I(N__6090));
    Span4Mux_v I__1053 (
            .O(N__6106),
            .I(N__6090));
    Span4Mux_h I__1052 (
            .O(N__6101),
            .I(N__6083));
    LocalMux I__1051 (
            .O(N__6098),
            .I(N__6083));
    LocalMux I__1050 (
            .O(N__6095),
            .I(N__6083));
    Span4Mux_v I__1049 (
            .O(N__6090),
            .I(N__6080));
    Span4Mux_v I__1048 (
            .O(N__6083),
            .I(N__6077));
    Sp12to4 I__1047 (
            .O(N__6080),
            .I(N__6072));
    Sp12to4 I__1046 (
            .O(N__6077),
            .I(N__6072));
    Span12Mux_h I__1045 (
            .O(N__6072),
            .I(N__6069));
    Span12Mux_v I__1044 (
            .O(N__6069),
            .I(N__6066));
    Odrv12 I__1043 (
            .O(N__6066),
            .I(A_c_19));
    InMux I__1042 (
            .O(N__6063),
            .I(N__6059));
    InMux I__1041 (
            .O(N__6062),
            .I(N__6056));
    LocalMux I__1040 (
            .O(N__6059),
            .I(ATA_BASE_3));
    LocalMux I__1039 (
            .O(N__6056),
            .I(ATA_BASE_3));
    CascadeMux I__1038 (
            .O(N__6051),
            .I(N__6048));
    InMux I__1037 (
            .O(N__6048),
            .I(N__6042));
    InMux I__1036 (
            .O(N__6047),
            .I(N__6039));
    InMux I__1035 (
            .O(N__6046),
            .I(N__6036));
    InMux I__1034 (
            .O(N__6045),
            .I(N__6033));
    LocalMux I__1033 (
            .O(N__6042),
            .I(N__6029));
    LocalMux I__1032 (
            .O(N__6039),
            .I(N__6022));
    LocalMux I__1031 (
            .O(N__6036),
            .I(N__6022));
    LocalMux I__1030 (
            .O(N__6033),
            .I(N__6022));
    CascadeMux I__1029 (
            .O(N__6032),
            .I(N__6019));
    Span4Mux_v I__1028 (
            .O(N__6029),
            .I(N__6016));
    Span4Mux_v I__1027 (
            .O(N__6022),
            .I(N__6013));
    InMux I__1026 (
            .O(N__6019),
            .I(N__6010));
    Sp12to4 I__1025 (
            .O(N__6016),
            .I(N__6003));
    Sp12to4 I__1024 (
            .O(N__6013),
            .I(N__6003));
    LocalMux I__1023 (
            .O(N__6010),
            .I(N__6003));
    Span12Mux_h I__1022 (
            .O(N__6003),
            .I(N__6000));
    Span12Mux_v I__1021 (
            .O(N__6000),
            .I(N__5997));
    Odrv12 I__1020 (
            .O(N__5997),
            .I(A_c_18));
    InMux I__1019 (
            .O(N__5994),
            .I(N__5991));
    LocalMux I__1018 (
            .O(N__5991),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2 ));
    InMux I__1017 (
            .O(N__5988),
            .I(N__5985));
    LocalMux I__1016 (
            .O(N__5985),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1 ));
    CascadeMux I__1015 (
            .O(N__5982),
            .I(N__5977));
    InMux I__1014 (
            .O(N__5981),
            .I(N__5974));
    InMux I__1013 (
            .O(N__5980),
            .I(N__5971));
    InMux I__1012 (
            .O(N__5977),
            .I(N__5968));
    LocalMux I__1011 (
            .O(N__5974),
            .I(N__5965));
    LocalMux I__1010 (
            .O(N__5971),
            .I(N__5962));
    LocalMux I__1009 (
            .O(N__5968),
            .I(N__5959));
    Span4Mux_v I__1008 (
            .O(N__5965),
            .I(N__5956));
    Span4Mux_h I__1007 (
            .O(N__5962),
            .I(N__5953));
    Span12Mux_v I__1006 (
            .O(N__5959),
            .I(N__5950));
    Sp12to4 I__1005 (
            .O(N__5956),
            .I(N__5947));
    Span4Mux_v I__1004 (
            .O(N__5953),
            .I(N__5944));
    Odrv12 I__1003 (
            .O(N__5950),
            .I(A_c_31));
    Odrv12 I__1002 (
            .O(N__5947),
            .I(A_c_31));
    Odrv4 I__1001 (
            .O(N__5944),
            .I(A_c_31));
    InMux I__1000 (
            .O(N__5937),
            .I(N__5934));
    LocalMux I__999 (
            .O(N__5934),
            .I(N_120));
    CascadeMux I__998 (
            .O(N__5931),
            .I(\U409_ADDRESS_DECODE.PORTSIZEZ0Z_0_cascade_ ));
    IoInMux I__997 (
            .O(N__5928),
            .I(N__5925));
    LocalMux I__996 (
            .O(N__5925),
            .I(N__5922));
    Span4Mux_s2_v I__995 (
            .O(N__5922),
            .I(N__5919));
    Span4Mux_h I__994 (
            .O(N__5919),
            .I(N__5916));
    Span4Mux_v I__993 (
            .O(N__5916),
            .I(N__5913));
    Span4Mux_v I__992 (
            .O(N__5913),
            .I(N__5910));
    Odrv4 I__991 (
            .O(N__5910),
            .I(PORTSIZE_0_i));
    InMux I__990 (
            .O(N__5907),
            .I(N__5904));
    LocalMux I__989 (
            .O(N__5904),
            .I(N__5899));
    CascadeMux I__988 (
            .O(N__5903),
            .I(N__5896));
    InMux I__987 (
            .O(N__5902),
            .I(N__5893));
    Span4Mux_v I__986 (
            .O(N__5899),
            .I(N__5890));
    InMux I__985 (
            .O(N__5896),
            .I(N__5887));
    LocalMux I__984 (
            .O(N__5893),
            .I(N__5884));
    Span4Mux_h I__983 (
            .O(N__5890),
            .I(N__5879));
    LocalMux I__982 (
            .O(N__5887),
            .I(N__5879));
    Span4Mux_v I__981 (
            .O(N__5884),
            .I(N__5876));
    Span4Mux_h I__980 (
            .O(N__5879),
            .I(N__5873));
    Sp12to4 I__979 (
            .O(N__5876),
            .I(N__5870));
    Span4Mux_v I__978 (
            .O(N__5873),
            .I(N__5867));
    Odrv12 I__977 (
            .O(N__5870),
            .I(A_c_30));
    Odrv4 I__976 (
            .O(N__5867),
            .I(A_c_30));
    CascadeMux I__975 (
            .O(N__5862),
            .I(N__5859));
    InMux I__974 (
            .O(N__5859),
            .I(N__5856));
    LocalMux I__973 (
            .O(N__5856),
            .I(N__5853));
    Span4Mux_h I__972 (
            .O(N__5853),
            .I(N__5849));
    InMux I__971 (
            .O(N__5852),
            .I(N__5846));
    Span4Mux_h I__970 (
            .O(N__5849),
            .I(N__5840));
    LocalMux I__969 (
            .O(N__5846),
            .I(N__5840));
    InMux I__968 (
            .O(N__5845),
            .I(N__5837));
    Span4Mux_v I__967 (
            .O(N__5840),
            .I(N__5834));
    LocalMux I__966 (
            .O(N__5837),
            .I(N__5831));
    Span4Mux_v I__965 (
            .O(N__5834),
            .I(N__5828));
    Span12Mux_v I__964 (
            .O(N__5831),
            .I(N__5823));
    Sp12to4 I__963 (
            .O(N__5828),
            .I(N__5823));
    Odrv12 I__962 (
            .O(N__5823),
            .I(A_c_29));
    InMux I__961 (
            .O(N__5820),
            .I(N__5817));
    LocalMux I__960 (
            .O(N__5817),
            .I(\U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_0 ));
    IoInMux I__959 (
            .O(N__5814),
            .I(N__5811));
    LocalMux I__958 (
            .O(N__5811),
            .I(N__5808));
    Span12Mux_s10_v I__957 (
            .O(N__5808),
            .I(N__5805));
    Span12Mux_h I__956 (
            .O(N__5805),
            .I(N__5801));
    InMux I__955 (
            .O(N__5804),
            .I(N__5798));
    Odrv12 I__954 (
            .O(N__5801),
            .I(CONFIGENn_c));
    LocalMux I__953 (
            .O(N__5798),
            .I(CONFIGENn_c));
    InMux I__952 (
            .O(N__5793),
            .I(N__5786));
    InMux I__951 (
            .O(N__5792),
            .I(N__5777));
    InMux I__950 (
            .O(N__5791),
            .I(N__5777));
    InMux I__949 (
            .O(N__5790),
            .I(N__5777));
    InMux I__948 (
            .O(N__5789),
            .I(N__5777));
    LocalMux I__947 (
            .O(N__5786),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    LocalMux I__946 (
            .O(N__5777),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    InMux I__945 (
            .O(N__5772),
            .I(N__5765));
    InMux I__944 (
            .O(N__5771),
            .I(N__5756));
    InMux I__943 (
            .O(N__5770),
            .I(N__5756));
    InMux I__942 (
            .O(N__5769),
            .I(N__5756));
    InMux I__941 (
            .O(N__5768),
            .I(N__5756));
    LocalMux I__940 (
            .O(N__5765),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    LocalMux I__939 (
            .O(N__5756),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    InMux I__938 (
            .O(N__5751),
            .I(N__5746));
    InMux I__937 (
            .O(N__5750),
            .I(N__5741));
    InMux I__936 (
            .O(N__5749),
            .I(N__5741));
    LocalMux I__935 (
            .O(N__5746),
            .I(N__5738));
    LocalMux I__934 (
            .O(N__5741),
            .I(N__5735));
    Span4Mux_v I__933 (
            .O(N__5738),
            .I(N__5729));
    Span4Mux_v I__932 (
            .O(N__5735),
            .I(N__5729));
    InMux I__931 (
            .O(N__5734),
            .I(N__5726));
    Sp12to4 I__930 (
            .O(N__5729),
            .I(N__5721));
    LocalMux I__929 (
            .O(N__5726),
            .I(N__5721));
    Span12Mux_h I__928 (
            .O(N__5721),
            .I(N__5718));
    Span12Mux_v I__927 (
            .O(N__5718),
            .I(N__5715));
    Odrv12 I__926 (
            .O(N__5715),
            .I(TM_c_0));
    InMux I__925 (
            .O(N__5712),
            .I(N__5707));
    CascadeMux I__924 (
            .O(N__5711),
            .I(N__5700));
    InMux I__923 (
            .O(N__5710),
            .I(N__5697));
    LocalMux I__922 (
            .O(N__5707),
            .I(N__5694));
    InMux I__921 (
            .O(N__5706),
            .I(N__5689));
    InMux I__920 (
            .O(N__5705),
            .I(N__5689));
    InMux I__919 (
            .O(N__5704),
            .I(N__5686));
    InMux I__918 (
            .O(N__5703),
            .I(N__5683));
    InMux I__917 (
            .O(N__5700),
            .I(N__5680));
    LocalMux I__916 (
            .O(N__5697),
            .I(CONFIGURED));
    Odrv4 I__915 (
            .O(N__5694),
            .I(CONFIGURED));
    LocalMux I__914 (
            .O(N__5689),
            .I(CONFIGURED));
    LocalMux I__913 (
            .O(N__5686),
            .I(CONFIGURED));
    LocalMux I__912 (
            .O(N__5683),
            .I(CONFIGURED));
    LocalMux I__911 (
            .O(N__5680),
            .I(CONFIGURED));
    InMux I__910 (
            .O(N__5667),
            .I(N__5660));
    InMux I__909 (
            .O(N__5666),
            .I(N__5660));
    CascadeMux I__908 (
            .O(N__5665),
            .I(N__5657));
    LocalMux I__907 (
            .O(N__5660),
            .I(N__5653));
    InMux I__906 (
            .O(N__5657),
            .I(N__5650));
    InMux I__905 (
            .O(N__5656),
            .I(N__5647));
    Span4Mux_v I__904 (
            .O(N__5653),
            .I(N__5642));
    LocalMux I__903 (
            .O(N__5650),
            .I(N__5642));
    LocalMux I__902 (
            .O(N__5647),
            .I(N__5639));
    Span4Mux_h I__901 (
            .O(N__5642),
            .I(N__5636));
    Span12Mux_h I__900 (
            .O(N__5639),
            .I(N__5631));
    Sp12to4 I__899 (
            .O(N__5636),
            .I(N__5631));
    Span12Mux_v I__898 (
            .O(N__5631),
            .I(N__5628));
    Odrv12 I__897 (
            .O(N__5628),
            .I(TM_c_1));
    InMux I__896 (
            .O(N__5625),
            .I(N__5621));
    InMux I__895 (
            .O(N__5624),
            .I(N__5618));
    LocalMux I__894 (
            .O(N__5621),
            .I(N__5614));
    LocalMux I__893 (
            .O(N__5618),
            .I(N__5611));
    InMux I__892 (
            .O(N__5617),
            .I(N__5607));
    Span4Mux_v I__891 (
            .O(N__5614),
            .I(N__5604));
    Span4Mux_v I__890 (
            .O(N__5611),
            .I(N__5601));
    InMux I__889 (
            .O(N__5610),
            .I(N__5598));
    LocalMux I__888 (
            .O(N__5607),
            .I(N__5595));
    Sp12to4 I__887 (
            .O(N__5604),
            .I(N__5588));
    Sp12to4 I__886 (
            .O(N__5601),
            .I(N__5588));
    LocalMux I__885 (
            .O(N__5598),
            .I(N__5588));
    Span12Mux_v I__884 (
            .O(N__5595),
            .I(N__5585));
    Span12Mux_h I__883 (
            .O(N__5588),
            .I(N__5582));
    Span12Mux_v I__882 (
            .O(N__5585),
            .I(N__5579));
    Span12Mux_v I__881 (
            .O(N__5582),
            .I(N__5576));
    Odrv12 I__880 (
            .O(N__5579),
            .I(A_c_17));
    Odrv12 I__879 (
            .O(N__5576),
            .I(A_c_17));
    CascadeMux I__878 (
            .O(N__5571),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1_cascade_ ));
    InMux I__877 (
            .O(N__5568),
            .I(N__5564));
    InMux I__876 (
            .O(N__5567),
            .I(N__5561));
    LocalMux I__875 (
            .O(N__5564),
            .I(ATA_BASE_1));
    LocalMux I__874 (
            .O(N__5561),
            .I(ATA_BASE_1));
    CascadeMux I__873 (
            .O(N__5556),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_4_cascade_ ));
    CascadeMux I__872 (
            .O(N__5553),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_ ));
    CascadeMux I__871 (
            .O(N__5550),
            .I(N__5546));
    CascadeMux I__870 (
            .O(N__5549),
            .I(N__5540));
    InMux I__869 (
            .O(N__5546),
            .I(N__5536));
    InMux I__868 (
            .O(N__5545),
            .I(N__5531));
    InMux I__867 (
            .O(N__5544),
            .I(N__5531));
    InMux I__866 (
            .O(N__5543),
            .I(N__5526));
    InMux I__865 (
            .O(N__5540),
            .I(N__5526));
    InMux I__864 (
            .O(N__5539),
            .I(N__5523));
    LocalMux I__863 (
            .O(N__5536),
            .I(N__5520));
    LocalMux I__862 (
            .O(N__5531),
            .I(N__5517));
    LocalMux I__861 (
            .O(N__5526),
            .I(N__5512));
    LocalMux I__860 (
            .O(N__5523),
            .I(N__5512));
    Span4Mux_v I__859 (
            .O(N__5520),
            .I(N__5507));
    Span4Mux_v I__858 (
            .O(N__5517),
            .I(N__5507));
    Span4Mux_v I__857 (
            .O(N__5512),
            .I(N__5504));
    Sp12to4 I__856 (
            .O(N__5507),
            .I(N__5499));
    Sp12to4 I__855 (
            .O(N__5504),
            .I(N__5499));
    Span12Mux_h I__854 (
            .O(N__5499),
            .I(N__5496));
    Span12Mux_v I__853 (
            .O(N__5496),
            .I(N__5493));
    Odrv12 I__852 (
            .O(N__5493),
            .I(RnW_c));
    InMux I__851 (
            .O(N__5490),
            .I(N__5487));
    LocalMux I__850 (
            .O(N__5487),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2Z0Z_4 ));
    CascadeMux I__849 (
            .O(N__5484),
            .I(N__5481));
    InMux I__848 (
            .O(N__5481),
            .I(N__5473));
    InMux I__847 (
            .O(N__5480),
            .I(N__5473));
    CascadeMux I__846 (
            .O(N__5479),
            .I(N__5467));
    CascadeMux I__845 (
            .O(N__5478),
            .I(N__5464));
    LocalMux I__844 (
            .O(N__5473),
            .I(N__5461));
    InMux I__843 (
            .O(N__5472),
            .I(N__5456));
    InMux I__842 (
            .O(N__5471),
            .I(N__5456));
    InMux I__841 (
            .O(N__5470),
            .I(N__5451));
    InMux I__840 (
            .O(N__5467),
            .I(N__5451));
    InMux I__839 (
            .O(N__5464),
            .I(N__5448));
    Span4Mux_v I__838 (
            .O(N__5461),
            .I(N__5445));
    LocalMux I__837 (
            .O(N__5456),
            .I(N__5438));
    LocalMux I__836 (
            .O(N__5451),
            .I(N__5438));
    LocalMux I__835 (
            .O(N__5448),
            .I(N__5438));
    Span4Mux_h I__834 (
            .O(N__5445),
            .I(N__5435));
    Span4Mux_v I__833 (
            .O(N__5438),
            .I(N__5432));
    Odrv4 I__832 (
            .O(N__5435),
            .I(\U409_ADDRESS_DECODE.Z2_SPACE ));
    Odrv4 I__831 (
            .O(N__5432),
            .I(\U409_ADDRESS_DECODE.Z2_SPACE ));
    IoInMux I__830 (
            .O(N__5427),
            .I(N__5424));
    LocalMux I__829 (
            .O(N__5424),
            .I(N__5421));
    IoSpan4Mux I__828 (
            .O(N__5421),
            .I(N__5418));
    Span4Mux_s1_h I__827 (
            .O(N__5418),
            .I(N__5415));
    Sp12to4 I__826 (
            .O(N__5415),
            .I(N__5412));
    Span12Mux_s6_h I__825 (
            .O(N__5412),
            .I(N__5409));
    Span12Mux_h I__824 (
            .O(N__5409),
            .I(N__5406));
    Span12Mux_v I__823 (
            .O(N__5406),
            .I(N__5403));
    Odrv12 I__822 (
            .O(N__5403),
            .I(N_120_i));
    IoInMux I__821 (
            .O(N__5400),
            .I(N__5397));
    LocalMux I__820 (
            .O(N__5397),
            .I(N__5394));
    IoSpan4Mux I__819 (
            .O(N__5394),
            .I(N__5391));
    Span4Mux_s3_v I__818 (
            .O(N__5391),
            .I(N__5388));
    Span4Mux_h I__817 (
            .O(N__5388),
            .I(N__5385));
    Sp12to4 I__816 (
            .O(N__5385),
            .I(N__5382));
    Span12Mux_v I__815 (
            .O(N__5382),
            .I(N__5379));
    Odrv12 I__814 (
            .O(N__5379),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn_i));
    InMux I__813 (
            .O(N__5376),
            .I(N__5370));
    InMux I__812 (
            .O(N__5375),
            .I(N__5370));
    LocalMux I__811 (
            .O(N__5370),
            .I(N__5367));
    Odrv4 I__810 (
            .O(N__5367),
            .I(\U409_ADDRESS_DECODE.N_102 ));
    InMux I__809 (
            .O(N__5364),
            .I(N__5358));
    InMux I__808 (
            .O(N__5363),
            .I(N__5358));
    LocalMux I__807 (
            .O(N__5358),
            .I(N__5355));
    Odrv4 I__806 (
            .O(N__5355),
            .I(\U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3Z0Z_0 ));
    InMux I__805 (
            .O(N__5352),
            .I(N__5349));
    LocalMux I__804 (
            .O(N__5349),
            .I(N__5346));
    Span4Mux_v I__803 (
            .O(N__5346),
            .I(N__5342));
    InMux I__802 (
            .O(N__5345),
            .I(N__5339));
    Odrv4 I__801 (
            .O(N__5342),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ));
    LocalMux I__800 (
            .O(N__5339),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ));
    InMux I__799 (
            .O(N__5334),
            .I(N__5330));
    CascadeMux I__798 (
            .O(N__5333),
            .I(N__5327));
    LocalMux I__797 (
            .O(N__5330),
            .I(N__5324));
    InMux I__796 (
            .O(N__5327),
            .I(N__5321));
    Odrv4 I__795 (
            .O(N__5324),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ));
    LocalMux I__794 (
            .O(N__5321),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ));
    IoInMux I__793 (
            .O(N__5316),
            .I(N__5313));
    LocalMux I__792 (
            .O(N__5313),
            .I(N__5310));
    Span12Mux_s5_v I__791 (
            .O(N__5310),
            .I(N__5307));
    Odrv12 I__790 (
            .O(N__5307),
            .I(U409_AUTOCONFIG_D_OUT_0_i_1));
    InMux I__789 (
            .O(N__5304),
            .I(N__5300));
    InMux I__788 (
            .O(N__5303),
            .I(N__5297));
    LocalMux I__787 (
            .O(N__5300),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2 ));
    LocalMux I__786 (
            .O(N__5297),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2 ));
    CascadeMux I__785 (
            .O(N__5292),
            .I(N__5289));
    InMux I__784 (
            .O(N__5289),
            .I(N__5286));
    LocalMux I__783 (
            .O(N__5286),
            .I(N__5282));
    CascadeMux I__782 (
            .O(N__5285),
            .I(N__5279));
    Span4Mux_v I__781 (
            .O(N__5282),
            .I(N__5276));
    InMux I__780 (
            .O(N__5279),
            .I(N__5273));
    Odrv4 I__779 (
            .O(N__5276),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ));
    LocalMux I__778 (
            .O(N__5273),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ));
    IoInMux I__777 (
            .O(N__5268),
            .I(N__5265));
    LocalMux I__776 (
            .O(N__5265),
            .I(N__5262));
    Span12Mux_s10_v I__775 (
            .O(N__5262),
            .I(N__5259));
    Odrv12 I__774 (
            .O(N__5259),
            .I(U409_AUTOCONFIG_D_OUT_0_i_2));
    InMux I__773 (
            .O(N__5256),
            .I(N__5252));
    InMux I__772 (
            .O(N__5255),
            .I(N__5249));
    LocalMux I__771 (
            .O(N__5252),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ));
    LocalMux I__770 (
            .O(N__5249),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ));
    CascadeMux I__769 (
            .O(N__5244),
            .I(N__5241));
    InMux I__768 (
            .O(N__5241),
            .I(N__5238));
    LocalMux I__767 (
            .O(N__5238),
            .I(N__5235));
    Span4Mux_v I__766 (
            .O(N__5235),
            .I(N__5231));
    InMux I__765 (
            .O(N__5234),
            .I(N__5228));
    Odrv4 I__764 (
            .O(N__5231),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ));
    LocalMux I__763 (
            .O(N__5228),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ));
    IoInMux I__762 (
            .O(N__5223),
            .I(N__5220));
    LocalMux I__761 (
            .O(N__5220),
            .I(N__5217));
    Span4Mux_s2_v I__760 (
            .O(N__5217),
            .I(N__5214));
    Sp12to4 I__759 (
            .O(N__5214),
            .I(N__5211));
    Span12Mux_h I__758 (
            .O(N__5211),
            .I(N__5208));
    Span12Mux_v I__757 (
            .O(N__5208),
            .I(N__5205));
    Odrv12 I__756 (
            .O(N__5205),
            .I(U409_AUTOCONFIG_D_OUT_0_i_3));
    InMux I__755 (
            .O(N__5202),
            .I(N__5199));
    LocalMux I__754 (
            .O(N__5199),
            .I(N__5196));
    Odrv12 I__753 (
            .O(N__5196),
            .I(\U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0Z0Z_0 ));
    CascadeMux I__752 (
            .O(N__5193),
            .I(N__5189));
    CascadeMux I__751 (
            .O(N__5192),
            .I(N__5185));
    InMux I__750 (
            .O(N__5189),
            .I(N__5175));
    InMux I__749 (
            .O(N__5188),
            .I(N__5175));
    InMux I__748 (
            .O(N__5185),
            .I(N__5175));
    InMux I__747 (
            .O(N__5184),
            .I(N__5175));
    LocalMux I__746 (
            .O(N__5175),
            .I(\U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa ));
    InMux I__745 (
            .O(N__5172),
            .I(N__5169));
    LocalMux I__744 (
            .O(N__5169),
            .I(N__5166));
    Odrv4 I__743 (
            .O(N__5166),
            .I(\U409_ADDRESS_DECODE.HIROMZ0 ));
    CascadeMux I__742 (
            .O(N__5163),
            .I(\U409_ADDRESS_DECODE.LOWROMZ0Z_2_cascade_ ));
    IoInMux I__741 (
            .O(N__5160),
            .I(N__5157));
    LocalMux I__740 (
            .O(N__5157),
            .I(N__5152));
    IoInMux I__739 (
            .O(N__5156),
            .I(N__5149));
    IoInMux I__738 (
            .O(N__5155),
            .I(N__5146));
    IoSpan4Mux I__737 (
            .O(N__5152),
            .I(N__5139));
    LocalMux I__736 (
            .O(N__5149),
            .I(N__5139));
    LocalMux I__735 (
            .O(N__5146),
            .I(N__5139));
    IoSpan4Mux I__734 (
            .O(N__5139),
            .I(N__5136));
    Span4Mux_s2_v I__733 (
            .O(N__5136),
            .I(N__5132));
    IoInMux I__732 (
            .O(N__5135),
            .I(N__5129));
    Sp12to4 I__731 (
            .O(N__5132),
            .I(N__5124));
    LocalMux I__730 (
            .O(N__5129),
            .I(N__5124));
    Span12Mux_s10_v I__729 (
            .O(N__5124),
            .I(N__5121));
    Odrv12 I__728 (
            .O(N__5121),
            .I(D_1_i));
    InMux I__727 (
            .O(N__5118),
            .I(N__5115));
    LocalMux I__726 (
            .O(N__5115),
            .I(\U409_AUTOCONFIG.AC_STARTZ0 ));
    CascadeMux I__725 (
            .O(N__5112),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2Z0Z_1_cascade_ ));
    CascadeMux I__724 (
            .O(N__5109),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2Z0Z_4_cascade_ ));
    InMux I__723 (
            .O(N__5106),
            .I(N__5103));
    LocalMux I__722 (
            .O(N__5103),
            .I(N__5100));
    Odrv4 I__721 (
            .O(N__5100),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_10 ));
    CascadeMux I__720 (
            .O(N__5097),
            .I(N_120_cascade_));
    InMux I__719 (
            .O(N__5094),
            .I(N__5091));
    LocalMux I__718 (
            .O(N__5091),
            .I(N__5088));
    Span12Mux_h I__717 (
            .O(N__5088),
            .I(N__5085));
    Odrv12 I__716 (
            .O(N__5085),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_11 ));
    InMux I__715 (
            .O(N__5082),
            .I(N__5079));
    LocalMux I__714 (
            .O(N__5079),
            .I(N__5076));
    Span4Mux_h I__713 (
            .O(N__5076),
            .I(N__5073));
    Odrv4 I__712 (
            .O(N__5073),
            .I(\U409_AUTOCONFIG.N_31 ));
    InMux I__711 (
            .O(N__5070),
            .I(N__5067));
    LocalMux I__710 (
            .O(N__5067),
            .I(N__5064));
    Span4Mux_h I__709 (
            .O(N__5064),
            .I(N__5061));
    Odrv4 I__708 (
            .O(N__5061),
            .I(\U409_AUTOCONFIG.N_22 ));
    InMux I__707 (
            .O(N__5058),
            .I(N__5055));
    LocalMux I__706 (
            .O(N__5055),
            .I(N__5052));
    Odrv12 I__705 (
            .O(N__5052),
            .I(\U409_AUTOCONFIG.LIDE_CONF_1_sqmuxa_0_a2_0Z0Z_2 ));
    InMux I__704 (
            .O(N__5049),
            .I(N__5046));
    LocalMux I__703 (
            .O(N__5046),
            .I(N__5043));
    Odrv4 I__702 (
            .O(N__5043),
            .I(\U409_AUTOCONFIG.N_20 ));
    InMux I__701 (
            .O(N__5040),
            .I(N__5037));
    LocalMux I__700 (
            .O(N__5037),
            .I(N__5034));
    Span12Mux_v I__699 (
            .O(N__5034),
            .I(N__5031));
    Odrv12 I__698 (
            .O(N__5031),
            .I(CPUCONFn_c));
    InMux I__697 (
            .O(N__5028),
            .I(N__5025));
    LocalMux I__696 (
            .O(N__5025),
            .I(\U409_AUTOCONFIG.N_52 ));
    CascadeMux I__695 (
            .O(N__5022),
            .I(\U409_AUTOCONFIG.N_52_cascade_ ));
    InMux I__694 (
            .O(N__5019),
            .I(N__5011));
    InMux I__693 (
            .O(N__5018),
            .I(N__5011));
    InMux I__692 (
            .O(N__5017),
            .I(N__5006));
    InMux I__691 (
            .O(N__5016),
            .I(N__5006));
    LocalMux I__690 (
            .O(N__5011),
            .I(\U409_AUTOCONFIG.N_56 ));
    LocalMux I__689 (
            .O(N__5006),
            .I(\U409_AUTOCONFIG.N_56 ));
    CascadeMux I__688 (
            .O(N__5001),
            .I(N__4997));
    InMux I__687 (
            .O(N__5000),
            .I(N__4994));
    InMux I__686 (
            .O(N__4997),
            .I(N__4991));
    LocalMux I__685 (
            .O(N__4994),
            .I(N__4988));
    LocalMux I__684 (
            .O(N__4991),
            .I(N__4985));
    Odrv12 I__683 (
            .O(N__4988),
            .I(\U409_AUTOCONFIG.N_67 ));
    Odrv4 I__682 (
            .O(N__4985),
            .I(\U409_AUTOCONFIG.N_67 ));
    CascadeMux I__681 (
            .O(N__4980),
            .I(\U409_AUTOCONFIG.N_56_cascade_ ));
    CascadeMux I__680 (
            .O(N__4977),
            .I(N__4971));
    CascadeMux I__679 (
            .O(N__4976),
            .I(N__4968));
    CascadeMux I__678 (
            .O(N__4975),
            .I(N__4965));
    CascadeMux I__677 (
            .O(N__4974),
            .I(N__4961));
    InMux I__676 (
            .O(N__4971),
            .I(N__4955));
    InMux I__675 (
            .O(N__4968),
            .I(N__4950));
    InMux I__674 (
            .O(N__4965),
            .I(N__4950));
    InMux I__673 (
            .O(N__4964),
            .I(N__4942));
    InMux I__672 (
            .O(N__4961),
            .I(N__4942));
    InMux I__671 (
            .O(N__4960),
            .I(N__4939));
    InMux I__670 (
            .O(N__4959),
            .I(N__4934));
    InMux I__669 (
            .O(N__4958),
            .I(N__4934));
    LocalMux I__668 (
            .O(N__4955),
            .I(N__4929));
    LocalMux I__667 (
            .O(N__4950),
            .I(N__4929));
    InMux I__666 (
            .O(N__4949),
            .I(N__4926));
    InMux I__665 (
            .O(N__4948),
            .I(N__4921));
    InMux I__664 (
            .O(N__4947),
            .I(N__4921));
    LocalMux I__663 (
            .O(N__4942),
            .I(N__4918));
    LocalMux I__662 (
            .O(N__4939),
            .I(N__4913));
    LocalMux I__661 (
            .O(N__4934),
            .I(N__4913));
    Span4Mux_v I__660 (
            .O(N__4929),
            .I(N__4910));
    LocalMux I__659 (
            .O(N__4926),
            .I(N__4905));
    LocalMux I__658 (
            .O(N__4921),
            .I(N__4905));
    Span4Mux_v I__657 (
            .O(N__4918),
            .I(N__4901));
    Span4Mux_v I__656 (
            .O(N__4913),
            .I(N__4898));
    Span4Mux_h I__655 (
            .O(N__4910),
            .I(N__4893));
    Span4Mux_v I__654 (
            .O(N__4905),
            .I(N__4893));
    InMux I__653 (
            .O(N__4904),
            .I(N__4890));
    Sp12to4 I__652 (
            .O(N__4901),
            .I(N__4881));
    Sp12to4 I__651 (
            .O(N__4898),
            .I(N__4881));
    Sp12to4 I__650 (
            .O(N__4893),
            .I(N__4881));
    LocalMux I__649 (
            .O(N__4890),
            .I(N__4881));
    Odrv12 I__648 (
            .O(N__4881),
            .I(A_c_4));
    InMux I__647 (
            .O(N__4878),
            .I(N__4875));
    LocalMux I__646 (
            .O(N__4875),
            .I(N__4868));
    InMux I__645 (
            .O(N__4874),
            .I(N__4863));
    InMux I__644 (
            .O(N__4873),
            .I(N__4863));
    CascadeMux I__643 (
            .O(N__4872),
            .I(N__4859));
    CascadeMux I__642 (
            .O(N__4871),
            .I(N__4856));
    Span4Mux_v I__641 (
            .O(N__4868),
            .I(N__4853));
    LocalMux I__640 (
            .O(N__4863),
            .I(N__4848));
    CascadeMux I__639 (
            .O(N__4862),
            .I(N__4845));
    InMux I__638 (
            .O(N__4859),
            .I(N__4838));
    InMux I__637 (
            .O(N__4856),
            .I(N__4838));
    Span4Mux_h I__636 (
            .O(N__4853),
            .I(N__4835));
    InMux I__635 (
            .O(N__4852),
            .I(N__4830));
    InMux I__634 (
            .O(N__4851),
            .I(N__4830));
    Span4Mux_v I__633 (
            .O(N__4848),
            .I(N__4827));
    InMux I__632 (
            .O(N__4845),
            .I(N__4820));
    InMux I__631 (
            .O(N__4844),
            .I(N__4820));
    InMux I__630 (
            .O(N__4843),
            .I(N__4820));
    LocalMux I__629 (
            .O(N__4838),
            .I(N__4817));
    Sp12to4 I__628 (
            .O(N__4835),
            .I(N__4808));
    LocalMux I__627 (
            .O(N__4830),
            .I(N__4808));
    Sp12to4 I__626 (
            .O(N__4827),
            .I(N__4808));
    LocalMux I__625 (
            .O(N__4820),
            .I(N__4808));
    Span4Mux_v I__624 (
            .O(N__4817),
            .I(N__4805));
    Span12Mux_h I__623 (
            .O(N__4808),
            .I(N__4802));
    Span4Mux_h I__622 (
            .O(N__4805),
            .I(N__4799));
    Span12Mux_v I__621 (
            .O(N__4802),
            .I(N__4796));
    Sp12to4 I__620 (
            .O(N__4799),
            .I(N__4793));
    Odrv12 I__619 (
            .O(N__4796),
            .I(A_c_2));
    Odrv12 I__618 (
            .O(N__4793),
            .I(A_c_2));
    InMux I__617 (
            .O(N__4788),
            .I(N__4785));
    LocalMux I__616 (
            .O(N__4785),
            .I(\U409_AUTOCONFIG.N_44 ));
    InMux I__615 (
            .O(N__4782),
            .I(N__4779));
    LocalMux I__614 (
            .O(N__4779),
            .I(N__4775));
    InMux I__613 (
            .O(N__4778),
            .I(N__4772));
    Span4Mux_v I__612 (
            .O(N__4775),
            .I(N__4765));
    LocalMux I__611 (
            .O(N__4772),
            .I(N__4762));
    InMux I__610 (
            .O(N__4771),
            .I(N__4757));
    InMux I__609 (
            .O(N__4770),
            .I(N__4757));
    InMux I__608 (
            .O(N__4769),
            .I(N__4752));
    InMux I__607 (
            .O(N__4768),
            .I(N__4752));
    Odrv4 I__606 (
            .O(N__4765),
            .I(\U409_AUTOCONFIG.N_86 ));
    Odrv4 I__605 (
            .O(N__4762),
            .I(\U409_AUTOCONFIG.N_86 ));
    LocalMux I__604 (
            .O(N__4757),
            .I(\U409_AUTOCONFIG.N_86 ));
    LocalMux I__603 (
            .O(N__4752),
            .I(\U409_AUTOCONFIG.N_86 ));
    InMux I__602 (
            .O(N__4743),
            .I(N__4730));
    InMux I__601 (
            .O(N__4742),
            .I(N__4730));
    InMux I__600 (
            .O(N__4741),
            .I(N__4730));
    InMux I__599 (
            .O(N__4740),
            .I(N__4730));
    CascadeMux I__598 (
            .O(N__4739),
            .I(N__4727));
    LocalMux I__597 (
            .O(N__4730),
            .I(N__4720));
    InMux I__596 (
            .O(N__4727),
            .I(N__4717));
    InMux I__595 (
            .O(N__4726),
            .I(N__4712));
    InMux I__594 (
            .O(N__4725),
            .I(N__4712));
    InMux I__593 (
            .O(N__4724),
            .I(N__4709));
    InMux I__592 (
            .O(N__4723),
            .I(N__4706));
    Span4Mux_v I__591 (
            .O(N__4720),
            .I(N__4702));
    LocalMux I__590 (
            .O(N__4717),
            .I(N__4695));
    LocalMux I__589 (
            .O(N__4712),
            .I(N__4695));
    LocalMux I__588 (
            .O(N__4709),
            .I(N__4695));
    LocalMux I__587 (
            .O(N__4706),
            .I(N__4692));
    InMux I__586 (
            .O(N__4705),
            .I(N__4689));
    Span4Mux_h I__585 (
            .O(N__4702),
            .I(N__4684));
    Span4Mux_v I__584 (
            .O(N__4695),
            .I(N__4684));
    Span4Mux_h I__583 (
            .O(N__4692),
            .I(N__4679));
    LocalMux I__582 (
            .O(N__4689),
            .I(N__4679));
    Sp12to4 I__581 (
            .O(N__4684),
            .I(N__4676));
    Sp12to4 I__580 (
            .O(N__4679),
            .I(N__4673));
    Span12Mux_s5_h I__579 (
            .O(N__4676),
            .I(N__4670));
    Span12Mux_v I__578 (
            .O(N__4673),
            .I(N__4667));
    Span12Mux_v I__577 (
            .O(N__4670),
            .I(N__4664));
    Odrv12 I__576 (
            .O(N__4667),
            .I(A_c_3));
    Odrv12 I__575 (
            .O(N__4664),
            .I(A_c_3));
    InMux I__574 (
            .O(N__4659),
            .I(N__4656));
    LocalMux I__573 (
            .O(N__4656),
            .I(\U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_1_85_i_i_0 ));
    InMux I__572 (
            .O(N__4653),
            .I(N__4649));
    InMux I__571 (
            .O(N__4652),
            .I(N__4646));
    LocalMux I__570 (
            .O(N__4649),
            .I(N_121));
    LocalMux I__569 (
            .O(N__4646),
            .I(N_121));
    CascadeMux I__568 (
            .O(N__4641),
            .I(N_121_cascade_));
    IoInMux I__567 (
            .O(N__4638),
            .I(N__4635));
    LocalMux I__566 (
            .O(N__4635),
            .I(N__4631));
    InMux I__565 (
            .O(N__4634),
            .I(N__4627));
    IoSpan4Mux I__564 (
            .O(N__4631),
            .I(N__4623));
    InMux I__563 (
            .O(N__4630),
            .I(N__4620));
    LocalMux I__562 (
            .O(N__4627),
            .I(N__4617));
    InMux I__561 (
            .O(N__4626),
            .I(N__4614));
    Span4Mux_s0_h I__560 (
            .O(N__4623),
            .I(N__4611));
    LocalMux I__559 (
            .O(N__4620),
            .I(N__4608));
    Span4Mux_v I__558 (
            .O(N__4617),
            .I(N__4603));
    LocalMux I__557 (
            .O(N__4614),
            .I(N__4603));
    Sp12to4 I__556 (
            .O(N__4611),
            .I(N__4600));
    Span4Mux_v I__555 (
            .O(N__4608),
            .I(N__4597));
    Span4Mux_v I__554 (
            .O(N__4603),
            .I(N__4594));
    Span12Mux_v I__553 (
            .O(N__4600),
            .I(N__4591));
    Sp12to4 I__552 (
            .O(N__4597),
            .I(N__4588));
    Span4Mux_v I__551 (
            .O(N__4594),
            .I(N__4585));
    Span12Mux_h I__550 (
            .O(N__4591),
            .I(N__4582));
    Span12Mux_h I__549 (
            .O(N__4588),
            .I(N__4579));
    Span4Mux_v I__548 (
            .O(N__4585),
            .I(N__4576));
    Span12Mux_h I__547 (
            .O(N__4582),
            .I(N__4569));
    Span12Mux_v I__546 (
            .O(N__4579),
            .I(N__4569));
    Sp12to4 I__545 (
            .O(N__4576),
            .I(N__4569));
    Odrv12 I__544 (
            .O(N__4569),
            .I(A_c_16));
    InMux I__543 (
            .O(N__4566),
            .I(N__4563));
    LocalMux I__542 (
            .O(N__4563),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_1 ));
    InMux I__541 (
            .O(N__4560),
            .I(N__4557));
    LocalMux I__540 (
            .O(N__4557),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2 ));
    InMux I__539 (
            .O(N__4554),
            .I(N__4551));
    LocalMux I__538 (
            .O(N__4551),
            .I(N__4548));
    Span4Mux_v I__537 (
            .O(N__4548),
            .I(N__4545));
    Odrv4 I__536 (
            .O(N__4545),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_7 ));
    InMux I__535 (
            .O(N__4542),
            .I(N__4538));
    InMux I__534 (
            .O(N__4541),
            .I(N__4535));
    LocalMux I__533 (
            .O(N__4538),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_0 ));
    LocalMux I__532 (
            .O(N__4535),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_0 ));
    IoInMux I__531 (
            .O(N__4530),
            .I(N__4527));
    LocalMux I__530 (
            .O(N__4527),
            .I(N__4524));
    Span12Mux_s4_v I__529 (
            .O(N__4524),
            .I(N__4521));
    Odrv12 I__528 (
            .O(N__4521),
            .I(U409_AUTOCONFIG_D_OUT_0_i_0));
    InMux I__527 (
            .O(N__4518),
            .I(N__4515));
    LocalMux I__526 (
            .O(N__4515),
            .I(N__4512));
    Span4Mux_v I__525 (
            .O(N__4512),
            .I(N__4509));
    Odrv4 I__524 (
            .O(N__4509),
            .I(\U409_AUTOCONFIG.N_27 ));
    CascadeMux I__523 (
            .O(N__4506),
            .I(N__4502));
    InMux I__522 (
            .O(N__4505),
            .I(N__4497));
    InMux I__521 (
            .O(N__4502),
            .I(N__4497));
    LocalMux I__520 (
            .O(N__4497),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ));
    InMux I__519 (
            .O(N__4494),
            .I(N__4491));
    LocalMux I__518 (
            .O(N__4491),
            .I(N__4487));
    InMux I__517 (
            .O(N__4490),
            .I(N__4484));
    Odrv4 I__516 (
            .O(N__4487),
            .I(\U409_AUTOCONFIG.N_111 ));
    LocalMux I__515 (
            .O(N__4484),
            .I(\U409_AUTOCONFIG.N_111 ));
    InMux I__514 (
            .O(N__4479),
            .I(N__4474));
    InMux I__513 (
            .O(N__4478),
            .I(N__4471));
    InMux I__512 (
            .O(N__4477),
            .I(N__4468));
    LocalMux I__511 (
            .O(N__4474),
            .I(\U409_AUTOCONFIG.N_41 ));
    LocalMux I__510 (
            .O(N__4471),
            .I(\U409_AUTOCONFIG.N_41 ));
    LocalMux I__509 (
            .O(N__4468),
            .I(\U409_AUTOCONFIG.N_41 ));
    InMux I__508 (
            .O(N__4461),
            .I(N__4458));
    LocalMux I__507 (
            .O(N__4458),
            .I(\U409_AUTOCONFIG.N_43 ));
    InMux I__506 (
            .O(N__4455),
            .I(N__4452));
    LocalMux I__505 (
            .O(N__4452),
            .I(\U409_AUTOCONFIG.N_66 ));
    CascadeMux I__504 (
            .O(N__4449),
            .I(\U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_i_1_cascade_ ));
    InMux I__503 (
            .O(N__4446),
            .I(N__4443));
    LocalMux I__502 (
            .O(N__4443),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_4 ));
    CascadeMux I__501 (
            .O(N__4440),
            .I(\U409_ADDRESS_DECODE.N_112_cascade_ ));
    InMux I__500 (
            .O(N__4437),
            .I(N__4434));
    LocalMux I__499 (
            .O(N__4434),
            .I(\U409_ADDRESS_DECODE.N_112 ));
    CascadeMux I__498 (
            .O(N__4431),
            .I(\U409_AUTOCONFIG.N_74_cascade_ ));
    InMux I__497 (
            .O(N__4428),
            .I(N__4425));
    LocalMux I__496 (
            .O(N__4425),
            .I(\U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_i_0 ));
    InMux I__495 (
            .O(N__4422),
            .I(N__4419));
    LocalMux I__494 (
            .O(N__4419),
            .I(N__4416));
    Span4Mux_h I__493 (
            .O(N__4416),
            .I(N__4413));
    Odrv4 I__492 (
            .O(N__4413),
            .I(N_89_1));
    CascadeMux I__491 (
            .O(N__4410),
            .I(N_89_1_cascade_));
    InMux I__490 (
            .O(N__4407),
            .I(N__4404));
    LocalMux I__489 (
            .O(N__4404),
            .I(N__4401));
    Odrv4 I__488 (
            .O(N__4401),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_3 ));
    InMux I__487 (
            .O(N__4398),
            .I(N__4394));
    InMux I__486 (
            .O(N__4397),
            .I(N__4391));
    LocalMux I__485 (
            .O(N__4394),
            .I(N__4388));
    LocalMux I__484 (
            .O(N__4391),
            .I(N__4385));
    Span4Mux_v I__483 (
            .O(N__4388),
            .I(N__4382));
    Span4Mux_v I__482 (
            .O(N__4385),
            .I(N__4379));
    Sp12to4 I__481 (
            .O(N__4382),
            .I(N__4374));
    Sp12to4 I__480 (
            .O(N__4379),
            .I(N__4374));
    Odrv12 I__479 (
            .O(N__4374),
            .I(A_c_25));
    InMux I__478 (
            .O(N__4371),
            .I(N__4368));
    LocalMux I__477 (
            .O(N__4368),
            .I(N__4365));
    Span12Mux_h I__476 (
            .O(N__4365),
            .I(N__4362));
    Odrv12 I__475 (
            .O(N__4362),
            .I(TT_c_0));
    CascadeMux I__474 (
            .O(N__4359),
            .I(N__4356));
    InMux I__473 (
            .O(N__4356),
            .I(N__4353));
    LocalMux I__472 (
            .O(N__4353),
            .I(N__4350));
    Span4Mux_h I__471 (
            .O(N__4350),
            .I(N__4347));
    Sp12to4 I__470 (
            .O(N__4347),
            .I(N__4344));
    Odrv12 I__469 (
            .O(N__4344),
            .I(TT_c_1));
    CascadeMux I__468 (
            .O(N__4341),
            .I(N__4338));
    InMux I__467 (
            .O(N__4338),
            .I(N__4335));
    LocalMux I__466 (
            .O(N__4335),
            .I(N__4332));
    Odrv4 I__465 (
            .O(N__4332),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_9 ));
    InMux I__464 (
            .O(N__4329),
            .I(N__4323));
    InMux I__463 (
            .O(N__4328),
            .I(N__4323));
    LocalMux I__462 (
            .O(N__4323),
            .I(\U409_AUTOCONFIG.N_38 ));
    InMux I__461 (
            .O(N__4320),
            .I(N__4317));
    LocalMux I__460 (
            .O(N__4317),
            .I(\U409_AUTOCONFIG.N_48 ));
    CascadeMux I__459 (
            .O(N__4314),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_1_0_cascade_ ));
    InMux I__458 (
            .O(N__4311),
            .I(N__4305));
    InMux I__457 (
            .O(N__4310),
            .I(N__4305));
    LocalMux I__456 (
            .O(N__4305),
            .I(N__4302));
    Odrv4 I__455 (
            .O(N__4302),
            .I(\U409_AUTOCONFIG.N_62 ));
    CascadeMux I__454 (
            .O(N__4299),
            .I(\U409_ADDRESS_DECODE.N_54_cascade_ ));
    InMux I__453 (
            .O(N__4296),
            .I(N__4288));
    InMux I__452 (
            .O(N__4295),
            .I(N__4288));
    InMux I__451 (
            .O(N__4294),
            .I(N__4283));
    InMux I__450 (
            .O(N__4293),
            .I(N__4283));
    LocalMux I__449 (
            .O(N__4288),
            .I(N__4280));
    LocalMux I__448 (
            .O(N__4283),
            .I(N__4275));
    Span4Mux_v I__447 (
            .O(N__4280),
            .I(N__4272));
    InMux I__446 (
            .O(N__4279),
            .I(N__4269));
    InMux I__445 (
            .O(N__4278),
            .I(N__4266));
    Span4Mux_v I__444 (
            .O(N__4275),
            .I(N__4263));
    Sp12to4 I__443 (
            .O(N__4272),
            .I(N__4254));
    LocalMux I__442 (
            .O(N__4269),
            .I(N__4254));
    LocalMux I__441 (
            .O(N__4266),
            .I(N__4254));
    Sp12to4 I__440 (
            .O(N__4263),
            .I(N__4254));
    Odrv12 I__439 (
            .O(N__4254),
            .I(A_c_5));
    CascadeMux I__438 (
            .O(N__4251),
            .I(N__4247));
    InMux I__437 (
            .O(N__4250),
            .I(N__4242));
    InMux I__436 (
            .O(N__4247),
            .I(N__4242));
    LocalMux I__435 (
            .O(N__4242),
            .I(N__4238));
    InMux I__434 (
            .O(N__4241),
            .I(N__4235));
    Odrv4 I__433 (
            .O(N__4238),
            .I(\U409_AUTOCONFIG.N_92 ));
    LocalMux I__432 (
            .O(N__4235),
            .I(\U409_AUTOCONFIG.N_92 ));
    CascadeMux I__431 (
            .O(N__4230),
            .I(\U409_AUTOCONFIG.N_86_cascade_ ));
    InMux I__430 (
            .O(N__4227),
            .I(N__4224));
    LocalMux I__429 (
            .O(N__4224),
            .I(\U409_AUTOCONFIG.N_57 ));
    InMux I__428 (
            .O(N__4221),
            .I(N__4218));
    LocalMux I__427 (
            .O(N__4218),
            .I(N__4215));
    Span4Mux_v I__426 (
            .O(N__4215),
            .I(N__4209));
    InMux I__425 (
            .O(N__4214),
            .I(N__4202));
    InMux I__424 (
            .O(N__4213),
            .I(N__4202));
    InMux I__423 (
            .O(N__4212),
            .I(N__4202));
    Sp12to4 I__422 (
            .O(N__4209),
            .I(N__4197));
    LocalMux I__421 (
            .O(N__4202),
            .I(N__4197));
    Odrv12 I__420 (
            .O(N__4197),
            .I(A_c_7));
    InMux I__419 (
            .O(N__4194),
            .I(N__4185));
    InMux I__418 (
            .O(N__4193),
            .I(N__4185));
    InMux I__417 (
            .O(N__4192),
            .I(N__4185));
    LocalMux I__416 (
            .O(N__4185),
            .I(N__4181));
    CascadeMux I__415 (
            .O(N__4184),
            .I(N__4178));
    Span4Mux_v I__414 (
            .O(N__4181),
            .I(N__4175));
    InMux I__413 (
            .O(N__4178),
            .I(N__4172));
    Sp12to4 I__412 (
            .O(N__4175),
            .I(N__4167));
    LocalMux I__411 (
            .O(N__4172),
            .I(N__4167));
    Odrv12 I__410 (
            .O(N__4167),
            .I(A_c_6));
    CascadeMux I__409 (
            .O(N__4164),
            .I(\U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4_cascade_ ));
    CascadeMux I__408 (
            .O(N__4161),
            .I(N__4157));
    InMux I__407 (
            .O(N__4160),
            .I(N__4154));
    InMux I__406 (
            .O(N__4157),
            .I(N__4151));
    LocalMux I__405 (
            .O(N__4154),
            .I(N__4146));
    LocalMux I__404 (
            .O(N__4151),
            .I(N__4146));
    Sp12to4 I__403 (
            .O(N__4146),
            .I(N__4143));
    Span12Mux_v I__402 (
            .O(N__4143),
            .I(N__4140));
    Odrv12 I__401 (
            .O(N__4140),
            .I(A_c_24));
    InMux I__400 (
            .O(N__4137),
            .I(N__4131));
    InMux I__399 (
            .O(N__4136),
            .I(N__4131));
    LocalMux I__398 (
            .O(N__4131),
            .I(N__4128));
    Sp12to4 I__397 (
            .O(N__4128),
            .I(N__4125));
    Span12Mux_v I__396 (
            .O(N__4125),
            .I(N__4122));
    Odrv12 I__395 (
            .O(N__4122),
            .I(A_c_26));
    InMux I__394 (
            .O(N__4119),
            .I(N__4113));
    InMux I__393 (
            .O(N__4118),
            .I(N__4113));
    LocalMux I__392 (
            .O(N__4113),
            .I(N__4110));
    Span4Mux_v I__391 (
            .O(N__4110),
            .I(N__4107));
    Sp12to4 I__390 (
            .O(N__4107),
            .I(N__4104));
    Odrv12 I__389 (
            .O(N__4104),
            .I(A_c_27));
    InMux I__388 (
            .O(N__4101),
            .I(N__4098));
    LocalMux I__387 (
            .O(N__4098),
            .I(\U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_5 ));
    InMux I__386 (
            .O(N__4095),
            .I(N__4092));
    LocalMux I__385 (
            .O(N__4092),
            .I(N__4089));
    Odrv4 I__384 (
            .O(N__4089),
            .I(\U409_AUTOCONFIG.N_42 ));
    CascadeMux I__383 (
            .O(N__4086),
            .I(\U409_AUTOCONFIG.N_111_cascade_ ));
    CascadeMux I__382 (
            .O(N__4083),
            .I(\U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0_a3_0Z0Z_2_cascade_ ));
    IoInMux I__381 (
            .O(N__4080),
            .I(N__4077));
    LocalMux I__380 (
            .O(N__4077),
            .I(N__4074));
    IoSpan4Mux I__379 (
            .O(N__4074),
            .I(N__4071));
    Span4Mux_s3_h I__378 (
            .O(N__4071),
            .I(N__4068));
    Sp12to4 I__377 (
            .O(N__4068),
            .I(N__4065));
    Span12Mux_h I__376 (
            .O(N__4065),
            .I(N__4062));
    Span12Mux_h I__375 (
            .O(N__4062),
            .I(N__4059));
    Odrv12 I__374 (
            .O(N__4059),
            .I(A_c_15));
    IoInMux I__373 (
            .O(N__4056),
            .I(N__4053));
    LocalMux I__372 (
            .O(N__4053),
            .I(N__4050));
    Span4Mux_s3_h I__371 (
            .O(N__4050),
            .I(N__4047));
    Span4Mux_v I__370 (
            .O(N__4047),
            .I(N__4044));
    Sp12to4 I__369 (
            .O(N__4044),
            .I(N__4041));
    Span12Mux_h I__368 (
            .O(N__4041),
            .I(N__4038));
    Span12Mux_h I__367 (
            .O(N__4038),
            .I(N__4035));
    Odrv12 I__366 (
            .O(N__4035),
            .I(A_c_14));
    ClkMux I__365 (
            .O(N__4032),
            .I(N__3990));
    ClkMux I__364 (
            .O(N__4031),
            .I(N__3990));
    ClkMux I__363 (
            .O(N__4030),
            .I(N__3990));
    ClkMux I__362 (
            .O(N__4029),
            .I(N__3990));
    ClkMux I__361 (
            .O(N__4028),
            .I(N__3990));
    ClkMux I__360 (
            .O(N__4027),
            .I(N__3990));
    ClkMux I__359 (
            .O(N__4026),
            .I(N__3990));
    ClkMux I__358 (
            .O(N__4025),
            .I(N__3990));
    ClkMux I__357 (
            .O(N__4024),
            .I(N__3990));
    ClkMux I__356 (
            .O(N__4023),
            .I(N__3990));
    ClkMux I__355 (
            .O(N__4022),
            .I(N__3990));
    ClkMux I__354 (
            .O(N__4021),
            .I(N__3990));
    ClkMux I__353 (
            .O(N__4020),
            .I(N__3990));
    ClkMux I__352 (
            .O(N__4019),
            .I(N__3990));
    GlobalMux I__351 (
            .O(N__3990),
            .I(CLK80_OUT));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .I(N__4029));
    INV \INVU409_TRANSFER_ACK.LASTCLK_1C  (
            .O(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .I(N__4021));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .I(N__4026));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .I(N__4024));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .I(N__4022));
    INV \INVU409_TRANSFER_ACK.CIA_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .I(N__4020));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .I(N__4019));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .I(N__4027));
    INV \INVU409_TRANSFER_ACK.TACK_OUTnC  (
            .O(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .I(N__4025));
    INV \INVU409_TRANSFER_ACK.TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.TACK_ENC_net ),
            .I(N__4023));
    INV \INVU409_TRANSFER_ACK.ROMENn_nessC  (
            .O(\INVU409_TRANSFER_ACK.ROMENn_nessC_net ),
            .I(N__4032));
    INV \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC  (
            .O(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .I(N__4028));
    INV \INVU409_AUTOCONFIG.ATA_BASE_2C  (
            .O(\INVU409_AUTOCONFIG.ATA_BASE_2C_net ),
            .I(N__8262));
    INV \INVU409_AUTOCONFIG.ATA_BASE_4C  (
            .O(\INVU409_AUTOCONFIG.ATA_BASE_4C_net ),
            .I(N__8263));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .I(N__4031));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net ),
            .I(N__4030));
    INV \INVU409_AUTOCONFIG.CONFIGENnC  (
            .O(\INVU409_AUTOCONFIG.CONFIGENnC_net ),
            .I(N__8267));
    INV \INVU409_AUTOCONFIG.LIDE_CONFC  (
            .O(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .I(N__8266));
    INV \INVU409_AUTOCONFIG.BRIDGE_OUT_1C  (
            .O(\INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net ),
            .I(N__8268));
    INV \INVU409_AUTOCONFIG.BRIDGE_OUT_0C  (
            .O(\INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ),
            .I(N__8270));
    INV \INVU409_AUTOCONFIG.LIDE_OUT_3C  (
            .O(\INVU409_AUTOCONFIG.LIDE_OUT_3C_net ),
            .I(N__8269));
    defparam IN_MUX_bfv_13_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_6_0_));
    defparam IN_MUX_bfv_13_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_7_0_ (
            .carryinitin(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .carryinitout(bfn_13_7_0_));
    defparam IN_MUX_bfv_14_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_5_0_));
    defparam IN_MUX_bfv_14_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_6_0_ (
            .carryinitin(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .carryinitout(bfn_14_6_0_));
    defparam IN_MUX_bfv_16_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_7_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__8169),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_4_0_LC_3_10_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_4_0_LC_3_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_4_0_LC_3_10_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_4_0_LC_3_10_1  (
            .in0(N__4192),
            .in1(N__4212),
            .in2(_gnd_net_),
            .in3(N__4725),
            .lcout(\U409_AUTOCONFIG.N_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_11_3_i_o3_LC_3_10_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_11_3_i_o3_LC_3_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_11_3_i_o3_LC_3_10_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U409_AUTOCONFIG.un1_A_11_3_i_o3_LC_3_10_2  (
            .in0(N__4214),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4194),
            .lcout(\U409_AUTOCONFIG.N_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0_a3_0_2_LC_3_10_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0_a3_0_2_LC_3_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0_a3_0_2_LC_3_10_4 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0_a3_0_2_LC_3_10_4  (
            .in0(N__4726),
            .in1(N__6342),
            .in2(N__4872),
            .in3(N__4948),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0_a3_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0_0_LC_3_10_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0_0_LC_3_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0_0_LC_3_10_5 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0_0_LC_3_10_5  (
            .in0(N__4294),
            .in1(N__4949),
            .in2(N__4083),
            .in3(N__10187),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_3_10_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_3_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_3_10_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_3_10_6  (
            .in0(N__4241),
            .in1(N__4293),
            .in2(N__4871),
            .in3(N__4947),
            .lcout(\U409_AUTOCONFIG.N_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_1_sqmuxa_0_a2_0_2_LC_3_10_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_1_sqmuxa_0_a2_0_2_LC_3_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_1_sqmuxa_0_a2_0_2_LC_3_10_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_1_sqmuxa_0_a2_0_2_LC_3_10_7  (
            .in0(N__4193),
            .in1(N__4782),
            .in2(N__4739),
            .in3(N__4213),
            .lcout(\U409_AUTOCONFIG.LIDE_CONF_1_sqmuxa_0_a2_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_5_0_LC_3_11_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_5_0_LC_3_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_5_0_LC_3_11_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_5_0_LC_3_11_4  (
            .in0(N__4221),
            .in1(N__6341),
            .in2(N__4184),
            .in3(N__4724),
            .lcout(\U409_AUTOCONFIG.N_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_3_14_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_3_14_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_3_14_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_3_14_3  (
            .in0(N__7027),
            .in1(N__5852),
            .in2(_gnd_net_),
            .in3(N__4160),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_3_14_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_3_14_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_3_14_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_3_14_4  (
            .in0(N__4397),
            .in1(N__10191),
            .in2(N__4164),
            .in3(N__4101),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACE ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_7_LC_3_15_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_7_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_7_LC_3_15_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_7_LC_3_15_1  (
            .in0(N__4119),
            .in1(N__4422),
            .in2(N__4161),
            .in3(N__4137),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_5_LC_3_15_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_5_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_5_LC_3_15_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_5_LC_3_15_6  (
            .in0(N__4136),
            .in1(N__5980),
            .in2(N__5903),
            .in3(N__4118),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_4_LC_5_10_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_4_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_4_LC_5_10_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_4_LC_5_10_1  (
            .in0(N__6114),
            .in1(N__5610),
            .in2(N__6032),
            .in3(N__4626),
            .lcout(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_o2_0_LC_5_10_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_o2_0_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_o2_0_LC_5_10_3 .LUT_INIT=16'b0011011100110011;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_o2_0_LC_5_10_3  (
            .in0(N__6359),
            .in1(N__10148),
            .in2(N__5001),
            .in3(N__4769),
            .lcout(\U409_AUTOCONFIG.N_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_6_0_LC_5_10_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_6_0_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_6_0_LC_5_10_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_6_0_LC_5_10_4  (
            .in0(N__4873),
            .in1(N__4311),
            .in2(_gnd_net_),
            .in3(N__4295),
            .lcout(\U409_AUTOCONFIG.N_111 ),
            .ltout(\U409_AUTOCONFIG.N_111_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_5_10_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_5_10_5 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_5_10_5  (
            .in0(N__6358),
            .in1(N__4095),
            .in2(N__4086),
            .in3(N__4960),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_5_10_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_5_10_6 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_5_10_6  (
            .in0(N__4768),
            .in1(N__4477),
            .in2(N__4314),
            .in3(N__4310),
            .lcout(\U409_AUTOCONFIG.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_3_1_LC_5_10_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_3_1_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_3_1_LC_5_10_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_3_1_LC_5_10_7  (
            .in0(N__4296),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4874),
            .lcout(\U409_AUTOCONFIG.N_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.HIROM_2_i_o3_LC_5_11_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.HIROM_2_i_o3_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.HIROM_2_i_o3_LC_5_11_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U409_ADDRESS_DECODE.HIROM_2_i_o3_LC_5_11_0  (
            .in0(N__6481),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7150),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.N_54_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.HIROM_LC_5_11_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.HIROM_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.HIROM_LC_5_11_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.HIROM_LC_5_11_1  (
            .in0(N__6115),
            .in1(N__6924),
            .in2(N__4299),
            .in3(N__6574),
            .lcout(\U409_ADDRESS_DECODE.HIROMZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_5_11_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_5_11_2 .LUT_INIT=16'b0001000001000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_5_11_2  (
            .in0(N__4705),
            .in1(N__6352),
            .in2(N__4862),
            .in3(N__4959),
            .lcout(\U409_AUTOCONFIG.N_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_5_11_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_5_11_3 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_5_11_3  (
            .in0(N__4478),
            .in1(N__4278),
            .in2(N__4251),
            .in3(N__4843),
            .lcout(\U409_AUTOCONFIG.N_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_3_0_LC_5_11_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_3_0_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_3_0_LC_5_11_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_3_0_LC_5_11_4  (
            .in0(N__4844),
            .in1(N__4279),
            .in2(_gnd_net_),
            .in3(N__4958),
            .lcout(\U409_AUTOCONFIG.N_86 ),
            .ltout(\U409_AUTOCONFIG.N_86_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_5_11_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_5_11_5 .LUT_INIT=16'b1111111110110011;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_5_11_5  (
            .in0(N__4250),
            .in1(N__10149),
            .in2(N__4230),
            .in3(N__4227),
            .lcout(\U409_AUTOCONFIG.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_3_LC_5_12_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_3_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_3_LC_5_12_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_3_LC_5_12_5  (
            .in0(N__4494),
            .in1(N__6351),
            .in2(_gnd_net_),
            .in3(N__4904),
            .lcout(\U409_AUTOCONFIG.N_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_3_LC_5_12_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_3_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_3_LC_5_12_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_3_LC_5_12_7  (
            .in0(N__6480),
            .in1(N__4652),
            .in2(N__7166),
            .in3(N__4634),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3_0_1_LC_5_13_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3_0_1_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3_0_1_LC_5_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3_0_1_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(N__6573),
            .in2(_gnd_net_),
            .in3(N__6925),
            .lcout(N_89_1),
            .ltout(N_89_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3_0_LC_5_13_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3_0_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3_0_LC_5_13_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3_0_LC_5_13_6  (
            .in0(N__4653),
            .in1(N__6479),
            .in2(N__4410),
            .in3(N__7146),
            .lcout(\U409_ADDRESS_DECODE.N_102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_11_LC_5_14_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_11_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_11_LC_5_14_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_11_LC_5_14_2  (
            .in0(N__4407),
            .in1(N__10176),
            .in2(N__4341),
            .in3(N__4398),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_9_LC_5_17_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_9_LC_5_17_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_9_LC_5_17_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_9_LC_5_17_3  (
            .in0(N__5902),
            .in1(N__4371),
            .in2(N__4359),
            .in3(N__5981),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_0_3_163_i_i_o2_LC_6_9_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_0_3_163_i_i_o2_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_0_3_163_i_i_o2_LC_6_9_1 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_0_3_163_i_i_o2_LC_6_9_1  (
            .in0(N__4778),
            .in1(N__10169),
            .in2(_gnd_net_),
            .in3(N__6372),
            .lcout(\U409_AUTOCONFIG.N_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_6_10_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_6_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_6_10_0 .LUT_INIT=16'b1111000100000001;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_3_LC_6_10_0  (
            .in0(N__4329),
            .in1(N__4461),
            .in2(N__5193),
            .in3(N__5234),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_3C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_6_10_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_6_10_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_6_10_1 .LUT_INIT=16'b1111000000010001;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_2_LC_6_10_1  (
            .in0(N__4788),
            .in1(N__4328),
            .in2(N__5285),
            .in3(N__5188),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_3C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_6_10_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_6_10_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_6_10_2 .LUT_INIT=16'b1111000100000001;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_0_LC_6_10_2  (
            .in0(N__4320),
            .in1(N__4659),
            .in2(N__5192),
            .in3(N__4541),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_3C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_2_LC_6_10_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_2_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_2_LC_6_10_3 .LUT_INIT=16'b1111111101001000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_2_LC_6_10_3  (
            .in0(N__6353),
            .in1(N__4490),
            .in2(N__4974),
            .in3(N__4479),
            .lcout(\U409_AUTOCONFIG.N_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_6_10_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_6_10_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_6_10_5  (
            .in0(N__4964),
            .in1(N__4878),
            .in2(N__6379),
            .in3(N__4723),
            .lcout(\U409_AUTOCONFIG.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_6_10_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_6_10_6 .LUT_INIT=16'b0101110101010101;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_6_10_6  (
            .in0(N__10170),
            .in1(N__4455),
            .in2(N__4977),
            .in3(N__6357),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_6_10_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_6_10_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_6_10_7 .LUT_INIT=16'b1100110000000101;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_1_LC_6_10_7  (
            .in0(N__4428),
            .in1(N__5345),
            .in2(N__4449),
            .in3(N__5184),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_3C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a2_LC_6_11_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a2_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a2_LC_6_11_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a2_LC_6_11_0  (
            .in0(N__6907),
            .in1(N__6487),
            .in2(_gnd_net_),
            .in3(N__7161),
            .lcout(\U409_ADDRESS_DECODE.N_112 ),
            .ltout(\U409_ADDRESS_DECODE.N_112_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_LC_6_11_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_LC_6_11_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_LC_6_11_1  (
            .in0(N__7189),
            .in1(N__4446),
            .in2(N__4440),
            .in3(N__6580),
            .lcout(AUTOCONFIG_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3_0_2_LC_6_11_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3_0_2_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3_0_2_LC_6_11_2 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3_0_2_LC_6_11_2  (
            .in0(N__6045),
            .in1(N__4437),
            .in2(_gnd_net_),
            .in3(N__6131),
            .lcout(\U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_6_11_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_6_11_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_6_11_3  (
            .in0(N__4743),
            .in1(N__6362),
            .in2(N__4976),
            .in3(N__4852),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.N_74_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_6_11_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_6_11_4 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_6_11_4  (
            .in0(N__6360),
            .in1(N__4770),
            .in2(N__4431),
            .in3(N__4740),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_6_11_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_6_11_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_6_11_5  (
            .in0(N__4741),
            .in1(N__6361),
            .in2(N__4975),
            .in3(N__4851),
            .lcout(\U409_AUTOCONFIG.N_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_6_11_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_6_11_6 .LUT_INIT=16'b0101010111011101;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_6_11_6  (
            .in0(N__10147),
            .in1(N__4771),
            .in2(_gnd_net_),
            .in3(N__4742),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_1_85_i_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a2_0_LC_6_12_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a2_0_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a2_0_LC_6_12_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a2_0_LC_6_12_2  (
            .in0(N__6046),
            .in1(N__6133),
            .in2(_gnd_net_),
            .in3(N__5617),
            .lcout(N_121),
            .ltout(N_121_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_1_LC_6_12_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_1_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_1_LC_6_12_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_1_LC_6_12_3  (
            .in0(N__6893),
            .in1(_gnd_net_),
            .in2(N__4641),
            .in3(N__4630),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_13_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_13_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_13_0  (
            .in0(N__4566),
            .in1(N__4560),
            .in2(N__5478),
            .in3(N__6485),
            .lcout(CIA_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_6_13_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_6_13_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_6_13_7  (
            .in0(N__7159),
            .in1(N__5734),
            .in2(N__5665),
            .in3(N__6575),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_10_LC_6_14_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_10_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_10_LC_6_14_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_10_LC_6_14_6  (
            .in0(N__7032),
            .in1(N__4554),
            .in2(_gnd_net_),
            .in3(N__5845),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIA2DB1_0_LC_7_9_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIA2DB1_0_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIA2DB1_0_LC_7_9_2 .LUT_INIT=16'b1111101011001010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNIA2DB1_0_LC_7_9_2  (
            .in0(N__4542),
            .in1(N__4505),
            .in2(N__6230),
            .in3(N__5710),
            .lcout(U409_AUTOCONFIG_D_OUT_0_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_7_9_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_7_9_3 .LUT_INIT=16'b1101000101010101;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_7_9_3  (
            .in0(N__4518),
            .in1(N__10153),
            .in2(N__4506),
            .in3(N__5018),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_7_9_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_7_9_6 .LUT_INIT=16'b1011001100010011;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_7_9_6  (
            .in0(N__5019),
            .in1(N__5082),
            .in2(N__10177),
            .in3(N__5255),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_7_10_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_7_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_7_10_0 .LUT_INIT=16'b1101000101010101;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_7_10_0  (
            .in0(N__5070),
            .in1(N__10160),
            .in2(N__5333),
            .in3(N__5016),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_0_LC_7_10_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_0_LC_7_10_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.STATE_0_LC_7_10_1 .LUT_INIT=16'b0010000011110000;
    LogicCell40 \U409_AUTOCONFIG.STATE_0_LC_7_10_1  (
            .in0(N__5791),
            .in1(N__5770),
            .in2(N__10180),
            .in3(N__5028),
            .lcout(\U409_AUTOCONFIG.STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNIU6QK1_0_LC_7_10_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNIU6QK1_0_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNIU6QK1_0_LC_7_10_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNIU6QK1_0_LC_7_10_2  (
            .in0(N__5769),
            .in1(N__5058),
            .in2(_gnd_net_),
            .in3(N__5790),
            .lcout(\U409_AUTOCONFIG.N_122 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_7_10_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_7_10_3 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_7_10_3 .LUT_INIT=16'b1011001100010011;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_7_10_3  (
            .in0(N__5017),
            .in1(N__5049),
            .in2(N__10179),
            .in3(N__5303),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_1_LC_7_10_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_1_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.STATE_1_LC_7_10_4 .LUT_INIT=16'b0100010000001000;
    LogicCell40 \U409_AUTOCONFIG.STATE_1_LC_7_10_4  (
            .in0(N__5771),
            .in1(N__10167),
            .in2(N__5549),
            .in3(N__5792),
            .lcout(\U409_AUTOCONFIG.STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_ns_1_0__m2_0_o2_LC_7_10_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_ns_1_0__m2_0_o2_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_ns_1_0__m2_0_o2_LC_7_10_5 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \U409_AUTOCONFIG.STATE_ns_1_0__m2_0_o2_LC_7_10_5  (
            .in0(N__5040),
            .in1(N__5768),
            .in2(_gnd_net_),
            .in3(N__5118),
            .lcout(\U409_AUTOCONFIG.N_52 ),
            .ltout(\U409_AUTOCONFIG.N_52_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNIBM2Q1_1_LC_7_10_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNIBM2Q1_1_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNIBM2Q1_1_LC_7_10_6 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNIBM2Q1_1_LC_7_10_6  (
            .in0(N__5543),
            .in1(_gnd_net_),
            .in2(N__5022),
            .in3(N__5789),
            .lcout(\U409_AUTOCONFIG.N_56 ),
            .ltout(\U409_AUTOCONFIG.N_56_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNI7U5N3_1_LC_7_10_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNI7U5N3_1_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNI7U5N3_1_LC_7_10_7 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNI7U5N3_1_LC_7_10_7  (
            .in0(N__10168),
            .in1(N__5000),
            .in2(N__4980),
            .in3(N__5202),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.LOWROM_2_LC_7_11_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.LOWROM_2_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.LOWROM_2_LC_7_11_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.LOWROM_2_LC_7_11_4  (
            .in0(N__7162),
            .in1(N__6584),
            .in2(N__6492),
            .in3(N__6923),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.LOWROMZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_ROMEN_LC_7_11_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_ROMEN_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_ROMEN_LC_7_11_5 .LUT_INIT=16'b0101010100010101;
    LogicCell40 \U409_ADDRESS_DECODE.un1_ROMEN_LC_7_11_5  (
            .in0(N__5172),
            .in1(N__7077),
            .in2(N__5163),
            .in3(N__6132),
            .lcout(U409_ADDRESS_DECODE_un1_ROMEN_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_7_11_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_7_11_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \U409_ADDRESS_DECODE.D_1_i_LC_7_11_6  (
            .in0(N__5539),
            .in1(N__10268),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(D_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_START_LC_7_11_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_START_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.AC_START_LC_7_11_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_AUTOCONFIG.AC_START_LC_7_11_7  (
            .in0(N__10269),
            .in1(N__8349),
            .in2(_gnd_net_),
            .in3(N__5703),
            .lcout(\U409_AUTOCONFIG.AC_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8265),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_1_LC_7_12_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_1_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_1_LC_7_12_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_1_LC_7_12_0  (
            .in0(N__5667),
            .in1(N__5750),
            .in2(N__6590),
            .in3(N__5625),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_4_LC_7_12_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_4_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_4_LC_7_12_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_4_LC_7_12_1  (
            .in0(N__6134),
            .in1(N__6486),
            .in2(N__5112),
            .in3(N__6047),
            .lcout(\U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2Z0Z_4 ),
            .ltout(\U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_7_12_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_7_12_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_7_12_2  (
            .in0(N__5472),
            .in1(N__6906),
            .in2(N__5109),
            .in3(N__7160),
            .lcout(N_120),
            .ltout(N_120_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_7_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_7_12_3 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_7_12_3  (
            .in0(N__5106),
            .in1(_gnd_net_),
            .in2(N__5097),
            .in3(N__5094),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_1_0_a2_LC_7_12_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_1_0_a2_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_1_0_a2_LC_7_12_7 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_1_0_a2_LC_7_12_7  (
            .in0(N__5749),
            .in1(N__5666),
            .in2(_gnd_net_),
            .in3(N__5471),
            .lcout(U409_ADDRESS_DECODE_ROMEN_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_7_13_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_7_13_6 .LUT_INIT=16'b0011000111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_7_13_6  (
            .in0(N__5364),
            .in1(N__5376),
            .in2(N__6589),
            .in3(N__5470),
            .lcout(U409_ADDRESS_DECODE_un1_REGSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_7_13_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_7_13_7 .LUT_INIT=16'b1010000011100000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_7_13_7  (
            .in0(N__5375),
            .in1(N__5363),
            .in2(N__5479),
            .in3(N__6576),
            .lcout(U409_ADDRESS_DECODE_un1_REGSPACEn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIC4DB1_1_LC_8_8_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIC4DB1_1_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIC4DB1_1_LC_8_8_4 .LUT_INIT=16'b1111101011001010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNIC4DB1_1_LC_8_8_4  (
            .in0(N__5352),
            .in1(N__5334),
            .in2(N__6231),
            .in3(N__5712),
            .lcout(U409_AUTOCONFIG_D_OUT_0_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIE6DB1_2_LC_8_9_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIE6DB1_2_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIE6DB1_2_LC_8_9_0 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNIE6DB1_2_LC_8_9_0  (
            .in0(N__5304),
            .in1(N__5705),
            .in2(N__5292),
            .in3(N__6211),
            .lcout(U409_AUTOCONFIG_D_OUT_0_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_LC_8_9_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_LC_8_9_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_LC_8_9_2  (
            .in0(N__6383),
            .in1(N__6210),
            .in2(_gnd_net_),
            .in3(N__6163),
            .lcout(\U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIG8DB1_3_LC_8_9_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIG8DB1_3_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIG8DB1_3_LC_8_9_4 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNIG8DB1_3_LC_8_9_4  (
            .in0(N__5256),
            .in1(N__5706),
            .in2(N__5244),
            .in3(N__6212),
            .lcout(U409_AUTOCONFIG_D_OUT_0_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_8_10_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_8_10_0 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_LC_8_10_0  (
            .in0(N__6215),
            .in1(N__6371),
            .in2(_gnd_net_),
            .in3(N__6166),
            .lcout(\U409_AUTOCONFIG.LIDE_CONFZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .ce(),
            .sr(N__9028));
    defparam \U409_AUTOCONFIG.CONFIGURED_LC_8_10_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.CONFIGURED_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.CONFIGURED_LC_8_10_1 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \U409_AUTOCONFIG.CONFIGURED_LC_8_10_1  (
            .in0(N__6167),
            .in1(N__6216),
            .in2(N__6382),
            .in3(N__5704),
            .lcout(CONFIGURED),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .ce(),
            .sr(N__9028));
    defparam \U409_AUTOCONFIG.AC_TACK_LC_8_10_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_TACK_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.AC_TACK_LC_8_10_2 .LUT_INIT=16'b1110111011001000;
    LogicCell40 \U409_AUTOCONFIG.AC_TACK_LC_8_10_2  (
            .in0(N__5793),
            .in1(N__5772),
            .in2(N__5550),
            .in3(N__7544),
            .lcout(AC_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .ce(),
            .sr(N__9028));
    defparam \U409_AUTOCONFIG.ATA_BASE_3_LC_8_10_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_3_LC_8_10_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.ATA_BASE_3_LC_8_10_4 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_3_LC_8_10_4  (
            .in0(N__7326),
            .in1(N__7292),
            .in2(N__6708),
            .in3(N__6063),
            .lcout(ATA_BASE_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .ce(),
            .sr(N__9028));
    defparam \U409_AUTOCONFIG.ATA_BASE_1_LC_8_10_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_1_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.ATA_BASE_1_LC_8_10_6 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_1_LC_8_10_6  (
            .in0(N__7325),
            .in1(N__7291),
            .in2(N__7432),
            .in3(N__5568),
            .lcout(ATA_BASE_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .ce(),
            .sr(N__9028));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_8_11_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_8_11_0 .LUT_INIT=16'b0101000010100000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_8_11_0  (
            .in0(N__5751),
            .in1(_gnd_net_),
            .in2(N__5711),
            .in3(N__5656),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1 ),
            .ltout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_4_LC_8_11_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_4_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_4_LC_8_11_1 .LUT_INIT=16'b1000000001000000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_4_LC_8_11_1  (
            .in0(N__5624),
            .in1(N__5480),
            .in2(N__5571),
            .in3(N__5567),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_LC_8_11_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_LC_8_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_LC_8_11_2  (
            .in0(N__6390),
            .in1(N__5994),
            .in2(N__5556),
            .in3(N__6846),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACEZ0 ),
            .ltout(\U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_LC_8_11_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_LC_8_11_3 .SEQ_MODE=4'b1000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_LC_8_11_3 .LUT_INIT=16'b1100110001000000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_LC_8_11_3  (
            .in0(N__5544),
            .in1(N__10178),
            .in2(N__5553),
            .in3(N__6805),
            .lcout(\U409_ADDRESS_DECODE.ATA_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8264),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_0_a3_LC_8_11_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_0_a3_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_0_a3_LC_8_11_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_0_a3_LC_8_11_4  (
            .in0(N__10279),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5545),
            .lcout(un1_AUTOCONFIG_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.N_120_i_LC_8_11_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.N_120_i_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.N_120_i_LC_8_11_6 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \U409_ADDRESS_DECODE.N_120_i_LC_8_11_6  (
            .in0(N__5490),
            .in1(N__7167),
            .in2(N__5484),
            .in3(N__6932),
            .lcout(N_120_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_1_LC_8_12_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_1_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_1_LC_8_12_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_1_LC_8_12_0  (
            .in0(N__7624),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7913),
            .lcout(\U409_TRANSFER_ACK.CO1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_3_LC_8_12_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_3_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_3_LC_8_12_2 .LUT_INIT=16'b1000010000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_3_LC_8_12_2  (
            .in0(N__6663),
            .in1(N__5988),
            .in2(N__5982),
            .in3(N__5820),
            .lcout(\U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_1_LC_8_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_1_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_1_LC_8_12_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_1_LC_8_12_3  (
            .in0(N__7599),
            .in1(N__7622),
            .in2(N__7921),
            .in3(N__7865),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.LOWROM_3_LC_8_12_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.LOWROM_3_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.LOWROM_3_LC_8_12_4 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \U409_ADDRESS_DECODE.LOWROM_3_LC_8_12_4  (
            .in0(N__6588),
            .in1(N__6491),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_ADDRESS_DECODE.LOWROMZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_1_LC_8_12_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_1_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_1_LC_8_12_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_1_LC_8_12_6  (
            .in0(N__7623),
            .in1(N__7598),
            .in2(N__7876),
            .in3(N__7909),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_LC_8_13_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_LC_8_13_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_0_LC_8_13_3  (
            .in0(N__10231),
            .in1(N__10288),
            .in2(_gnd_net_),
            .in3(N__5937),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.PORTSIZEZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNI4345U_LC_8_13_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNI4345U_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNI4345U_LC_8_13_4 .LUT_INIT=16'b1110111111001111;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_RNI4345U_LC_8_13_4  (
            .in0(N__7760),
            .in1(N__7724),
            .in2(N__5931),
            .in3(N__6810),
            .lcout(PORTSIZE_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_0_LC_8_13_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_0_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_0_LC_8_13_5 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_0_LC_8_13_5  (
            .in0(N__6648),
            .in1(N__5907),
            .in2(N__5862),
            .in3(N__6627),
            .lcout(\U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_9_9_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_9_9_0 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_9_9_0 .LUT_INIT=16'b1000101010101010;
    LogicCell40 \U409_AUTOCONFIG.CONFIGENn_LC_9_9_0  (
            .in0(N__5804),
            .in1(N__6384),
            .in2(N__6226),
            .in3(N__6171),
            .lcout(CONFIGENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.CONFIGENnC_net ),
            .ce(),
            .sr(N__9029));
    defparam \U409_AUTOCONFIG.ATA_BASE_7_LC_9_9_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_7_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.ATA_BASE_7_LC_9_9_1 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_7_LC_9_9_1  (
            .in0(N__7346),
            .in1(N__7386),
            .in2(N__6697),
            .in3(N__6504),
            .lcout(ATA_BASE_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.CONFIGENnC_net ),
            .ce(),
            .sr(N__9029));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_9_9_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_9_9_3 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_9_9_3 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_9_9_3  (
            .in0(N__7352),
            .in1(N__6609),
            .in2(N__6698),
            .in3(N__6659),
            .lcout(BRIDGE_BASE_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.CONFIGENnC_net ),
            .ce(),
            .sr(N__9029));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_9_9_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_9_9_4 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_9_9_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_9_9_4  (
            .in0(N__7264),
            .in1(N__7351),
            .in2(N__6644),
            .in3(N__6608),
            .lcout(BRIDGE_BASE_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.CONFIGENnC_net ),
            .ce(),
            .sr(N__9029));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_9_9_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_9_9_5 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_9_9_5 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_9_9_5  (
            .in0(N__6606),
            .in1(N__7439),
            .in2(N__7356),
            .in3(N__6620),
            .lcout(BRIDGE_BASE_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.CONFIGENnC_net ),
            .ce(),
            .sr(N__9029));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_9_9_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_9_9_6 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_9_9_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_9_9_6  (
            .in0(N__7484),
            .in1(N__7347),
            .in2(N__6986),
            .in3(N__6607),
            .lcout(BRIDGE_BASE_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.CONFIGENnC_net ),
            .ce(),
            .sr(N__9029));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_9_10_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_9_10_2 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_9_10_2  (
            .in0(N__6591),
            .in1(N__6503),
            .in2(N__6478),
            .in3(N__7367),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_1_LC_9_10_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_1_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_1_LC_9_10_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_1_LC_9_10_3  (
            .in0(N__6381),
            .in1(N__6214),
            .in2(_gnd_net_),
            .in3(N__6165),
            .lcout(\U409_AUTOCONFIG.LIDE_CONF_RNIUPP42Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_0_LC_9_10_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_0_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_0_LC_9_10_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_0_LC_9_10_7  (
            .in0(N__6380),
            .in1(N__6213),
            .in2(_gnd_net_),
            .in3(N__6164),
            .lcout(\U409_AUTOCONFIG.LIDE_CONF_RNIUPP42Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_9_11_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_9_11_0 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_9_11_0  (
            .in0(N__6135),
            .in1(N__6062),
            .in2(N__6051),
            .in3(N__7232),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_1_0_LC_9_11_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_1_0_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_1_0_LC_9_11_1 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_1_0_LC_9_11_1  (
            .in0(N__7168),
            .in1(N__7397),
            .in2(N__6936),
            .in3(N__7460),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACE_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_9_11_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_9_11_4 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_9_11_4  (
            .in0(N__7202),
            .in1(N__7066),
            .in2(N__7221),
            .in3(N__7169),
            .lcout(U409_ADDRESS_DECODE_un1_RAMSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_9_11_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_9_11_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_9_11_5  (
            .in0(N__6819),
            .in1(N__8367),
            .in2(N__8306),
            .in3(N__7203),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNI206O6_LC_9_11_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNI206O6_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNI206O6_LC_9_11_7 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_RNI206O6_LC_9_11_7  (
            .in0(N__7753),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6806),
            .lcout(U409_ADDRESS_DECODE_un1_ATA_ENn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_9_12_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_9_12_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_9_12_1 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_9_12_1  (
            .in0(N__7601),
            .in1(N__6768),
            .in2(N__6720),
            .in3(N__7869),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net ),
            .ce(),
            .sr(N__9023));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_9_12_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_9_12_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_9_12_2 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_9_12_2  (
            .in0(N__6767),
            .in1(N__6716),
            .in2(_gnd_net_),
            .in3(N__7602),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net ),
            .ce(),
            .sr(N__9023));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_9_12_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_9_12_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_9_12_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(N__7914),
            .in2(_gnd_net_),
            .in3(N__7626),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net ),
            .ce(),
            .sr(N__9023));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_9_13_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_9_13_1 .LUT_INIT=16'b0000111000000101;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_9_13_1  (
            .in0(N__7925),
            .in1(N__6747),
            .in2(N__6735),
            .in3(N__6759),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__9019));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIL9Q68_1_LC_9_13_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIL9Q68_1_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIL9Q68_1_LC_9_13_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIL9Q68_1_LC_9_13_5  (
            .in0(N__6758),
            .in1(N__6746),
            .in2(_gnd_net_),
            .in3(N__6731),
            .lcout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0 ),
            .ltout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_ness_RNO_LC_9_13_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_ness_RNO_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_ness_RNO_LC_9_13_6 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_ness_RNO_LC_9_13_6  (
            .in0(N__9033),
            .in1(_gnd_net_),
            .in2(N__7497),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.ATA_BASE_4_LC_10_10_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_4_LC_10_10_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.ATA_BASE_4_LC_10_10_2 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_4_LC_10_10_2  (
            .in0(N__7353),
            .in1(N__7383),
            .in2(N__7494),
            .in3(N__7461),
            .lcout(ATA_BASE_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_4C_net ),
            .ce(),
            .sr(N__9026));
    defparam \U409_AUTOCONFIG.ATA_BASE_5_LC_10_10_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_5_LC_10_10_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.ATA_BASE_5_LC_10_10_4 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_5_LC_10_10_4  (
            .in0(N__7354),
            .in1(N__7384),
            .in2(N__7449),
            .in3(N__7398),
            .lcout(ATA_BASE_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_4C_net ),
            .ce(),
            .sr(N__9026));
    defparam \U409_AUTOCONFIG.ATA_BASE_6_LC_10_10_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_6_LC_10_10_6 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.ATA_BASE_6_LC_10_10_6 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_6_LC_10_10_6  (
            .in0(N__7355),
            .in1(N__7385),
            .in2(N__7277),
            .in3(N__7368),
            .lcout(ATA_BASE_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_4C_net ),
            .ce(),
            .sr(N__9026));
    defparam \U409_AUTOCONFIG.ATA_BASE_2_LC_10_11_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_2_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.ATA_BASE_2_LC_10_11_1 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_2_LC_10_11_1  (
            .in0(N__7338),
            .in1(N__7293),
            .in2(N__7278),
            .in3(N__7233),
            .lcout(ATA_BASE_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_2C_net ),
            .ce(),
            .sr(N__9024));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_10_12_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_10_12_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_10_12_1  (
            .in0(N__7220),
            .in1(N__7196),
            .in2(N__7173),
            .in3(N__7073),
            .lcout(U409_ADDRESS_DECODE_un1_RAMSPACEn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_12_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_12_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_12_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_12_2  (
            .in0(N__8303),
            .in1(N__8368),
            .in2(N__7817),
            .in3(N__7829),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_LC_10_12_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_LC_10_12_3 .LUT_INIT=16'b0111101111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_LC_10_12_3  (
            .in0(N__7031),
            .in1(N__10080),
            .in2(N__6990),
            .in3(N__6969),
            .lcout(U409_ADDRESS_DECODE_un1_BRIDGE_ENn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_10_12_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_10_12_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_10_12_7  (
            .in0(_gnd_net_),
            .in1(N__7625),
            .in2(_gnd_net_),
            .in3(N__7600),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_ness_LC_10_14_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_ness_LC_10_14_1 .SEQ_MODE=4'b1001;
    defparam \U409_TRANSFER_ACK.ROMENn_ness_LC_10_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_ness_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7878),
            .lcout(ROMENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROMENn_nessC_net ),
            .ce(N__7560),
            .sr(N__9016));
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_11_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_11_10_0 .LUT_INIT=16'b0111000001110001;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_LC_11_10_0  (
            .in0(N__7515),
            .in1(N__8004),
            .in2(N__10324),
            .in3(N__7527),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_ENC_net ),
            .ce(),
            .sr(N__9025));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_11_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_11_11_0 .LUT_INIT=16'b0000101011111010;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_LC_11_11_0  (
            .in0(N__7946),
            .in1(_gnd_net_),
            .in2(N__10146),
            .in3(N__7932),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_11_2 .LUT_INIT=16'b0101000010100000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_11_2  (
            .in0(N__8002),
            .in1(_gnd_net_),
            .in2(N__10145),
            .in3(N__7513),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_11_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_11_4 .LUT_INIT=16'b0100000001010000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_11_4  (
            .in0(N__8003),
            .in1(N__7514),
            .in2(N__10144),
            .in3(N__7526),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_11_11_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_11_11_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__8153),
            .in2(_gnd_net_),
            .in3(N__7793),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_11_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_11_11_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_11_11_6  (
            .in0(N__7548),
            .in1(N__7841),
            .in2(N__7530),
            .in3(N__8015),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER6 ),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_11_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_11_7 .LUT_INIT=16'b0000000111011101;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_11_7  (
            .in0(N__7512),
            .in1(N__8001),
            .in2(N__7986),
            .in3(N__7945),
            .lcout(\U409_TRANSFER_ACK.TACK_OUTn_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_12_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_12_1 .LUT_INIT=16'b0011101010101010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_12_1  (
            .in0(N__7842),
            .in1(N__7926),
            .in2(N__7887),
            .in3(N__7877),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .ce(),
            .sr(N__9017));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_11_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_11_12_3 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_11_12_3  (
            .in0(N__7689),
            .in1(N__7830),
            .in2(N__7818),
            .in3(N__7794),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .ce(),
            .sr(N__9017));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_11_13_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_11_13_1 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_11_13_1  (
            .in0(N__7782),
            .in1(N__10094),
            .in2(N__7737),
            .in3(N__7713),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.LV_SPACE_LC_11_13_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.LV_SPACE_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.LV_SPACE_LC_11_13_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.LV_SPACE_LC_11_13_5  (
            .in0(N__7764),
            .in1(N__10295),
            .in2(N__7736),
            .in3(N__7712),
            .lcout(BUFENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_11_14_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_11_14_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_11_14_2  (
            .in0(N__8369),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8301),
            .lcout(\U409_TRANSFER_ACK.N_119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_1.C_ON=1'b0;
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_1.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8305),
            .lcout(GB_BUFFER_CLK40_IN_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_1_LC_12_7_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_1_LC_12_7_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_1_LC_12_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER60_1_LC_12_7_0  (
            .in0(_gnd_net_),
            .in1(N__8585),
            .in2(_gnd_net_),
            .in3(N__8421),
            .lcout(\U409_TICK.COUNTER60Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9606),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_7_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_7_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_7_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_9_LC_12_8_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_9_LC_12_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_9_LC_12_8_1 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \U409_TICK.COUNTER60_9_LC_12_8_1  (
            .in0(N__9369),
            .in1(N__8385),
            .in2(N__9336),
            .in3(N__9399),
            .lcout(\U409_TICK.COUNTER60Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9608),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_12_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_12_9_0 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_12_9_0  (
            .in0(N__8519),
            .in1(_gnd_net_),
            .in2(N__8562),
            .in3(N__8304),
            .lcout(\U409_TRANSFER_ACK.N_17_mux ),
            .ltout(\U409_TRANSFER_ACK.N_17_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_12_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_12_9_1 .LUT_INIT=16'b0001110100111111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_12_9_1  (
            .in0(N__8536),
            .in1(N__8057),
            .in2(N__8091),
            .in3(N__8548),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_12_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_12_9_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_12_9_2 .LUT_INIT=16'b0000010010001100;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_0_LC_12_9_2  (
            .in0(N__8033),
            .in1(N__10061),
            .in2(N__8088),
            .in3(N__8082),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_9_4 .LUT_INIT=16'b0001000000011111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_9_4  (
            .in0(N__8549),
            .in1(N__8537),
            .in2(N__8066),
            .in3(N__8076),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.N_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_9_5 .LUT_INIT=16'b0010101000001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_9_5  (
            .in0(N__10062),
            .in1(N__8032),
            .in2(N__8085),
            .in3(N__8064),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_12_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_12_9_6 .LUT_INIT=16'b0001111100010000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_12_9_6  (
            .in0(N__8550),
            .in1(N__8535),
            .in2(N__8067),
            .in3(N__8075),
            .lcout(\U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_12_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_12_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_12_9_7  (
            .in0(_gnd_net_),
            .in1(N__8558),
            .in2(_gnd_net_),
            .in3(N__8518),
            .lcout(\U409_TRANSFER_ACK.N_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_12_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_12_10_5 .LUT_INIT=16'b0101111100001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_LC_12_10_5  (
            .in0(N__8065),
            .in1(N__8040),
            .in2(N__8034),
            .in3(N__8016),
            .lcout(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__9018));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_12_11_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_12_11_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_12_11_1 .LUT_INIT=16'b0100010011111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_12_11_1  (
            .in0(N__8205),
            .in1(N__8154),
            .in2(_gnd_net_),
            .in3(N__8118),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .ce(),
            .sr(N__8773));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_12_12_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_12_12_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_12_12_0  (
            .in0(N__8964),
            .in1(N__8945),
            .in2(N__8192),
            .in3(N__8101),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_12_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_12_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__8924),
            .in2(_gnd_net_),
            .in3(N__8865),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_12_12_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_12_12_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_12_12_2  (
            .in0(N__8965),
            .in1(N__8946),
            .in2(N__8193),
            .in3(N__8102),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_12_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_12_12_3 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_12_12_3  (
            .in0(N__8893),
            .in1(N__8798),
            .in2(N__8142),
            .in3(N__8135),
            .lcout(\U409_TRANSFER_ACK.N_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_12_12_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_12_12_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_12_12_4  (
            .in0(N__8797),
            .in1(N__8892),
            .in2(N__8139),
            .in3(N__8127),
            .lcout(\U409_TRANSFER_ACK.N_87 ),
            .ltout(\U409_TRANSFER_ACK.N_87_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_3_LC_12_12_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_3_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_3_LC_12_12_5 .LUT_INIT=16'b0100000011111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_3_LC_12_12_5  (
            .in0(N__8370),
            .in1(N__8302),
            .in2(N__8121),
            .in3(N__8117),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_12_12_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_12_12_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_12_12_6 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_12_12_6  (
            .in0(N__8190),
            .in1(N__8103),
            .in2(N__8106),
            .in3(N__8982),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .ce(),
            .sr(N__8777));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_13_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_13_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_13_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_13_1  (
            .in0(N__8928),
            .in1(N__8899),
            .in2(_gnd_net_),
            .in3(N__8832),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__8766));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_13_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_13_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_13_2 .LUT_INIT=16'b0011111111000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(N__8927),
            .in2(N__8904),
            .in3(N__8868),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__8766));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_13_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_13_5 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_13_5 .LUT_INIT=16'b1101110000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_13_5  (
            .in0(N__8348),
            .in1(N__8898),
            .in2(N__8307),
            .in3(N__8204),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__8766));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_12_13_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_12_13_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_12_13_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_12_13_7  (
            .in0(N__8981),
            .in1(N__8191),
            .in2(_gnd_net_),
            .in3(N__8831),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__8766));
    defparam RESETn_ibuf_RNIM9SF_LC_12_15_2.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_15_2.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_15_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10027),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_5_LC_13_5_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_5_LC_13_5_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_5_LC_13_5_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_5_LC_13_5_0  (
            .in0(N__9736),
            .in1(N__9783),
            .in2(N__9690),
            .in3(N__9069),
            .lcout(\U409_TICK.COUNTER50Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9598),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_13_5_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_13_5_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER50_RNIUHF01_16_LC_13_5_1  (
            .in0(N__9054),
            .in1(N__8729),
            .in2(N__9093),
            .in3(N__9227),
            .lcout(\U409_TICK.TICK503_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_0_LC_13_5_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_0_LC_13_5_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_0_LC_13_5_4 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U409_TICK.COUNTER50_0_LC_13_5_4  (
            .in0(N__9735),
            .in1(N__9686),
            .in2(N__9128),
            .in3(N__9784),
            .lcout(\U409_TICK.COUNTER50Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9598),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_6_0 .C_ON=1'b1;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_6_0  (
            .in0(_gnd_net_),
            .in1(N__8419),
            .in2(N__8589),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_6_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_2_LC_13_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_2_LC_13_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_2_LC_13_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_2_LC_13_6_1  (
            .in0(_gnd_net_),
            .in1(N__8447),
            .in2(_gnd_net_),
            .in3(N__8157),
            .lcout(\U409_TICK.COUNTER60Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .clk(N__9600),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_3_LC_13_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_3_LC_13_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_3_LC_13_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_3_LC_13_6_2  (
            .in0(_gnd_net_),
            .in1(N__8603),
            .in2(_gnd_net_),
            .in3(N__8403),
            .lcout(\U409_TICK.COUNTER60Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .clk(N__9600),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_13_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_13_6_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_13_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_4_LC_13_6_3  (
            .in0(_gnd_net_),
            .in1(N__8643),
            .in2(_gnd_net_),
            .in3(N__8400),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_5_LC_13_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_5_LC_13_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_5_LC_13_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_5_LC_13_6_4  (
            .in0(_gnd_net_),
            .in1(N__8654),
            .in2(_gnd_net_),
            .in3(N__8397),
            .lcout(\U409_TICK.COUNTER60Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .clk(N__9600),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_13_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_13_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_13_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_6_LC_13_6_5  (
            .in0(_gnd_net_),
            .in1(N__9507),
            .in2(_gnd_net_),
            .in3(N__8394),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_7_LC_13_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_7_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_7_LC_13_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_7_LC_13_6_6  (
            .in0(_gnd_net_),
            .in1(N__8708),
            .in2(_gnd_net_),
            .in3(N__8391),
            .lcout(\U409_TICK.COUNTER60Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .clk(N__9600),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_13_6_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_13_6_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_13_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_8_LC_13_6_7  (
            .in0(_gnd_net_),
            .in1(N__9416),
            .in2(_gnd_net_),
            .in3(N__8388),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_13_7_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_13_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_9_LC_13_7_0  (
            .in0(_gnd_net_),
            .in1(N__9518),
            .in2(_gnd_net_),
            .in3(N__8379),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_13_7_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_10_LC_13_7_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_10_LC_13_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_10_LC_13_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_10_LC_13_7_1  (
            .in0(_gnd_net_),
            .in1(N__8696),
            .in2(_gnd_net_),
            .in3(N__8376),
            .lcout(\U409_TICK.COUNTER60Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .clk(N__9602),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_11_LC_13_7_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_11_LC_13_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_11_LC_13_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_11_LC_13_7_2  (
            .in0(_gnd_net_),
            .in1(N__8621),
            .in2(_gnd_net_),
            .in3(N__8373),
            .lcout(\U409_TICK.COUNTER60Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .clk(N__9602),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_12_LC_13_7_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_12_LC_13_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_12_LC_13_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_12_LC_13_7_3  (
            .in0(_gnd_net_),
            .in1(N__8462),
            .in2(_gnd_net_),
            .in3(N__8505),
            .lcout(\U409_TICK.COUNTER60Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .clk(N__9602),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_13_LC_13_7_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_13_LC_13_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_13_LC_13_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_13_LC_13_7_4  (
            .in0(_gnd_net_),
            .in1(N__8681),
            .in2(_gnd_net_),
            .in3(N__8502),
            .lcout(\U409_TICK.COUNTER60Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .clk(N__9602),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_13_7_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_13_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_14_LC_13_7_5  (
            .in0(_gnd_net_),
            .in1(N__9482),
            .in2(_gnd_net_),
            .in3(N__8499),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_13_7_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_13_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_15_LC_13_7_6  (
            .in0(_gnd_net_),
            .in1(N__8669),
            .in2(_gnd_net_),
            .in3(N__8496),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_16_LC_13_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_16_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_16_LC_13_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER60_16_LC_13_7_7  (
            .in0(_gnd_net_),
            .in1(N__8435),
            .in2(_gnd_net_),
            .in3(N__8493),
            .lcout(\U409_TICK.COUNTER60Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9602),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_6_LC_13_8_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_6_LC_13_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_6_LC_13_8_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_6_LC_13_8_0  (
            .in0(N__9395),
            .in1(N__9365),
            .in2(N__9334),
            .in3(N__8490),
            .lcout(\U409_TICK.COUNTER60Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9605),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_15_LC_13_8_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_15_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_15_LC_13_8_1 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_15_LC_13_8_1  (
            .in0(N__9363),
            .in1(N__9393),
            .in2(N__8481),
            .in3(N__9325),
            .lcout(\U409_TICK.COUNTER60Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9605),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_4_LC_13_8_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_4_LC_13_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_4_LC_13_8_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_4_LC_13_8_2  (
            .in0(N__9394),
            .in1(N__9364),
            .in2(N__9333),
            .in3(N__8472),
            .lcout(\U409_TICK.COUNTER60Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9605),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_8_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_8_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_8_3  (
            .in0(N__8463),
            .in1(N__8451),
            .in2(N__8436),
            .in3(N__8420),
            .lcout(\U409_TICK.TICK603_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_13_8_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_13_8_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_TICK.COUNTER60_RNI2USG_10_LC_13_8_4  (
            .in0(N__8712),
            .in1(N__8697),
            .in2(N__8685),
            .in3(N__8670),
            .lcout(\U409_TICK.TICK603_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_13_8_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_13_8_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_TICK.COUNTER60_RNIHJU51_4_LC_13_8_5  (
            .in0(N__8658),
            .in1(N__8642),
            .in2(_gnd_net_),
            .in3(N__8583),
            .lcout(),
            .ltout(\U409_TICK.TICK603_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_13_8_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_13_8_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER60_RNI335G2_11_LC_13_8_6  (
            .in0(N__8628),
            .in1(N__8622),
            .in2(N__8610),
            .in3(N__8607),
            .lcout(\U409_TICK.TICK603_14 ),
            .ltout(\U409_TICK.TICK603_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_0_LC_13_8_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_0_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_0_LC_13_8_7 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \U409_TICK.COUNTER60_0_LC_13_8_7  (
            .in0(N__9362),
            .in1(N__9318),
            .in2(N__8592),
            .in3(N__8584),
            .lcout(\U409_TICK.COUNTER60Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9605),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_13_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_13_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_1_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8520),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .ce(),
            .sr(N__9027));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_13_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_13_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_13_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8538),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .ce(),
            .sr(N__9027));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_13_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_13_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_13_9_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_13_9_3  (
            .in0(_gnd_net_),
            .in1(N__10060),
            .in2(_gnd_net_),
            .in3(N__9974),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .ce(),
            .sr(N__9027));
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_13_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_13_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_13_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_0_LC_13_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9200),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .ce(),
            .sr(N__9027));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_13_13_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_13_13_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_13_13_0  (
            .in0(N__8966),
            .in1(N__8866),
            .in2(N__8805),
            .in3(N__8947),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_13_13_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_13_13_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(N__8894),
            .in2(N__8985),
            .in3(N__8925),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_13_13_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_13_13_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_13_13_3  (
            .in0(N__8948),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8802),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_13_13_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_13_13_4 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_13_13_4 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_13_13_4  (
            .in0(N__8967),
            .in1(N__8834),
            .in2(N__8970),
            .in3(N__8846),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__8778));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_13_13_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_13_13_5 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_13_13_5 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_13_13_5  (
            .in0(N__8949),
            .in1(N__8804),
            .in2(N__8847),
            .in3(N__8833),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__8778));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_13_13_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_13_13_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_13_13_6  (
            .in0(N__8926),
            .in1(_gnd_net_),
            .in2(N__8903),
            .in3(N__8867),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_13_13_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_13_13_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_13_13_7 .LUT_INIT=16'b0001010000010100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_13_13_7  (
            .in0(N__8835),
            .in1(N__8803),
            .in2(N__8808),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__8778));
    defparam \U409_TICK.COUNTER50_1_LC_14_4_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_1_LC_14_4_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_1_LC_14_4_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER50_1_LC_14_4_0  (
            .in0(_gnd_net_),
            .in1(N__9120),
            .in2(_gnd_net_),
            .in3(N__8730),
            .lcout(\U409_TICK.COUNTER50Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9599),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_5_0 .C_ON=1'b1;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_5_0  (
            .in0(_gnd_net_),
            .in1(N__8728),
            .in2(N__9124),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_5_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_2_LC_14_5_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_2_LC_14_5_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_2_LC_14_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_2_LC_14_5_1  (
            .in0(_gnd_net_),
            .in1(N__9089),
            .in2(_gnd_net_),
            .in3(N__9078),
            .lcout(\U409_TICK.COUNTER50Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .clk(N__9601),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_3_LC_14_5_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_3_LC_14_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_3_LC_14_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_3_LC_14_5_2  (
            .in0(_gnd_net_),
            .in1(N__9140),
            .in2(_gnd_net_),
            .in3(N__9075),
            .lcout(\U409_TICK.COUNTER50Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .clk(N__9601),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_4_LC_14_5_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_4_LC_14_5_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_4_LC_14_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_4_LC_14_5_3  (
            .in0(_gnd_net_),
            .in1(N__9851),
            .in2(_gnd_net_),
            .in3(N__9072),
            .lcout(\U409_TICK.COUNTER50Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .clk(N__9601),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_14_5_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_14_5_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_5_LC_14_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9164),
            .in3(N__9063),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_14_5_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_14_5_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_14_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_6_LC_14_5_5  (
            .in0(_gnd_net_),
            .in1(N__9878),
            .in2(_gnd_net_),
            .in3(N__9060),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_7_LC_14_5_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_7_LC_14_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_7_LC_14_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_7_LC_14_5_6  (
            .in0(_gnd_net_),
            .in1(N__9866),
            .in2(_gnd_net_),
            .in3(N__9057),
            .lcout(\U409_TICK.COUNTER50Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .clk(N__9601),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_8_LC_14_5_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_8_LC_14_5_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_8_LC_14_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_8_LC_14_5_7  (
            .in0(_gnd_net_),
            .in1(N__9053),
            .in2(_gnd_net_),
            .in3(N__9042),
            .lcout(\U409_TICK.COUNTER50Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .clk(N__9601),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_14_6_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_14_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_9_LC_14_6_0  (
            .in0(_gnd_net_),
            .in1(N__9263),
            .in2(_gnd_net_),
            .in3(N__9039),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_14_6_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_10_LC_14_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_10_LC_14_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_10_LC_14_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_10_LC_14_6_1  (
            .in0(_gnd_net_),
            .in1(N__9560),
            .in2(_gnd_net_),
            .in3(N__9036),
            .lcout(\U409_TICK.COUNTER50Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .clk(N__9603),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_14_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_14_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_11_LC_14_6_2  (
            .in0(_gnd_net_),
            .in1(N__9620),
            .in2(_gnd_net_),
            .in3(N__9246),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_12_LC_14_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_12_LC_14_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_12_LC_14_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_12_LC_14_6_3  (
            .in0(_gnd_net_),
            .in1(N__9533),
            .in2(_gnd_net_),
            .in3(N__9243),
            .lcout(\U409_TICK.COUNTER50Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .clk(N__9603),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_14_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_14_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_13_LC_14_6_4  (
            .in0(_gnd_net_),
            .in1(N__9833),
            .in2(_gnd_net_),
            .in3(N__9240),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_14_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_14_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_14_LC_14_6_5  (
            .in0(_gnd_net_),
            .in1(N__9797),
            .in2(_gnd_net_),
            .in3(N__9237),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_14_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_14_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_15_LC_14_6_6  (
            .in0(_gnd_net_),
            .in1(N__9815),
            .in2(_gnd_net_),
            .in3(N__9234),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_16_LC_14_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_16_LC_14_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_16_LC_14_6_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER50_16_LC_14_6_7  (
            .in0(_gnd_net_),
            .in1(N__9228),
            .in2(_gnd_net_),
            .in3(N__9231),
            .lcout(\U409_TICK.COUNTER50Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9603),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_14_7_0 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_14_7_0 .LUT_INIT=16'b0000000000011000;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_1_LC_14_7_0  (
            .in0(N__10587),
            .in1(N__10473),
            .in2(N__9199),
            .in3(N__10449),
            .lcout(),
            .ltout(\U409_CIA.CLK_CIA_r_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_LC_14_7_1 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_LC_14_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CLK_CIA_LC_14_7_1 .LUT_INIT=16'b1010101001101010;
    LogicCell40 \U409_CIA.CLK_CIA_LC_14_7_1  (
            .in0(N__9192),
            .in1(N__9567),
            .in2(N__9216),
            .in3(N__10423),
            .lcout(CLK_CIA_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10491),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_14_7_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_14_7_5 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \U409_TICK.COUNTER50_RNID6CP_3_LC_14_7_5  (
            .in0(N__9168),
            .in1(_gnd_net_),
            .in2(N__9147),
            .in3(N__9129),
            .lcout(),
            .ltout(\U409_TICK.TICK503_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_14_7_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_14_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_14_7_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_TICK.COUNTER50_RNITU182_10_LC_14_7_6  (
            .in0(N__9561),
            .in1(N__9549),
            .in2(N__9537),
            .in3(N__9534),
            .lcout(\U409_TICK.TICK503_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_14_8_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_14_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNICDC71_14_LC_14_8_1  (
            .in0(N__9522),
            .in1(N__9506),
            .in2(N__9417),
            .in3(N__9483),
            .lcout(\U409_TICK.TICK603_9 ),
            .ltout(\U409_TICK.TICK603_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_14_LC_14_8_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_14_LC_14_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_14_LC_14_8_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_14_LC_14_8_2  (
            .in0(N__9366),
            .in1(N__9396),
            .in2(N__9492),
            .in3(N__9489),
            .lcout(\U409_TICK.COUNTER60Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9609),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_9_LC_14_8_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_9_LC_14_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_9_LC_14_8_3 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_9_LC_14_8_3  (
            .in0(N__9684),
            .in1(N__9734),
            .in2(N__9471),
            .in3(N__9786),
            .lcout(\U409_TICK.COUNTER50Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9609),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK50_LC_14_8_5 .C_ON=1'b0;
    defparam \U409_TICK.TICK50_LC_14_8_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK50_LC_14_8_5 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK50_LC_14_8_5  (
            .in0(N__9685),
            .in1(N__9443),
            .in2(N__9741),
            .in3(N__9785),
            .lcout(TICK50_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9609),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_8_LC_14_8_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_8_LC_14_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_8_LC_14_8_6 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_8_LC_14_8_6  (
            .in0(N__9367),
            .in1(N__9397),
            .in2(N__9432),
            .in3(N__9329),
            .lcout(\U409_TICK.COUNTER60Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9609),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK60_LC_14_8_7 .C_ON=1'b0;
    defparam \U409_TICK.TICK60_LC_14_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK60_LC_14_8_7 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \U409_TICK.TICK60_LC_14_8_7  (
            .in0(N__9398),
            .in1(N__9368),
            .in2(N__9335),
            .in3(N__9275),
            .lcout(TICK60_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9609),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_15_5_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_15_5_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_15_5_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNIH14V_11_LC_15_5_1  (
            .in0(N__9621),
            .in1(N__9264),
            .in2(N__9882),
            .in3(N__9834),
            .lcout(\U409_TICK.TICK503_9 ),
            .ltout(\U409_TICK.TICK503_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_6_LC_15_5_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_6_LC_15_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_6_LC_15_5_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_6_LC_15_5_2  (
            .in0(N__9778),
            .in1(N__9740),
            .in2(N__9891),
            .in3(N__9888),
            .lcout(\U409_TICK.COUNTER50Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9604),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_15_5_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_15_5_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_15_5_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNII24V_14_LC_15_5_3  (
            .in0(N__9798),
            .in1(N__9867),
            .in2(N__9855),
            .in3(N__9816),
            .lcout(\U409_TICK.TICK503_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_13_LC_15_6_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_13_LC_15_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_13_LC_15_6_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_13_LC_15_6_4  (
            .in0(N__9730),
            .in1(N__9781),
            .in2(N__9682),
            .in3(N__9840),
            .lcout(\U409_TICK.COUNTER50Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9607),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_15_LC_15_6_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_15_LC_15_6_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_15_LC_15_6_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_15_LC_15_6_5  (
            .in0(N__9780),
            .in1(N__9733),
            .in2(N__9681),
            .in3(N__9822),
            .lcout(\U409_TICK.COUNTER50Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9607),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_14_LC_15_6_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_14_LC_15_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_14_LC_15_6_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_14_LC_15_6_6  (
            .in0(N__9731),
            .in1(N__9782),
            .in2(N__9683),
            .in3(N__9804),
            .lcout(\U409_TICK.COUNTER50Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9607),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_11_LC_15_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_11_LC_15_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_11_LC_15_6_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_11_LC_15_6_7  (
            .in0(N__9779),
            .in1(N__9732),
            .in2(N__9680),
            .in3(N__9627),
            .lcout(\U409_TICK.COUNTER50Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9607),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_15_7_0 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_15_7_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_0_LC_15_7_0  (
            .in0(N__10392),
            .in1(N__10546),
            .in2(N__10518),
            .in3(N__9917),
            .lcout(\U409_CIA.CLK_CIA6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_15_7_1 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_15_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_15_7_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_1_LC_15_7_1  (
            .in0(N__9919),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10393),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10489),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_15_7_2 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_15_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_15_7_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_15_7_2  (
            .in0(N__10547),
            .in1(N__10582),
            .in2(N__10517),
            .in3(N__9918),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_3 ),
            .ltout(\U409_CIA.CIA_CLK_COUNT11_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_15_7_3 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_15_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_15_7_3 .LUT_INIT=16'b0001010100101010;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_3_LC_15_7_3  (
            .in0(N__10472),
            .in1(N__9942),
            .in2(N__9945),
            .in3(N__10596),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10489),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_15_7_5 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_15_7_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_15_7_5  (
            .in0(N__10471),
            .in1(N__10445),
            .in2(N__10425),
            .in3(N__10391),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_2_0 ),
            .ltout(\U409_CIA.CIA_CLK_COUNT11_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_15_7_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_15_7_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_15_7_6 .LUT_INIT=16'b0001001101001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_5_LC_15_7_6  (
            .in0(N__9936),
            .in1(N__10422),
            .in2(N__9930),
            .in3(N__10557),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10489),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_1_LC_16_6_0 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_1_LC_16_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_1_LC_16_6_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_CIA.VMA_RNO_1_LC_16_6_0  (
            .in0(_gnd_net_),
            .in1(N__10515),
            .in2(_gnd_net_),
            .in3(N__10545),
            .lcout(),
            .ltout(\U409_CIA.CLK_CIA6_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_0_LC_16_6_1 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_0_LC_16_6_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_0_LC_16_6_1 .LUT_INIT=16'b0100000010000000;
    LogicCell40 \U409_CIA.VMA_RNO_0_LC_16_6_1  (
            .in0(N__10583),
            .in1(N__10365),
            .in2(N__9927),
            .in3(N__9920),
            .lcout(),
            .ltout(\U409_CIA.VMA_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_LC_16_6_2 .C_ON=1'b0;
    defparam \U409_CIA.VMA_LC_16_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.VMA_LC_16_6_2 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \U409_CIA.VMA_LC_16_6_2  (
            .in0(N__9921),
            .in1(N__10248),
            .in2(N__9924),
            .in3(N__9961),
            .lcout(\U409_CIA.VMAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10490),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_16_6_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_16_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_16_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_0_LC_16_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10394),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10490),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_16_7_0 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_16_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_16_7_0  (
            .in0(_gnd_net_),
            .in1(N__9916),
            .in2(N__10395),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_7_0_),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_16_7_1 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_16_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_16_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_2_LC_16_7_1  (
            .in0(_gnd_net_),
            .in1(N__10443),
            .in2(_gnd_net_),
            .in3(N__9894),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .clk(N__10488),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_16_7_2 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_16_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_16_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_16_7_2  (
            .in0(_gnd_net_),
            .in1(N__10469),
            .in2(_gnd_net_),
            .in3(N__10590),
            .lcout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_16_7_3 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_16_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_16_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_4_LC_16_7_3  (
            .in0(_gnd_net_),
            .in1(N__10581),
            .in2(_gnd_net_),
            .in3(N__10560),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .clk(N__10488),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_16_7_4 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_16_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_16_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_16_7_4  (
            .in0(_gnd_net_),
            .in1(N__10418),
            .in2(_gnd_net_),
            .in3(N__10551),
            .lcout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_16_7_5 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_16_7_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_16_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_6_LC_16_7_5  (
            .in0(_gnd_net_),
            .in1(N__10548),
            .in2(_gnd_net_),
            .in3(N__10524),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ),
            .clk(N__10488),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_16_7_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_16_7_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_16_7_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_7_LC_16_7_6  (
            .in0(_gnd_net_),
            .in1(N__10516),
            .in2(_gnd_net_),
            .in3(N__10521),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10488),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_2_LC_16_7_7 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_2_LC_16_7_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_2_LC_16_7_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_CIA.VMA_RNO_2_LC_16_7_7  (
            .in0(N__10470),
            .in1(N__10444),
            .in2(N__10424),
            .in3(N__10390),
            .lcout(\U409_CIA.un1_CIA_CLK_COUNT_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_16_13_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_16_13_4 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_16_13_4  (
            .in0(N__10337),
            .in1(N__10299),
            .in2(_gnd_net_),
            .in3(N__10238),
            .lcout(TCIn_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNI692L_0_LC_22_3_4 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNI692L_0_LC_22_3_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNI692L_0_LC_22_3_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_CIA.VMA_RNI692L_0_LC_22_3_4  (
            .in0(N__10005),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9975),
            .lcout(CIA_ENABLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_24_3_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_24_3_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_24_3_1 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_24_3_1  (
            .in0(N__10709),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10658),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS0n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_24_3_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_24_3_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_24_3_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_24_3_6  (
            .in0(N__10659),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10640),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS1n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U409_TOP

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     May 13 2025 19:08:48

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    DA : out std_logic_vector(2 downto 0);
    A : in std_logic_vector(20 downto 0);
    DBRn : in std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    TCIn : out std_logic;
    TBIn : out std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__12615\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12146\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12037\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \A_c_14\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.N_340\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_297_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_196_cascade_\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_95_i_a2_i_0\ : std_logic;
signal \U712_CHIP_RAM.N_556_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_202\ : std_logic;
signal \U712_CHIP_RAM.N_388_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_i_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto7_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lt7\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_417_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_1\ : std_logic;
signal \U712_CHIP_RAM.N_206\ : std_logic;
signal \U712_CHIP_RAM.N_457\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_i_1\ : std_logic;
signal \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\ : std_logic;
signal \LATCH_CLK_c\ : std_logic;
signal \TSn_c\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.N_414\ : std_logic;
signal \U712_CYCLE_TERM.N_452_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_312\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ1Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.START_RSTZ0\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \RASn_c\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\ : std_logic;
signal \U712_CHIP_RAM.N_346\ : std_logic;
signal \U712_CHIP_RAM.N_388\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA25_0_i_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_10_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_445\ : std_logic;
signal \U712_CHIP_RAM.N_208\ : std_logic;
signal \U712_CHIP_RAM.N_303\ : std_logic;
signal \U712_CHIP_RAM.N_443_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_204\ : std_logic;
signal \U712_CHIP_RAM.N_463_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_439\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_0_a2_1_0\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_cascade_\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_360\ : std_logic;
signal \U712_CHIP_RAM.N_418\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_5_0\ : std_logic;
signal \U712_REG_SM.N_400_cascade_\ : std_logic;
signal \U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_405\ : std_logic;
signal \bfn_10_12_0_\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \DBR_SYNC_i_1\ : std_logic;
signal \U712_REG_SM.N_307_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_3\ : std_logic;
signal \REGENn_c\ : std_logic;
signal \U712_REG_SM.REGENn_e_1\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.WRITE_CYCLEZ0\ : std_logic;
signal \A_c_12\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_551\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_10_0_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.N_555_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER16\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER16_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_556\ : std_logic;
signal \U712_CHIP_RAM.N_302\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER19\ : std_logic;
signal \U712_CHIP_RAM.N_355_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_389\ : std_logic;
signal \U712_CHIP_RAM.N_301\ : std_logic;
signal \U712_CHIP_RAM.N_289\ : std_logic;
signal \U712_CHIP_RAM.N_356\ : std_logic;
signal \U712_CHIP_RAM.N_356_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_448\ : std_logic;
signal \U712_CHIP_RAM.N_288_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_473\ : std_logic;
signal \U712_CHIP_RAM.N_473_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_i_1_0\ : std_logic;
signal \U712_CHIP_RAM.N_362\ : std_logic;
signal \U712_CHIP_RAM.N_463\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_0\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\ : std_logic;
signal \U712_REG_SM.N_306_cascade_\ : std_logic;
signal \U712_REG_SM.N_399_cascade_\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_5_iv_0_0\ : std_logic;
signal \U712_REG_SM.N_311\ : std_logic;
signal \U712_REG_SM.N_353_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_322\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_REG_SM.STATE_COUNTsr_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_7\ : std_logic;
signal \U712_REG_SM.N_307\ : std_logic;
signal \U712_REG_SM.N_553\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_4\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_5\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_6\ : std_logic;
signal \N_130_i\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0\ : std_logic;
signal \U712_CHIP_RAM.N_294_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_288\ : std_logic;
signal \U712_CHIP_RAM.N_469_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_557\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.N_555\ : std_logic;
signal \U712_CHIP_RAM.N_309_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_387\ : std_logic;
signal \U712_CHIP_RAM.N_200_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_309\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.N_285\ : std_logic;
signal \U712_CHIP_RAM.N_285_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_293\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_a2_0_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.N_200\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_2\ : std_logic;
signal \U712_BYTE_ENABLE.N_451\ : std_logic;
signal \N_211_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_410_cascade_\ : std_logic;
signal \N_148_i\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_a2Z0Z_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_8\ : std_logic;
signal \U712_REG_SM.N_95_cascade_\ : std_logic;
signal \U712_REG_SM.N_432\ : std_logic;
signal \LDSn_c\ : std_logic;
signal \U712_REG_SM.N_95\ : std_logic;
signal \UDSn_c\ : std_logic;
signal \U712_REG_SM.N_433\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.N_297\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\ : std_logic;
signal \U712_BYTE_ENABLE.N_409\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.N_95_0\ : std_logic;
signal \LLBEn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \CASn_c\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \N_146_i\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_406\ : std_logic;
signal \U712_BYTE_ENABLE.N_284_i\ : std_logic;
signal \N_374_i\ : std_logic;
signal \N_373_i\ : std_logic;
signal \A_c_1\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \UMBEn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_i_0_9\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA25_0_i_0\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \U712_BYTE_ENABLE.N_411\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \N_150_i\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_0\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \N_136_i\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \RnW_c\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \DMA_WRITE_CYCLE\ : std_logic;
signal \N_357\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \DA_wire\ : std_logic_vector(2 downto 0);
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    TBIn <= \TBIn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    ASn <= \ASn_wire\;
    DA <= \DA_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    TCIn <= \TCIn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__4376\,
            RESETB => \N__6917\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12615\,
            DIN => \N__12614\,
            DOUT => \N__12613\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12615\,
            PADOUT => \N__12614\,
            PADIN => \N__12613\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11093\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12606\,
            DIN => \N__12605\,
            DOUT => \N__12604\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12606\,
            PADOUT => \N__12605\,
            PADIN => \N__12604\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12597\,
            DIN => \N__12596\,
            DOUT => \N__12595\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12597\,
            PADOUT => \N__12596\,
            PADIN => \N__12595\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9083\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12588\,
            DIN => \N__12587\,
            DOUT => \N__12586\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12588\,
            PADOUT => \N__12587\,
            PADIN => \N__12586\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11651\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12579\,
            DIN => \N__12578\,
            DOUT => \N__12577\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12579\,
            PADOUT => \N__12578\,
            PADIN => \N__12577\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12570\,
            DIN => \N__12569\,
            DOUT => \N__12568\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12570\,
            PADOUT => \N__12569\,
            PADIN => \N__12568\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12561\,
            DIN => \N__12560\,
            DOUT => \N__12559\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12561\,
            PADOUT => \N__12560\,
            PADIN => \N__12559\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12552\,
            DIN => \N__12551\,
            DOUT => \N__12550\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12552\,
            PADOUT => \N__12551\,
            PADIN => \N__12550\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12543\,
            DIN => \N__12542\,
            DOUT => \N__12541\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12543\,
            PADOUT => \N__12542\,
            PADIN => \N__12541\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12534\,
            DIN => \N__12533\,
            DOUT => \N__12532\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12534\,
            PADOUT => \N__12533\,
            PADIN => \N__12532\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12525\,
            DIN => \N__12524\,
            DOUT => \N__12523\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12525\,
            PADOUT => \N__12524\,
            PADIN => \N__12523\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12516\,
            DIN => \N__12515\,
            DOUT => \N__12514\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12516\,
            PADOUT => \N__12515\,
            PADIN => \N__12514\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4673\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12507\,
            DIN => \N__12506\,
            DOUT => \N__12505\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12507\,
            PADOUT => \N__12506\,
            PADIN => \N__12505\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11633\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12498\,
            DIN => \N__12497\,
            DOUT => \N__12496\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12498\,
            PADOUT => \N__12497\,
            PADIN => \N__12496\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12489\,
            DIN => \N__12488\,
            DOUT => \N__12487\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12489\,
            PADOUT => \N__12488\,
            PADIN => \N__12487\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12480\,
            DIN => \N__12479\,
            DOUT => \N__12478\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12480\,
            PADOUT => \N__12479\,
            PADIN => \N__12478\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12471\,
            DIN => \N__12470\,
            DOUT => \N__12469\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12471\,
            PADOUT => \N__12470\,
            PADIN => \N__12469\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4406\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12462\,
            DIN => \N__12461\,
            DOUT => \N__12460\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12462\,
            PADOUT => \N__12461\,
            PADIN => \N__12460\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12453\,
            DIN => \N__12452\,
            DOUT => \N__12451\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12453\,
            PADOUT => \N__12452\,
            PADIN => \N__12451\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12444\,
            DIN => \N__12443\,
            DOUT => \N__12442\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12444\,
            PADOUT => \N__12443\,
            PADIN => \N__12442\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5354\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12435\,
            DIN => \N__12434\,
            DOUT => \N__12433\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12435\,
            PADOUT => \N__12434\,
            PADIN => \N__12433\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12426\,
            DIN => \N__12425\,
            DOUT => \N__12424\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12426\,
            PADOUT => \N__12425\,
            PADIN => \N__12424\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5393\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12417\,
            DIN => \N__12416\,
            DOUT => \N__12415\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12417\,
            PADOUT => \N__12416\,
            PADIN => \N__12415\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12408\,
            DIN => \N__12407\,
            DOUT => \N__12406\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12408\,
            PADOUT => \N__12407\,
            PADIN => \N__12406\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9242\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12399\,
            DIN => \N__12398\,
            DOUT => \N__12397\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12399\,
            PADOUT => \N__12398\,
            PADIN => \N__12397\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4486\,
            DIN0 => OPEN,
            DOUT0 => \N__5248\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12390\,
            DIN => \N__12389\,
            DOUT => \N__12388\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12390\,
            PADOUT => \N__12389\,
            PADIN => \N__12388\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12381\,
            DIN => \N__12380\,
            DOUT => \N__12379\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12381\,
            PADOUT => \N__12380\,
            PADIN => \N__12379\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12372\,
            DIN => \N__12371\,
            DOUT => \N__12370\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12372\,
            PADOUT => \N__12371\,
            PADIN => \N__12370\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12363\,
            DIN => \N__12362\,
            DOUT => \N__12361\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12363\,
            PADOUT => \N__12362\,
            PADIN => \N__12361\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12354\,
            DIN => \N__12353\,
            DOUT => \N__12352\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12354\,
            PADOUT => \N__12353\,
            PADIN => \N__12352\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12345\,
            DIN => \N__12344\,
            DOUT => \N__12343\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12345\,
            PADOUT => \N__12344\,
            PADIN => \N__12343\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6647\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12336\,
            DIN => \N__12335\,
            DOUT => \N__12334\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12336\,
            PADOUT => \N__12335\,
            PADIN => \N__12334\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12327\,
            DIN => \N__12326\,
            DOUT => \N__12325\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12327\,
            PADOUT => \N__12326\,
            PADIN => \N__12325\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12318\,
            DIN => \N__12317\,
            DOUT => \N__12316\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12318\,
            PADOUT => \N__12317\,
            PADIN => \N__12316\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12309\,
            DIN => \N__12308\,
            DOUT => \N__12307\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12309\,
            PADOUT => \N__12308\,
            PADIN => \N__12307\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12300\,
            DIN => \N__12299\,
            DOUT => \N__12298\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12300\,
            PADOUT => \N__12299\,
            PADIN => \N__12298\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12291\,
            DIN => \N__12290\,
            DOUT => \N__12289\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12291\,
            PADOUT => \N__12290\,
            PADIN => \N__12289\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5372\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12282\,
            DIN => \N__12281\,
            DOUT => \N__12280\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12282\,
            PADOUT => \N__12281\,
            PADIN => \N__12280\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12273\,
            DIN => \N__12272\,
            DOUT => \N__12271\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12273\,
            PADOUT => \N__12272\,
            PADIN => \N__12271\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12264\,
            DIN => \N__12263\,
            DOUT => \N__12262\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12264\,
            PADOUT => \N__12263\,
            PADIN => \N__12262\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9266\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12255\,
            DIN => \N__12254\,
            DOUT => \N__12253\,
            PACKAGEPIN => \DA_wire\(0)
        );

    \DA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12255\,
            PADOUT => \N__12254\,
            PADIN => \N__12253\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5318\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12246\,
            DIN => \N__12245\,
            DOUT => \N__12244\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12246\,
            PADOUT => \N__12245\,
            PADIN => \N__12244\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12237\,
            DIN => \N__12236\,
            DOUT => \N__12235\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12237\,
            PADOUT => \N__12236\,
            PADIN => \N__12235\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5342\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12228\,
            DIN => \N__12227\,
            DOUT => \N__12226\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12228\,
            PADOUT => \N__12227\,
            PADIN => \N__12226\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8597\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12219\,
            DIN => \N__12218\,
            DOUT => \N__12217\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12219\,
            PADOUT => \N__12218\,
            PADIN => \N__12217\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6137\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12210\,
            DIN => \N__12209\,
            DOUT => \N__12208\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12210\,
            PADOUT => \N__12209\,
            PADIN => \N__12208\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12201\,
            DIN => \N__12200\,
            DOUT => \N__12199\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12201\,
            PADOUT => \N__12200\,
            PADIN => \N__12199\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12192\,
            DIN => \N__12191\,
            DOUT => \N__12190\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12192\,
            PADOUT => \N__12191\,
            PADIN => \N__12190\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11021\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12183\,
            DIN => \N__12182\,
            DOUT => \N__12181\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12183\,
            PADOUT => \N__12182\,
            PADIN => \N__12181\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4487\,
            DIN0 => OPEN,
            DOUT0 => \N__5252\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12174\,
            DIN => \N__12173\,
            DOUT => \N__12172\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12174\,
            PADOUT => \N__12173\,
            PADIN => \N__12172\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6860\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12165\,
            DIN => \N__12164\,
            DOUT => \N__12163\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12165\,
            PADOUT => \N__12164\,
            PADIN => \N__12163\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6407\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12156\,
            DIN => \N__12155\,
            DOUT => \N__12154\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12156\,
            PADOUT => \N__12155\,
            PADIN => \N__12154\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8369\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12147\,
            DIN => \N__12146\,
            DOUT => \N__12145\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12147\,
            PADOUT => \N__12146\,
            PADIN => \N__12145\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12138\,
            DIN => \N__12137\,
            DOUT => \N__12136\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12138\,
            PADOUT => \N__12137\,
            PADIN => \N__12136\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12129\,
            DIN => \N__12128\,
            DOUT => \N__12127\,
            PACKAGEPIN => \DA_wire\(2)
        );

    \DA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12129\,
            PADOUT => \N__12128\,
            PADIN => \N__12127\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6047\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12120\,
            DIN => \N__12119\,
            DOUT => \N__12118\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12120\,
            PADOUT => \N__12119\,
            PADIN => \N__12118\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12111\,
            DIN => \N__12110\,
            DOUT => \N__12109\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12111\,
            PADOUT => \N__12110\,
            PADIN => \N__12109\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12102\,
            DIN => \N__12101\,
            DOUT => \N__12100\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12102\,
            PADOUT => \N__12101\,
            PADIN => \N__12100\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4556\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12093\,
            DIN => \N__12092\,
            DOUT => \N__12091\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12093\,
            PADOUT => \N__12092\,
            PADIN => \N__12091\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9413\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12084\,
            DIN => \N__12083\,
            DOUT => \N__12082\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12084\,
            PADOUT => \N__12083\,
            PADIN => \N__12082\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12075\,
            DIN => \N__12074\,
            DOUT => \N__12073\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12075\,
            PADOUT => \N__12074\,
            PADIN => \N__12073\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9551\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12066\,
            DIN => \N__12065\,
            DOUT => \N__12064\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12066\,
            PADOUT => \N__12065\,
            PADIN => \N__12064\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4461\,
            DIN0 => OPEN,
            DOUT0 => \N__5241\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12057\,
            DIN => \N__12056\,
            DOUT => \N__12055\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12057\,
            PADOUT => \N__12056\,
            PADIN => \N__12055\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5330\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12048\,
            DIN => \N__12047\,
            DOUT => \N__12046\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12048\,
            PADOUT => \N__12047\,
            PADIN => \N__12046\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12039\,
            DIN => \N__12038\,
            DOUT => \N__12037\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12039\,
            PADOUT => \N__12038\,
            PADIN => \N__12037\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12030\,
            DIN => \N__12029\,
            DOUT => \N__12028\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12030\,
            PADOUT => \N__12029\,
            PADIN => \N__12028\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4652\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12021\,
            DIN => \N__12020\,
            DOUT => \N__12019\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12021\,
            PADOUT => \N__12020\,
            PADIN => \N__12019\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12012\,
            DIN => \N__12011\,
            DOUT => \N__12010\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12012\,
            PADOUT => \N__12011\,
            PADIN => \N__12010\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12003\,
            DIN => \N__12002\,
            DOUT => \N__12001\,
            PACKAGEPIN => \DA_wire\(1)
        );

    \DA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12003\,
            PADOUT => \N__12002\,
            PADIN => \N__12001\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4730\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11994\,
            DIN => \N__11993\,
            DOUT => \N__11992\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11994\,
            PADOUT => \N__11993\,
            PADIN => \N__11992\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11985\,
            DIN => \N__11984\,
            DOUT => \N__11983\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11985\,
            PADOUT => \N__11984\,
            PADIN => \N__11983\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11976\,
            DIN => \N__11975\,
            DOUT => \N__11974\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11976\,
            PADOUT => \N__11975\,
            PADIN => \N__11974\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4529\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11967\,
            DIN => \N__11966\,
            DOUT => \N__11965\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11967\,
            PADOUT => \N__11966\,
            PADIN => \N__11965\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8672\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11958\,
            DIN => \N__11957\,
            DOUT => \N__11956\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11958\,
            PADOUT => \N__11957\,
            PADIN => \N__11956\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11288\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11949\,
            DIN => \N__11948\,
            DOUT => \N__11947\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11949\,
            PADOUT => \N__11948\,
            PADIN => \N__11947\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5717\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11940\,
            DIN => \N__11939\,
            DOUT => \N__11938\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11940\,
            PADOUT => \N__11939\,
            PADIN => \N__11938\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11931\,
            DIN => \N__11930\,
            DOUT => \N__11929\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11931\,
            PADOUT => \N__11930\,
            PADIN => \N__11929\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11922\,
            DIN => \N__11921\,
            DOUT => \N__11920\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11922\,
            PADOUT => \N__11921\,
            PADIN => \N__11920\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8459\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11913\,
            DIN => \N__11912\,
            DOUT => \N__11911\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11913\,
            PADOUT => \N__11912\,
            PADIN => \N__11911\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11904\,
            DIN => \N__11903\,
            DOUT => \N__11902\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11904\,
            PADOUT => \N__11903\,
            PADIN => \N__11902\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11895\,
            DIN => \N__11894\,
            DOUT => \N__11893\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11895\,
            PADOUT => \N__11894\,
            PADIN => \N__11893\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5048\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11886\,
            DIN => \N__11885\,
            DOUT => \N__11884\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11886\,
            PADOUT => \N__11885\,
            PADIN => \N__11884\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8174\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11877\,
            DIN => \N__11876\,
            DOUT => \N__11875\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11877\,
            PADOUT => \N__11876\,
            PADIN => \N__11875\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9482\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11868\,
            DIN => \N__11867\,
            DOUT => \N__11866\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11868\,
            PADOUT => \N__11867\,
            PADIN => \N__11866\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11859\,
            DIN => \N__11858\,
            DOUT => \N__11857\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11859\,
            PADOUT => \N__11858\,
            PADIN => \N__11857\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9471\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11850\,
            DIN => \N__11849\,
            DOUT => \N__11848\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11850\,
            PADOUT => \N__11849\,
            PADIN => \N__11848\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4430\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11841\,
            DIN => \N__11840\,
            DOUT => \N__11839\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11841\,
            PADOUT => \N__11840\,
            PADIN => \N__11839\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8618\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11832\,
            DIN => \N__11831\,
            DOUT => \N__11830\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11832\,
            PADOUT => \N__11831\,
            PADIN => \N__11830\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11823\,
            DIN => \N__11822\,
            DOUT => \N__11821\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11823\,
            PADOUT => \N__11822\,
            PADIN => \N__11821\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11814\,
            DIN => \N__11813\,
            DOUT => \N__11812\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11814\,
            PADOUT => \N__11813\,
            PADIN => \N__11812\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11805\,
            DIN => \N__11804\,
            DOUT => \N__11803\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11805\,
            PADOUT => \N__11804\,
            PADIN => \N__11803\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11796\,
            DIN => \N__11795\,
            DOUT => \N__11794\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11796\,
            PADOUT => \N__11795\,
            PADIN => \N__11794\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9481\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11787\,
            DIN => \N__11786\,
            DOUT => \N__11785\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11787\,
            PADOUT => \N__11786\,
            PADIN => \N__11785\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9917\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11778\,
            DIN => \N__11777\,
            DOUT => \N__11776\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11778\,
            PADOUT => \N__11777\,
            PADIN => \N__11776\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8393\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11769\,
            DIN => \N__11768\,
            DOUT => \N__11767\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11769\,
            PADOUT => \N__11768\,
            PADIN => \N__11767\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11243\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2838\ : InMux
    port map (
            O => \N__11750\,
            I => \N__11745\
        );

    \I__2837\ : InMux
    port map (
            O => \N__11749\,
            I => \N__11738\
        );

    \I__2836\ : InMux
    port map (
            O => \N__11748\,
            I => \N__11738\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__11745\,
            I => \N__11735\
        );

    \I__2834\ : InMux
    port map (
            O => \N__11744\,
            I => \N__11732\
        );

    \I__2833\ : CascadeMux
    port map (
            O => \N__11743\,
            I => \N__11728\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__11738\,
            I => \N__11725\
        );

    \I__2831\ : Sp12to4
    port map (
            O => \N__11735\,
            I => \N__11722\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__11732\,
            I => \N__11719\
        );

    \I__2829\ : InMux
    port map (
            O => \N__11731\,
            I => \N__11716\
        );

    \I__2828\ : InMux
    port map (
            O => \N__11728\,
            I => \N__11713\
        );

    \I__2827\ : Span12Mux_h
    port map (
            O => \N__11725\,
            I => \N__11710\
        );

    \I__2826\ : Span12Mux_v
    port map (
            O => \N__11722\,
            I => \N__11707\
        );

    \I__2825\ : Span12Mux_h
    port map (
            O => \N__11719\,
            I => \N__11700\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__11716\,
            I => \N__11700\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__11713\,
            I => \N__11700\
        );

    \I__2822\ : Span12Mux_v
    port map (
            O => \N__11710\,
            I => \N__11697\
        );

    \I__2821\ : Span12Mux_h
    port map (
            O => \N__11707\,
            I => \N__11692\
        );

    \I__2820\ : Span12Mux_v
    port map (
            O => \N__11700\,
            I => \N__11692\
        );

    \I__2819\ : Odrv12
    port map (
            O => \N__11697\,
            I => \CASLn_c\
        );

    \I__2818\ : Odrv12
    port map (
            O => \N__11692\,
            I => \CASLn_c\
        );

    \I__2817\ : InMux
    port map (
            O => \N__11687\,
            I => \N__11684\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__11684\,
            I => \N__11681\
        );

    \I__2815\ : Span4Mux_v
    port map (
            O => \N__11681\,
            I => \N__11678\
        );

    \I__2814\ : Sp12to4
    port map (
            O => \N__11678\,
            I => \N__11674\
        );

    \I__2813\ : InMux
    port map (
            O => \N__11677\,
            I => \N__11671\
        );

    \I__2812\ : Span12Mux_h
    port map (
            O => \N__11674\,
            I => \N__11665\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__11671\,
            I => \N__11665\
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__11670\,
            I => \N__11662\
        );

    \I__2809\ : Span12Mux_s11_v
    port map (
            O => \N__11665\,
            I => \N__11659\
        );

    \I__2808\ : InMux
    port map (
            O => \N__11662\,
            I => \N__11656\
        );

    \I__2807\ : Odrv12
    port map (
            O => \N__11659\,
            I => \DMA_WRITE_CYCLE\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__11656\,
            I => \DMA_WRITE_CYCLE\
        );

    \I__2805\ : IoInMux
    port map (
            O => \N__11651\,
            I => \N__11648\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__11648\,
            I => \N__11645\
        );

    \I__2803\ : IoSpan4Mux
    port map (
            O => \N__11645\,
            I => \N__11642\
        );

    \I__2802\ : Span4Mux_s3_v
    port map (
            O => \N__11642\,
            I => \N__11639\
        );

    \I__2801\ : Span4Mux_v
    port map (
            O => \N__11639\,
            I => \N__11636\
        );

    \I__2800\ : Odrv4
    port map (
            O => \N__11636\,
            I => \N_357\
        );

    \I__2799\ : IoInMux
    port map (
            O => \N__11633\,
            I => \N__11630\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__11630\,
            I => \N__11627\
        );

    \I__2797\ : Span4Mux_s3_v
    port map (
            O => \N__11627\,
            I => \N__11624\
        );

    \I__2796\ : Odrv4
    port map (
            O => \N__11624\,
            I => \N_373_i\
        );

    \I__2795\ : InMux
    port map (
            O => \N__11621\,
            I => \N__11615\
        );

    \I__2794\ : InMux
    port map (
            O => \N__11620\,
            I => \N__11615\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__11615\,
            I => \N__11606\
        );

    \I__2792\ : InMux
    port map (
            O => \N__11614\,
            I => \N__11599\
        );

    \I__2791\ : InMux
    port map (
            O => \N__11613\,
            I => \N__11599\
        );

    \I__2790\ : InMux
    port map (
            O => \N__11612\,
            I => \N__11599\
        );

    \I__2789\ : InMux
    port map (
            O => \N__11611\,
            I => \N__11596\
        );

    \I__2788\ : InMux
    port map (
            O => \N__11610\,
            I => \N__11591\
        );

    \I__2787\ : InMux
    port map (
            O => \N__11609\,
            I => \N__11591\
        );

    \I__2786\ : Span4Mux_v
    port map (
            O => \N__11606\,
            I => \N__11588\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__11599\,
            I => \N__11585\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__11596\,
            I => \N__11582\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__11591\,
            I => \N__11579\
        );

    \I__2782\ : Span4Mux_v
    port map (
            O => \N__11588\,
            I => \N__11574\
        );

    \I__2781\ : Span4Mux_v
    port map (
            O => \N__11585\,
            I => \N__11574\
        );

    \I__2780\ : Span4Mux_v
    port map (
            O => \N__11582\,
            I => \N__11571\
        );

    \I__2779\ : Span12Mux_v
    port map (
            O => \N__11579\,
            I => \N__11568\
        );

    \I__2778\ : Sp12to4
    port map (
            O => \N__11574\,
            I => \N__11563\
        );

    \I__2777\ : Sp12to4
    port map (
            O => \N__11571\,
            I => \N__11563\
        );

    \I__2776\ : Span12Mux_h
    port map (
            O => \N__11568\,
            I => \N__11560\
        );

    \I__2775\ : Span12Mux_h
    port map (
            O => \N__11563\,
            I => \N__11557\
        );

    \I__2774\ : Odrv12
    port map (
            O => \N__11560\,
            I => \A_c_1\
        );

    \I__2773\ : Odrv12
    port map (
            O => \N__11557\,
            I => \A_c_1\
        );

    \I__2772\ : InMux
    port map (
            O => \N__11552\,
            I => \N__11540\
        );

    \I__2771\ : InMux
    port map (
            O => \N__11551\,
            I => \N__11540\
        );

    \I__2770\ : InMux
    port map (
            O => \N__11550\,
            I => \N__11540\
        );

    \I__2769\ : InMux
    port map (
            O => \N__11549\,
            I => \N__11535\
        );

    \I__2768\ : InMux
    port map (
            O => \N__11548\,
            I => \N__11535\
        );

    \I__2767\ : InMux
    port map (
            O => \N__11547\,
            I => \N__11531\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__11540\,
            I => \N__11527\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__11535\,
            I => \N__11524\
        );

    \I__2764\ : InMux
    port map (
            O => \N__11534\,
            I => \N__11521\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__11531\,
            I => \N__11518\
        );

    \I__2762\ : InMux
    port map (
            O => \N__11530\,
            I => \N__11515\
        );

    \I__2761\ : Span4Mux_v
    port map (
            O => \N__11527\,
            I => \N__11510\
        );

    \I__2760\ : Span4Mux_v
    port map (
            O => \N__11524\,
            I => \N__11510\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__11521\,
            I => \N__11507\
        );

    \I__2758\ : Span4Mux_v
    port map (
            O => \N__11518\,
            I => \N__11503\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__11515\,
            I => \N__11500\
        );

    \I__2756\ : Span4Mux_h
    port map (
            O => \N__11510\,
            I => \N__11495\
        );

    \I__2755\ : Span4Mux_v
    port map (
            O => \N__11507\,
            I => \N__11495\
        );

    \I__2754\ : InMux
    port map (
            O => \N__11506\,
            I => \N__11492\
        );

    \I__2753\ : Sp12to4
    port map (
            O => \N__11503\,
            I => \N__11487\
        );

    \I__2752\ : Span12Mux_v
    port map (
            O => \N__11500\,
            I => \N__11487\
        );

    \I__2751\ : Sp12to4
    port map (
            O => \N__11495\,
            I => \N__11482\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__11492\,
            I => \N__11482\
        );

    \I__2749\ : Span12Mux_h
    port map (
            O => \N__11487\,
            I => \N__11479\
        );

    \I__2748\ : Span12Mux_h
    port map (
            O => \N__11482\,
            I => \N__11476\
        );

    \I__2747\ : Odrv12
    port map (
            O => \N__11479\,
            I => \A_c_0\
        );

    \I__2746\ : Odrv12
    port map (
            O => \N__11476\,
            I => \A_c_0\
        );

    \I__2745\ : InMux
    port map (
            O => \N__11471\,
            I => \N__11467\
        );

    \I__2744\ : InMux
    port map (
            O => \N__11470\,
            I => \N__11459\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__11467\,
            I => \N__11456\
        );

    \I__2742\ : InMux
    port map (
            O => \N__11466\,
            I => \N__11453\
        );

    \I__2741\ : InMux
    port map (
            O => \N__11465\,
            I => \N__11450\
        );

    \I__2740\ : CascadeMux
    port map (
            O => \N__11464\,
            I => \N__11447\
        );

    \I__2739\ : CascadeMux
    port map (
            O => \N__11463\,
            I => \N__11444\
        );

    \I__2738\ : CascadeMux
    port map (
            O => \N__11462\,
            I => \N__11441\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__11459\,
            I => \N__11437\
        );

    \I__2736\ : Span4Mux_v
    port map (
            O => \N__11456\,
            I => \N__11432\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__11453\,
            I => \N__11432\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__11450\,
            I => \N__11429\
        );

    \I__2733\ : InMux
    port map (
            O => \N__11447\,
            I => \N__11422\
        );

    \I__2732\ : InMux
    port map (
            O => \N__11444\,
            I => \N__11422\
        );

    \I__2731\ : InMux
    port map (
            O => \N__11441\,
            I => \N__11422\
        );

    \I__2730\ : InMux
    port map (
            O => \N__11440\,
            I => \N__11419\
        );

    \I__2729\ : Span4Mux_v
    port map (
            O => \N__11437\,
            I => \N__11416\
        );

    \I__2728\ : Span4Mux_h
    port map (
            O => \N__11432\,
            I => \N__11411\
        );

    \I__2727\ : Span4Mux_v
    port map (
            O => \N__11429\,
            I => \N__11411\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__11422\,
            I => \N__11406\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__11419\,
            I => \N__11406\
        );

    \I__2724\ : Span4Mux_v
    port map (
            O => \N__11416\,
            I => \N__11403\
        );

    \I__2723\ : Span4Mux_v
    port map (
            O => \N__11411\,
            I => \N__11398\
        );

    \I__2722\ : Span4Mux_h
    port map (
            O => \N__11406\,
            I => \N__11398\
        );

    \I__2721\ : Span4Mux_v
    port map (
            O => \N__11403\,
            I => \N__11395\
        );

    \I__2720\ : Span4Mux_v
    port map (
            O => \N__11398\,
            I => \N__11392\
        );

    \I__2719\ : Sp12to4
    port map (
            O => \N__11395\,
            I => \N__11387\
        );

    \I__2718\ : Sp12to4
    port map (
            O => \N__11392\,
            I => \N__11387\
        );

    \I__2717\ : Span12Mux_h
    port map (
            O => \N__11387\,
            I => \N__11384\
        );

    \I__2716\ : Odrv12
    port map (
            O => \N__11384\,
            I => \SIZ_c_0\
        );

    \I__2715\ : CascadeMux
    port map (
            O => \N__11381\,
            I => \N__11376\
        );

    \I__2714\ : InMux
    port map (
            O => \N__11380\,
            I => \N__11372\
        );

    \I__2713\ : InMux
    port map (
            O => \N__11379\,
            I => \N__11369\
        );

    \I__2712\ : InMux
    port map (
            O => \N__11376\,
            I => \N__11366\
        );

    \I__2711\ : InMux
    port map (
            O => \N__11375\,
            I => \N__11363\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__11372\,
            I => \N__11357\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__11369\,
            I => \N__11357\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__11366\,
            I => \N__11354\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__11363\,
            I => \N__11351\
        );

    \I__2706\ : CascadeMux
    port map (
            O => \N__11362\,
            I => \N__11345\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__11357\,
            I => \N__11342\
        );

    \I__2704\ : Span4Mux_h
    port map (
            O => \N__11354\,
            I => \N__11337\
        );

    \I__2703\ : Span4Mux_v
    port map (
            O => \N__11351\,
            I => \N__11337\
        );

    \I__2702\ : InMux
    port map (
            O => \N__11350\,
            I => \N__11329\
        );

    \I__2701\ : InMux
    port map (
            O => \N__11349\,
            I => \N__11329\
        );

    \I__2700\ : InMux
    port map (
            O => \N__11348\,
            I => \N__11329\
        );

    \I__2699\ : InMux
    port map (
            O => \N__11345\,
            I => \N__11326\
        );

    \I__2698\ : Span4Mux_v
    port map (
            O => \N__11342\,
            I => \N__11323\
        );

    \I__2697\ : Span4Mux_v
    port map (
            O => \N__11337\,
            I => \N__11320\
        );

    \I__2696\ : InMux
    port map (
            O => \N__11336\,
            I => \N__11317\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__11329\,
            I => \N__11312\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__11326\,
            I => \N__11312\
        );

    \I__2693\ : Span4Mux_v
    port map (
            O => \N__11323\,
            I => \N__11309\
        );

    \I__2692\ : Span4Mux_v
    port map (
            O => \N__11320\,
            I => \N__11306\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__11317\,
            I => \N__11301\
        );

    \I__2690\ : Sp12to4
    port map (
            O => \N__11312\,
            I => \N__11301\
        );

    \I__2689\ : Sp12to4
    port map (
            O => \N__11309\,
            I => \N__11294\
        );

    \I__2688\ : Sp12to4
    port map (
            O => \N__11306\,
            I => \N__11294\
        );

    \I__2687\ : Span12Mux_v
    port map (
            O => \N__11301\,
            I => \N__11294\
        );

    \I__2686\ : Span12Mux_h
    port map (
            O => \N__11294\,
            I => \N__11291\
        );

    \I__2685\ : Odrv12
    port map (
            O => \N__11291\,
            I => \SIZ_c_1\
        );

    \I__2684\ : IoInMux
    port map (
            O => \N__11288\,
            I => \N__11285\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__11285\,
            I => \N__11282\
        );

    \I__2682\ : Span4Mux_s2_v
    port map (
            O => \N__11282\,
            I => \N__11279\
        );

    \I__2681\ : Span4Mux_h
    port map (
            O => \N__11279\,
            I => \N__11276\
        );

    \I__2680\ : Span4Mux_v
    port map (
            O => \N__11276\,
            I => \N__11273\
        );

    \I__2679\ : Odrv4
    port map (
            O => \N__11273\,
            I => \UMBEn_c\
        );

    \I__2678\ : InMux
    port map (
            O => \N__11270\,
            I => \N__11267\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__11267\,
            I => \N__11264\
        );

    \I__2676\ : Odrv12
    port map (
            O => \N__11264\,
            I => \U712_CHIP_RAM.CMA_5_i_0_9\
        );

    \I__2675\ : InMux
    port map (
            O => \N__11261\,
            I => \N__11258\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__11258\,
            I => \N__11255\
        );

    \I__2673\ : Sp12to4
    port map (
            O => \N__11255\,
            I => \N__11252\
        );

    \I__2672\ : Span12Mux_v
    port map (
            O => \N__11252\,
            I => \N__11249\
        );

    \I__2671\ : Span12Mux_h
    port map (
            O => \N__11249\,
            I => \N__11246\
        );

    \I__2670\ : Odrv12
    port map (
            O => \N__11246\,
            I => \A_c_19\
        );

    \I__2669\ : IoInMux
    port map (
            O => \N__11243\,
            I => \N__11240\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__11240\,
            I => \N__11237\
        );

    \I__2667\ : IoSpan4Mux
    port map (
            O => \N__11237\,
            I => \N__11234\
        );

    \I__2666\ : IoSpan4Mux
    port map (
            O => \N__11234\,
            I => \N__11231\
        );

    \I__2665\ : Span4Mux_s2_h
    port map (
            O => \N__11231\,
            I => \N__11228\
        );

    \I__2664\ : Sp12to4
    port map (
            O => \N__11228\,
            I => \N__11225\
        );

    \I__2663\ : Odrv12
    port map (
            O => \N__11225\,
            I => \CMA_c_9\
        );

    \I__2662\ : CEMux
    port map (
            O => \N__11222\,
            I => \N__11219\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__11219\,
            I => \N__11214\
        );

    \I__2660\ : CEMux
    port map (
            O => \N__11218\,
            I => \N__11211\
        );

    \I__2659\ : CEMux
    port map (
            O => \N__11217\,
            I => \N__11208\
        );

    \I__2658\ : Span4Mux_v
    port map (
            O => \N__11214\,
            I => \N__11202\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__11211\,
            I => \N__11202\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__11208\,
            I => \N__11199\
        );

    \I__2655\ : CEMux
    port map (
            O => \N__11207\,
            I => \N__11196\
        );

    \I__2654\ : Sp12to4
    port map (
            O => \N__11202\,
            I => \N__11192\
        );

    \I__2653\ : Span4Mux_h
    port map (
            O => \N__11199\,
            I => \N__11187\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__11196\,
            I => \N__11187\
        );

    \I__2651\ : CEMux
    port map (
            O => \N__11195\,
            I => \N__11184\
        );

    \I__2650\ : Span12Mux_h
    port map (
            O => \N__11192\,
            I => \N__11179\
        );

    \I__2649\ : Sp12to4
    port map (
            O => \N__11187\,
            I => \N__11179\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__11184\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__2647\ : Odrv12
    port map (
            O => \N__11179\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__2646\ : CascadeMux
    port map (
            O => \N__11174\,
            I => \N__11169\
        );

    \I__2645\ : InMux
    port map (
            O => \N__11173\,
            I => \N__11165\
        );

    \I__2644\ : InMux
    port map (
            O => \N__11172\,
            I => \N__11160\
        );

    \I__2643\ : InMux
    port map (
            O => \N__11169\,
            I => \N__11157\
        );

    \I__2642\ : InMux
    port map (
            O => \N__11168\,
            I => \N__11154\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__11165\,
            I => \N__11150\
        );

    \I__2640\ : InMux
    port map (
            O => \N__11164\,
            I => \N__11147\
        );

    \I__2639\ : InMux
    port map (
            O => \N__11163\,
            I => \N__11144\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__11160\,
            I => \N__11141\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__11157\,
            I => \N__11138\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__11154\,
            I => \N__11135\
        );

    \I__2635\ : InMux
    port map (
            O => \N__11153\,
            I => \N__11132\
        );

    \I__2634\ : Span4Mux_h
    port map (
            O => \N__11150\,
            I => \N__11126\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__11147\,
            I => \N__11126\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__11144\,
            I => \N__11123\
        );

    \I__2631\ : Span4Mux_v
    port map (
            O => \N__11141\,
            I => \N__11118\
        );

    \I__2630\ : Span4Mux_v
    port map (
            O => \N__11138\,
            I => \N__11118\
        );

    \I__2629\ : Span4Mux_h
    port map (
            O => \N__11135\,
            I => \N__11113\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__11132\,
            I => \N__11113\
        );

    \I__2627\ : InMux
    port map (
            O => \N__11131\,
            I => \N__11110\
        );

    \I__2626\ : Odrv4
    port map (
            O => \N__11126\,
            I => \DMA_CYCLEm\
        );

    \I__2625\ : Odrv4
    port map (
            O => \N__11123\,
            I => \DMA_CYCLEm\
        );

    \I__2624\ : Odrv4
    port map (
            O => \N__11118\,
            I => \DMA_CYCLEm\
        );

    \I__2623\ : Odrv4
    port map (
            O => \N__11113\,
            I => \DMA_CYCLEm\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__11110\,
            I => \DMA_CYCLEm\
        );

    \I__2621\ : InMux
    port map (
            O => \N__11099\,
            I => \N__11096\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__11096\,
            I => \U712_BYTE_ENABLE.N_411\
        );

    \I__2619\ : IoInMux
    port map (
            O => \N__11093\,
            I => \N__11090\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__11090\,
            I => \N__11085\
        );

    \I__2617\ : InMux
    port map (
            O => \N__11089\,
            I => \N__11082\
        );

    \I__2616\ : InMux
    port map (
            O => \N__11088\,
            I => \N__11079\
        );

    \I__2615\ : Span4Mux_s2_v
    port map (
            O => \N__11085\,
            I => \N__11075\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__11082\,
            I => \N__11072\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__11079\,
            I => \N__11069\
        );

    \I__2612\ : InMux
    port map (
            O => \N__11078\,
            I => \N__11066\
        );

    \I__2611\ : Span4Mux_v
    port map (
            O => \N__11075\,
            I => \N__11063\
        );

    \I__2610\ : Span4Mux_v
    port map (
            O => \N__11072\,
            I => \N__11059\
        );

    \I__2609\ : Span4Mux_v
    port map (
            O => \N__11069\,
            I => \N__11056\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__11066\,
            I => \N__11053\
        );

    \I__2607\ : Sp12to4
    port map (
            O => \N__11063\,
            I => \N__11050\
        );

    \I__2606\ : InMux
    port map (
            O => \N__11062\,
            I => \N__11047\
        );

    \I__2605\ : Span4Mux_v
    port map (
            O => \N__11059\,
            I => \N__11043\
        );

    \I__2604\ : Span4Mux_h
    port map (
            O => \N__11056\,
            I => \N__11038\
        );

    \I__2603\ : Span4Mux_v
    port map (
            O => \N__11053\,
            I => \N__11038\
        );

    \I__2602\ : Span12Mux_h
    port map (
            O => \N__11050\,
            I => \N__11033\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__11047\,
            I => \N__11033\
        );

    \I__2600\ : InMux
    port map (
            O => \N__11046\,
            I => \N__11030\
        );

    \I__2599\ : Odrv4
    port map (
            O => \N__11043\,
            I => \DBENn_c\
        );

    \I__2598\ : Odrv4
    port map (
            O => \N__11038\,
            I => \DBENn_c\
        );

    \I__2597\ : Odrv12
    port map (
            O => \N__11033\,
            I => \DBENn_c\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__11030\,
            I => \DBENn_c\
        );

    \I__2595\ : IoInMux
    port map (
            O => \N__11021\,
            I => \N__11018\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__11018\,
            I => \N__11015\
        );

    \I__2593\ : Span4Mux_s1_h
    port map (
            O => \N__11015\,
            I => \N__11012\
        );

    \I__2592\ : Sp12to4
    port map (
            O => \N__11012\,
            I => \N__11009\
        );

    \I__2591\ : Span12Mux_v
    port map (
            O => \N__11009\,
            I => \N__11006\
        );

    \I__2590\ : Span12Mux_h
    port map (
            O => \N__11006\,
            I => \N__11003\
        );

    \I__2589\ : Odrv12
    port map (
            O => \N__11003\,
            I => \N_150_i\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__11000\,
            I => \N__10991\
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__10999\,
            I => \N__10987\
        );

    \I__2586\ : CascadeMux
    port map (
            O => \N__10998\,
            I => \N__10984\
        );

    \I__2585\ : CascadeMux
    port map (
            O => \N__10997\,
            I => \N__10975\
        );

    \I__2584\ : InMux
    port map (
            O => \N__10996\,
            I => \N__10972\
        );

    \I__2583\ : InMux
    port map (
            O => \N__10995\,
            I => \N__10969\
        );

    \I__2582\ : InMux
    port map (
            O => \N__10994\,
            I => \N__10954\
        );

    \I__2581\ : InMux
    port map (
            O => \N__10991\,
            I => \N__10954\
        );

    \I__2580\ : InMux
    port map (
            O => \N__10990\,
            I => \N__10954\
        );

    \I__2579\ : InMux
    port map (
            O => \N__10987\,
            I => \N__10954\
        );

    \I__2578\ : InMux
    port map (
            O => \N__10984\,
            I => \N__10954\
        );

    \I__2577\ : InMux
    port map (
            O => \N__10983\,
            I => \N__10954\
        );

    \I__2576\ : InMux
    port map (
            O => \N__10982\,
            I => \N__10954\
        );

    \I__2575\ : InMux
    port map (
            O => \N__10981\,
            I => \N__10949\
        );

    \I__2574\ : InMux
    port map (
            O => \N__10980\,
            I => \N__10949\
        );

    \I__2573\ : InMux
    port map (
            O => \N__10979\,
            I => \N__10946\
        );

    \I__2572\ : InMux
    port map (
            O => \N__10978\,
            I => \N__10942\
        );

    \I__2571\ : InMux
    port map (
            O => \N__10975\,
            I => \N__10939\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__10972\,
            I => \N__10924\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__10969\,
            I => \N__10924\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__10954\,
            I => \N__10924\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__10949\,
            I => \N__10924\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__10946\,
            I => \N__10921\
        );

    \I__2565\ : InMux
    port map (
            O => \N__10945\,
            I => \N__10918\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__10942\,
            I => \N__10915\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__10939\,
            I => \N__10912\
        );

    \I__2562\ : InMux
    port map (
            O => \N__10938\,
            I => \N__10905\
        );

    \I__2561\ : InMux
    port map (
            O => \N__10937\,
            I => \N__10905\
        );

    \I__2560\ : InMux
    port map (
            O => \N__10936\,
            I => \N__10905\
        );

    \I__2559\ : InMux
    port map (
            O => \N__10935\,
            I => \N__10902\
        );

    \I__2558\ : InMux
    port map (
            O => \N__10934\,
            I => \N__10899\
        );

    \I__2557\ : InMux
    port map (
            O => \N__10933\,
            I => \N__10896\
        );

    \I__2556\ : Span4Mux_v
    port map (
            O => \N__10924\,
            I => \N__10889\
        );

    \I__2555\ : Span4Mux_h
    port map (
            O => \N__10921\,
            I => \N__10889\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__10918\,
            I => \N__10889\
        );

    \I__2553\ : Span4Mux_v
    port map (
            O => \N__10915\,
            I => \N__10886\
        );

    \I__2552\ : Span12Mux_h
    port map (
            O => \N__10912\,
            I => \N__10879\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__10905\,
            I => \N__10879\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__10902\,
            I => \N__10879\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__10899\,
            I => \N__10872\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__10896\,
            I => \N__10872\
        );

    \I__2547\ : Sp12to4
    port map (
            O => \N__10889\,
            I => \N__10872\
        );

    \I__2546\ : Sp12to4
    port map (
            O => \N__10886\,
            I => \N__10869\
        );

    \I__2545\ : Span12Mux_h
    port map (
            O => \N__10879\,
            I => \N__10866\
        );

    \I__2544\ : Span12Mux_v
    port map (
            O => \N__10872\,
            I => \N__10863\
        );

    \I__2543\ : Span12Mux_h
    port map (
            O => \N__10869\,
            I => \N__10860\
        );

    \I__2542\ : Span12Mux_v
    port map (
            O => \N__10866\,
            I => \N__10855\
        );

    \I__2541\ : Span12Mux_h
    port map (
            O => \N__10863\,
            I => \N__10855\
        );

    \I__2540\ : Span12Mux_v
    port map (
            O => \N__10860\,
            I => \N__10852\
        );

    \I__2539\ : Odrv12
    port map (
            O => \N__10855\,
            I => \AGNUS_REV_c\
        );

    \I__2538\ : Odrv12
    port map (
            O => \N__10852\,
            I => \AGNUS_REV_c\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__10847\,
            I => \N__10842\
        );

    \I__2536\ : InMux
    port map (
            O => \N__10846\,
            I => \N__10839\
        );

    \I__2535\ : InMux
    port map (
            O => \N__10845\,
            I => \N__10836\
        );

    \I__2534\ : InMux
    port map (
            O => \N__10842\,
            I => \N__10833\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__10839\,
            I => \N__10829\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__10836\,
            I => \N__10824\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__10833\,
            I => \N__10824\
        );

    \I__2530\ : InMux
    port map (
            O => \N__10832\,
            I => \N__10821\
        );

    \I__2529\ : Span4Mux_h
    port map (
            O => \N__10829\,
            I => \N__10814\
        );

    \I__2528\ : Span4Mux_v
    port map (
            O => \N__10824\,
            I => \N__10814\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__10821\,
            I => \N__10814\
        );

    \I__2526\ : Span4Mux_h
    port map (
            O => \N__10814\,
            I => \N__10811\
        );

    \I__2525\ : Span4Mux_v
    port map (
            O => \N__10811\,
            I => \N__10808\
        );

    \I__2524\ : Sp12to4
    port map (
            O => \N__10808\,
            I => \N__10805\
        );

    \I__2523\ : Span12Mux_v
    port map (
            O => \N__10805\,
            I => \N__10802\
        );

    \I__2522\ : Odrv12
    port map (
            O => \N__10802\,
            I => \DRA_c_9\
        );

    \I__2521\ : InMux
    port map (
            O => \N__10799\,
            I => \N__10796\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__10796\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2519\ : ClkMux
    port map (
            O => \N__10793\,
            I => \N__10775\
        );

    \I__2518\ : ClkMux
    port map (
            O => \N__10792\,
            I => \N__10775\
        );

    \I__2517\ : ClkMux
    port map (
            O => \N__10791\,
            I => \N__10775\
        );

    \I__2516\ : ClkMux
    port map (
            O => \N__10790\,
            I => \N__10775\
        );

    \I__2515\ : ClkMux
    port map (
            O => \N__10789\,
            I => \N__10775\
        );

    \I__2514\ : ClkMux
    port map (
            O => \N__10788\,
            I => \N__10775\
        );

    \I__2513\ : GlobalMux
    port map (
            O => \N__10775\,
            I => \N__10772\
        );

    \I__2512\ : gio2CtrlBuf
    port map (
            O => \N__10772\,
            I => \C3_c_g\
        );

    \I__2511\ : CEMux
    port map (
            O => \N__10769\,
            I => \N__10742\
        );

    \I__2510\ : CEMux
    port map (
            O => \N__10768\,
            I => \N__10742\
        );

    \I__2509\ : CEMux
    port map (
            O => \N__10767\,
            I => \N__10742\
        );

    \I__2508\ : CEMux
    port map (
            O => \N__10766\,
            I => \N__10742\
        );

    \I__2507\ : CEMux
    port map (
            O => \N__10765\,
            I => \N__10742\
        );

    \I__2506\ : CEMux
    port map (
            O => \N__10764\,
            I => \N__10742\
        );

    \I__2505\ : CEMux
    port map (
            O => \N__10763\,
            I => \N__10742\
        );

    \I__2504\ : CEMux
    port map (
            O => \N__10762\,
            I => \N__10742\
        );

    \I__2503\ : CEMux
    port map (
            O => \N__10761\,
            I => \N__10742\
        );

    \I__2502\ : GlobalMux
    port map (
            O => \N__10742\,
            I => \N__10739\
        );

    \I__2501\ : gio2CtrlBuf
    port map (
            O => \N__10739\,
            I => \DBRn_c_i_0_g\
        );

    \I__2500\ : InMux
    port map (
            O => \N__10736\,
            I => \N__10726\
        );

    \I__2499\ : InMux
    port map (
            O => \N__10735\,
            I => \N__10719\
        );

    \I__2498\ : InMux
    port map (
            O => \N__10734\,
            I => \N__10719\
        );

    \I__2497\ : InMux
    port map (
            O => \N__10733\,
            I => \N__10719\
        );

    \I__2496\ : InMux
    port map (
            O => \N__10732\,
            I => \N__10716\
        );

    \I__2495\ : InMux
    port map (
            O => \N__10731\,
            I => \N__10711\
        );

    \I__2494\ : InMux
    port map (
            O => \N__10730\,
            I => \N__10711\
        );

    \I__2493\ : InMux
    port map (
            O => \N__10729\,
            I => \N__10708\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__10726\,
            I => \N__10704\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__10719\,
            I => \N__10691\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__10716\,
            I => \N__10683\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__10711\,
            I => \N__10676\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__10708\,
            I => \N__10658\
        );

    \I__2487\ : SRMux
    port map (
            O => \N__10707\,
            I => \N__10574\
        );

    \I__2486\ : Glb2LocalMux
    port map (
            O => \N__10704\,
            I => \N__10574\
        );

    \I__2485\ : SRMux
    port map (
            O => \N__10703\,
            I => \N__10574\
        );

    \I__2484\ : SRMux
    port map (
            O => \N__10702\,
            I => \N__10574\
        );

    \I__2483\ : SRMux
    port map (
            O => \N__10701\,
            I => \N__10574\
        );

    \I__2482\ : SRMux
    port map (
            O => \N__10700\,
            I => \N__10574\
        );

    \I__2481\ : SRMux
    port map (
            O => \N__10699\,
            I => \N__10574\
        );

    \I__2480\ : SRMux
    port map (
            O => \N__10698\,
            I => \N__10574\
        );

    \I__2479\ : SRMux
    port map (
            O => \N__10697\,
            I => \N__10574\
        );

    \I__2478\ : SRMux
    port map (
            O => \N__10696\,
            I => \N__10574\
        );

    \I__2477\ : SRMux
    port map (
            O => \N__10695\,
            I => \N__10574\
        );

    \I__2476\ : SRMux
    port map (
            O => \N__10694\,
            I => \N__10574\
        );

    \I__2475\ : Glb2LocalMux
    port map (
            O => \N__10691\,
            I => \N__10574\
        );

    \I__2474\ : SRMux
    port map (
            O => \N__10690\,
            I => \N__10574\
        );

    \I__2473\ : SRMux
    port map (
            O => \N__10689\,
            I => \N__10574\
        );

    \I__2472\ : SRMux
    port map (
            O => \N__10688\,
            I => \N__10574\
        );

    \I__2471\ : SRMux
    port map (
            O => \N__10687\,
            I => \N__10574\
        );

    \I__2470\ : SRMux
    port map (
            O => \N__10686\,
            I => \N__10574\
        );

    \I__2469\ : Glb2LocalMux
    port map (
            O => \N__10683\,
            I => \N__10574\
        );

    \I__2468\ : SRMux
    port map (
            O => \N__10682\,
            I => \N__10574\
        );

    \I__2467\ : SRMux
    port map (
            O => \N__10681\,
            I => \N__10574\
        );

    \I__2466\ : SRMux
    port map (
            O => \N__10680\,
            I => \N__10574\
        );

    \I__2465\ : SRMux
    port map (
            O => \N__10679\,
            I => \N__10574\
        );

    \I__2464\ : Glb2LocalMux
    port map (
            O => \N__10676\,
            I => \N__10574\
        );

    \I__2463\ : SRMux
    port map (
            O => \N__10675\,
            I => \N__10574\
        );

    \I__2462\ : SRMux
    port map (
            O => \N__10674\,
            I => \N__10574\
        );

    \I__2461\ : SRMux
    port map (
            O => \N__10673\,
            I => \N__10574\
        );

    \I__2460\ : SRMux
    port map (
            O => \N__10672\,
            I => \N__10574\
        );

    \I__2459\ : SRMux
    port map (
            O => \N__10671\,
            I => \N__10574\
        );

    \I__2458\ : SRMux
    port map (
            O => \N__10670\,
            I => \N__10574\
        );

    \I__2457\ : SRMux
    port map (
            O => \N__10669\,
            I => \N__10574\
        );

    \I__2456\ : SRMux
    port map (
            O => \N__10668\,
            I => \N__10574\
        );

    \I__2455\ : SRMux
    port map (
            O => \N__10667\,
            I => \N__10574\
        );

    \I__2454\ : SRMux
    port map (
            O => \N__10666\,
            I => \N__10574\
        );

    \I__2453\ : SRMux
    port map (
            O => \N__10665\,
            I => \N__10574\
        );

    \I__2452\ : SRMux
    port map (
            O => \N__10664\,
            I => \N__10574\
        );

    \I__2451\ : SRMux
    port map (
            O => \N__10663\,
            I => \N__10574\
        );

    \I__2450\ : SRMux
    port map (
            O => \N__10662\,
            I => \N__10574\
        );

    \I__2449\ : SRMux
    port map (
            O => \N__10661\,
            I => \N__10574\
        );

    \I__2448\ : Glb2LocalMux
    port map (
            O => \N__10658\,
            I => \N__10574\
        );

    \I__2447\ : SRMux
    port map (
            O => \N__10657\,
            I => \N__10574\
        );

    \I__2446\ : GlobalMux
    port map (
            O => \N__10574\,
            I => \N__10571\
        );

    \I__2445\ : gio2CtrlBuf
    port map (
            O => \N__10571\,
            I => \RESETn_c_i_g\
        );

    \I__2444\ : CascadeMux
    port map (
            O => \N__10568\,
            I => \N__10564\
        );

    \I__2443\ : InMux
    port map (
            O => \N__10567\,
            I => \N__10555\
        );

    \I__2442\ : InMux
    port map (
            O => \N__10564\,
            I => \N__10542\
        );

    \I__2441\ : InMux
    port map (
            O => \N__10563\,
            I => \N__10535\
        );

    \I__2440\ : InMux
    port map (
            O => \N__10562\,
            I => \N__10535\
        );

    \I__2439\ : InMux
    port map (
            O => \N__10561\,
            I => \N__10535\
        );

    \I__2438\ : InMux
    port map (
            O => \N__10560\,
            I => \N__10528\
        );

    \I__2437\ : InMux
    port map (
            O => \N__10559\,
            I => \N__10528\
        );

    \I__2436\ : InMux
    port map (
            O => \N__10558\,
            I => \N__10528\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__10555\,
            I => \N__10525\
        );

    \I__2434\ : InMux
    port map (
            O => \N__10554\,
            I => \N__10516\
        );

    \I__2433\ : InMux
    port map (
            O => \N__10553\,
            I => \N__10516\
        );

    \I__2432\ : InMux
    port map (
            O => \N__10552\,
            I => \N__10516\
        );

    \I__2431\ : InMux
    port map (
            O => \N__10551\,
            I => \N__10516\
        );

    \I__2430\ : InMux
    port map (
            O => \N__10550\,
            I => \N__10511\
        );

    \I__2429\ : InMux
    port map (
            O => \N__10549\,
            I => \N__10511\
        );

    \I__2428\ : InMux
    port map (
            O => \N__10548\,
            I => \N__10501\
        );

    \I__2427\ : InMux
    port map (
            O => \N__10547\,
            I => \N__10496\
        );

    \I__2426\ : InMux
    port map (
            O => \N__10546\,
            I => \N__10496\
        );

    \I__2425\ : InMux
    port map (
            O => \N__10545\,
            I => \N__10493\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__10542\,
            I => \N__10481\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__10535\,
            I => \N__10481\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__10528\,
            I => \N__10478\
        );

    \I__2421\ : Span4Mux_v
    port map (
            O => \N__10525\,
            I => \N__10471\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__10516\,
            I => \N__10471\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__10511\,
            I => \N__10471\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10510\,
            I => \N__10464\
        );

    \I__2417\ : InMux
    port map (
            O => \N__10509\,
            I => \N__10464\
        );

    \I__2416\ : InMux
    port map (
            O => \N__10508\,
            I => \N__10453\
        );

    \I__2415\ : InMux
    port map (
            O => \N__10507\,
            I => \N__10453\
        );

    \I__2414\ : InMux
    port map (
            O => \N__10506\,
            I => \N__10453\
        );

    \I__2413\ : InMux
    port map (
            O => \N__10505\,
            I => \N__10453\
        );

    \I__2412\ : InMux
    port map (
            O => \N__10504\,
            I => \N__10453\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__10501\,
            I => \N__10446\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__10496\,
            I => \N__10446\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__10493\,
            I => \N__10446\
        );

    \I__2408\ : InMux
    port map (
            O => \N__10492\,
            I => \N__10439\
        );

    \I__2407\ : InMux
    port map (
            O => \N__10491\,
            I => \N__10439\
        );

    \I__2406\ : InMux
    port map (
            O => \N__10490\,
            I => \N__10439\
        );

    \I__2405\ : InMux
    port map (
            O => \N__10489\,
            I => \N__10432\
        );

    \I__2404\ : InMux
    port map (
            O => \N__10488\,
            I => \N__10432\
        );

    \I__2403\ : InMux
    port map (
            O => \N__10487\,
            I => \N__10432\
        );

    \I__2402\ : InMux
    port map (
            O => \N__10486\,
            I => \N__10429\
        );

    \I__2401\ : Span4Mux_v
    port map (
            O => \N__10481\,
            I => \N__10417\
        );

    \I__2400\ : Span4Mux_v
    port map (
            O => \N__10478\,
            I => \N__10417\
        );

    \I__2399\ : Span4Mux_v
    port map (
            O => \N__10471\,
            I => \N__10417\
        );

    \I__2398\ : InMux
    port map (
            O => \N__10470\,
            I => \N__10414\
        );

    \I__2397\ : InMux
    port map (
            O => \N__10469\,
            I => \N__10409\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__10464\,
            I => \N__10406\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__10453\,
            I => \N__10395\
        );

    \I__2394\ : Span4Mux_v
    port map (
            O => \N__10446\,
            I => \N__10395\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__10439\,
            I => \N__10395\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__10432\,
            I => \N__10395\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__10429\,
            I => \N__10395\
        );

    \I__2390\ : InMux
    port map (
            O => \N__10428\,
            I => \N__10390\
        );

    \I__2389\ : InMux
    port map (
            O => \N__10427\,
            I => \N__10390\
        );

    \I__2388\ : InMux
    port map (
            O => \N__10426\,
            I => \N__10383\
        );

    \I__2387\ : InMux
    port map (
            O => \N__10425\,
            I => \N__10383\
        );

    \I__2386\ : InMux
    port map (
            O => \N__10424\,
            I => \N__10383\
        );

    \I__2385\ : Span4Mux_h
    port map (
            O => \N__10417\,
            I => \N__10380\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__10414\,
            I => \N__10377\
        );

    \I__2383\ : InMux
    port map (
            O => \N__10413\,
            I => \N__10372\
        );

    \I__2382\ : InMux
    port map (
            O => \N__10412\,
            I => \N__10372\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__10409\,
            I => \N__10369\
        );

    \I__2380\ : Span4Mux_v
    port map (
            O => \N__10406\,
            I => \N__10364\
        );

    \I__2379\ : Span4Mux_v
    port map (
            O => \N__10395\,
            I => \N__10364\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__10390\,
            I => \N__10359\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__10383\,
            I => \N__10359\
        );

    \I__2376\ : Span4Mux_h
    port map (
            O => \N__10380\,
            I => \N__10354\
        );

    \I__2375\ : Span4Mux_v
    port map (
            O => \N__10377\,
            I => \N__10354\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__10372\,
            I => \N__10351\
        );

    \I__2373\ : Span12Mux_v
    port map (
            O => \N__10369\,
            I => \N__10344\
        );

    \I__2372\ : Sp12to4
    port map (
            O => \N__10364\,
            I => \N__10344\
        );

    \I__2371\ : Span12Mux_v
    port map (
            O => \N__10359\,
            I => \N__10344\
        );

    \I__2370\ : Span4Mux_h
    port map (
            O => \N__10354\,
            I => \N__10341\
        );

    \I__2369\ : Span12Mux_h
    port map (
            O => \N__10351\,
            I => \N__10338\
        );

    \I__2368\ : Span12Mux_h
    port map (
            O => \N__10344\,
            I => \N__10335\
        );

    \I__2367\ : Span4Mux_h
    port map (
            O => \N__10341\,
            I => \N__10332\
        );

    \I__2366\ : Odrv12
    port map (
            O => \N__10338\,
            I => \RESETn_c\
        );

    \I__2365\ : Odrv12
    port map (
            O => \N__10335\,
            I => \RESETn_c\
        );

    \I__2364\ : Odrv4
    port map (
            O => \N__10332\,
            I => \RESETn_c\
        );

    \I__2363\ : InMux
    port map (
            O => \N__10325\,
            I => \N__10322\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__10322\,
            I => \N__10319\
        );

    \I__2361\ : Span12Mux_h
    port map (
            O => \N__10319\,
            I => \N__10316\
        );

    \I__2360\ : Odrv12
    port map (
            O => \N__10316\,
            I => \RAS1n_c\
        );

    \I__2359\ : InMux
    port map (
            O => \N__10313\,
            I => \N__10310\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__10310\,
            I => \N__10306\
        );

    \I__2357\ : InMux
    port map (
            O => \N__10309\,
            I => \N__10303\
        );

    \I__2356\ : Sp12to4
    port map (
            O => \N__10306\,
            I => \N__10300\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__10303\,
            I => \N__10297\
        );

    \I__2354\ : Span12Mux_v
    port map (
            O => \N__10300\,
            I => \N__10294\
        );

    \I__2353\ : Span12Mux_h
    port map (
            O => \N__10297\,
            I => \N__10291\
        );

    \I__2352\ : Odrv12
    port map (
            O => \N__10294\,
            I => \RAS0n_c\
        );

    \I__2351\ : Odrv12
    port map (
            O => \N__10291\,
            I => \RAS0n_c\
        );

    \I__2350\ : InMux
    port map (
            O => \N__10286\,
            I => \N__10283\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__10283\,
            I => \N__10280\
        );

    \I__2348\ : Span12Mux_v
    port map (
            O => \N__10280\,
            I => \N__10277\
        );

    \I__2347\ : Odrv12
    port map (
            O => \N__10277\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2346\ : InMux
    port map (
            O => \N__10274\,
            I => \N__10271\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__10271\,
            I => \N__10243\
        );

    \I__2344\ : ClkMux
    port map (
            O => \N__10270\,
            I => \N__10136\
        );

    \I__2343\ : ClkMux
    port map (
            O => \N__10269\,
            I => \N__10136\
        );

    \I__2342\ : ClkMux
    port map (
            O => \N__10268\,
            I => \N__10136\
        );

    \I__2341\ : ClkMux
    port map (
            O => \N__10267\,
            I => \N__10136\
        );

    \I__2340\ : ClkMux
    port map (
            O => \N__10266\,
            I => \N__10136\
        );

    \I__2339\ : ClkMux
    port map (
            O => \N__10265\,
            I => \N__10136\
        );

    \I__2338\ : ClkMux
    port map (
            O => \N__10264\,
            I => \N__10136\
        );

    \I__2337\ : ClkMux
    port map (
            O => \N__10263\,
            I => \N__10136\
        );

    \I__2336\ : ClkMux
    port map (
            O => \N__10262\,
            I => \N__10136\
        );

    \I__2335\ : ClkMux
    port map (
            O => \N__10261\,
            I => \N__10136\
        );

    \I__2334\ : ClkMux
    port map (
            O => \N__10260\,
            I => \N__10136\
        );

    \I__2333\ : ClkMux
    port map (
            O => \N__10259\,
            I => \N__10136\
        );

    \I__2332\ : ClkMux
    port map (
            O => \N__10258\,
            I => \N__10136\
        );

    \I__2331\ : ClkMux
    port map (
            O => \N__10257\,
            I => \N__10136\
        );

    \I__2330\ : ClkMux
    port map (
            O => \N__10256\,
            I => \N__10136\
        );

    \I__2329\ : ClkMux
    port map (
            O => \N__10255\,
            I => \N__10136\
        );

    \I__2328\ : ClkMux
    port map (
            O => \N__10254\,
            I => \N__10136\
        );

    \I__2327\ : ClkMux
    port map (
            O => \N__10253\,
            I => \N__10136\
        );

    \I__2326\ : ClkMux
    port map (
            O => \N__10252\,
            I => \N__10136\
        );

    \I__2325\ : ClkMux
    port map (
            O => \N__10251\,
            I => \N__10136\
        );

    \I__2324\ : ClkMux
    port map (
            O => \N__10250\,
            I => \N__10136\
        );

    \I__2323\ : ClkMux
    port map (
            O => \N__10249\,
            I => \N__10136\
        );

    \I__2322\ : ClkMux
    port map (
            O => \N__10248\,
            I => \N__10136\
        );

    \I__2321\ : ClkMux
    port map (
            O => \N__10247\,
            I => \N__10136\
        );

    \I__2320\ : ClkMux
    port map (
            O => \N__10246\,
            I => \N__10136\
        );

    \I__2319\ : Glb2LocalMux
    port map (
            O => \N__10243\,
            I => \N__10136\
        );

    \I__2318\ : ClkMux
    port map (
            O => \N__10242\,
            I => \N__10136\
        );

    \I__2317\ : ClkMux
    port map (
            O => \N__10241\,
            I => \N__10136\
        );

    \I__2316\ : ClkMux
    port map (
            O => \N__10240\,
            I => \N__10136\
        );

    \I__2315\ : ClkMux
    port map (
            O => \N__10239\,
            I => \N__10136\
        );

    \I__2314\ : ClkMux
    port map (
            O => \N__10238\,
            I => \N__10136\
        );

    \I__2313\ : ClkMux
    port map (
            O => \N__10237\,
            I => \N__10136\
        );

    \I__2312\ : ClkMux
    port map (
            O => \N__10236\,
            I => \N__10136\
        );

    \I__2311\ : ClkMux
    port map (
            O => \N__10235\,
            I => \N__10136\
        );

    \I__2310\ : ClkMux
    port map (
            O => \N__10234\,
            I => \N__10136\
        );

    \I__2309\ : ClkMux
    port map (
            O => \N__10233\,
            I => \N__10136\
        );

    \I__2308\ : ClkMux
    port map (
            O => \N__10232\,
            I => \N__10136\
        );

    \I__2307\ : ClkMux
    port map (
            O => \N__10231\,
            I => \N__10136\
        );

    \I__2306\ : ClkMux
    port map (
            O => \N__10230\,
            I => \N__10136\
        );

    \I__2305\ : ClkMux
    port map (
            O => \N__10229\,
            I => \N__10136\
        );

    \I__2304\ : ClkMux
    port map (
            O => \N__10228\,
            I => \N__10136\
        );

    \I__2303\ : ClkMux
    port map (
            O => \N__10227\,
            I => \N__10136\
        );

    \I__2302\ : ClkMux
    port map (
            O => \N__10226\,
            I => \N__10136\
        );

    \I__2301\ : ClkMux
    port map (
            O => \N__10225\,
            I => \N__10136\
        );

    \I__2300\ : GlobalMux
    port map (
            O => \N__10136\,
            I => \CLK80_PLL\
        );

    \I__2299\ : InMux
    port map (
            O => \N__10133\,
            I => \N__10130\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__10130\,
            I => \N__10127\
        );

    \I__2297\ : Span4Mux_v
    port map (
            O => \N__10127\,
            I => \N__10123\
        );

    \I__2296\ : InMux
    port map (
            O => \N__10126\,
            I => \N__10120\
        );

    \I__2295\ : Sp12to4
    port map (
            O => \N__10123\,
            I => \N__10117\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__10120\,
            I => \N__10114\
        );

    \I__2293\ : Span12Mux_h
    port map (
            O => \N__10117\,
            I => \N__10107\
        );

    \I__2292\ : Span12Mux_h
    port map (
            O => \N__10114\,
            I => \N__10107\
        );

    \I__2291\ : InMux
    port map (
            O => \N__10113\,
            I => \N__10104\
        );

    \I__2290\ : InMux
    port map (
            O => \N__10112\,
            I => \N__10101\
        );

    \I__2289\ : Odrv12
    port map (
            O => \N__10107\,
            I => \REG_CYCLEm\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__10104\,
            I => \REG_CYCLEm\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__10101\,
            I => \REG_CYCLEm\
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__10094\,
            I => \N__10091\
        );

    \I__2285\ : InMux
    port map (
            O => \N__10091\,
            I => \N__10086\
        );

    \I__2284\ : CascadeMux
    port map (
            O => \N__10090\,
            I => \N__10083\
        );

    \I__2283\ : CascadeMux
    port map (
            O => \N__10089\,
            I => \N__10080\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__10086\,
            I => \N__10076\
        );

    \I__2281\ : InMux
    port map (
            O => \N__10083\,
            I => \N__10071\
        );

    \I__2280\ : InMux
    port map (
            O => \N__10080\,
            I => \N__10071\
        );

    \I__2279\ : CascadeMux
    port map (
            O => \N__10079\,
            I => \N__10066\
        );

    \I__2278\ : Span4Mux_v
    port map (
            O => \N__10076\,
            I => \N__10063\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__10071\,
            I => \N__10060\
        );

    \I__2276\ : InMux
    port map (
            O => \N__10070\,
            I => \N__10056\
        );

    \I__2275\ : InMux
    port map (
            O => \N__10069\,
            I => \N__10053\
        );

    \I__2274\ : InMux
    port map (
            O => \N__10066\,
            I => \N__10046\
        );

    \I__2273\ : Sp12to4
    port map (
            O => \N__10063\,
            I => \N__10043\
        );

    \I__2272\ : Span4Mux_v
    port map (
            O => \N__10060\,
            I => \N__10038\
        );

    \I__2271\ : InMux
    port map (
            O => \N__10059\,
            I => \N__10035\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__10056\,
            I => \N__10030\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__10053\,
            I => \N__10030\
        );

    \I__2268\ : InMux
    port map (
            O => \N__10052\,
            I => \N__10025\
        );

    \I__2267\ : InMux
    port map (
            O => \N__10051\,
            I => \N__10020\
        );

    \I__2266\ : InMux
    port map (
            O => \N__10050\,
            I => \N__10020\
        );

    \I__2265\ : InMux
    port map (
            O => \N__10049\,
            I => \N__10017\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__10046\,
            I => \N__10013\
        );

    \I__2263\ : Span12Mux_s9_h
    port map (
            O => \N__10043\,
            I => \N__10007\
        );

    \I__2262\ : InMux
    port map (
            O => \N__10042\,
            I => \N__10002\
        );

    \I__2261\ : InMux
    port map (
            O => \N__10041\,
            I => \N__10002\
        );

    \I__2260\ : Span4Mux_h
    port map (
            O => \N__10038\,
            I => \N__9994\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__10035\,
            I => \N__9994\
        );

    \I__2258\ : Span4Mux_v
    port map (
            O => \N__10030\,
            I => \N__9989\
        );

    \I__2257\ : InMux
    port map (
            O => \N__10029\,
            I => \N__9984\
        );

    \I__2256\ : InMux
    port map (
            O => \N__10028\,
            I => \N__9984\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__10025\,
            I => \N__9977\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__10020\,
            I => \N__9977\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__10017\,
            I => \N__9977\
        );

    \I__2252\ : InMux
    port map (
            O => \N__10016\,
            I => \N__9974\
        );

    \I__2251\ : Span4Mux_h
    port map (
            O => \N__10013\,
            I => \N__9971\
        );

    \I__2250\ : InMux
    port map (
            O => \N__10012\,
            I => \N__9964\
        );

    \I__2249\ : InMux
    port map (
            O => \N__10011\,
            I => \N__9964\
        );

    \I__2248\ : InMux
    port map (
            O => \N__10010\,
            I => \N__9964\
        );

    \I__2247\ : Span12Mux_v
    port map (
            O => \N__10007\,
            I => \N__9959\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__10002\,
            I => \N__9959\
        );

    \I__2245\ : InMux
    port map (
            O => \N__10001\,
            I => \N__9952\
        );

    \I__2244\ : InMux
    port map (
            O => \N__10000\,
            I => \N__9952\
        );

    \I__2243\ : InMux
    port map (
            O => \N__9999\,
            I => \N__9952\
        );

    \I__2242\ : Span4Mux_v
    port map (
            O => \N__9994\,
            I => \N__9949\
        );

    \I__2241\ : InMux
    port map (
            O => \N__9993\,
            I => \N__9944\
        );

    \I__2240\ : InMux
    port map (
            O => \N__9992\,
            I => \N__9944\
        );

    \I__2239\ : Span4Mux_v
    port map (
            O => \N__9989\,
            I => \N__9937\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__9984\,
            I => \N__9937\
        );

    \I__2237\ : Span4Mux_v
    port map (
            O => \N__9977\,
            I => \N__9937\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__9974\,
            I => \N__9934\
        );

    \I__2235\ : Odrv4
    port map (
            O => \N__9971\,
            I => \CPU_CYCLEm\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__9964\,
            I => \CPU_CYCLEm\
        );

    \I__2233\ : Odrv12
    port map (
            O => \N__9959\,
            I => \CPU_CYCLEm\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__9952\,
            I => \CPU_CYCLEm\
        );

    \I__2231\ : Odrv4
    port map (
            O => \N__9949\,
            I => \CPU_CYCLEm\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__9944\,
            I => \CPU_CYCLEm\
        );

    \I__2229\ : Odrv4
    port map (
            O => \N__9937\,
            I => \CPU_CYCLEm\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__9934\,
            I => \CPU_CYCLEm\
        );

    \I__2227\ : IoInMux
    port map (
            O => \N__9917\,
            I => \N__9914\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__9914\,
            I => \N__9911\
        );

    \I__2225\ : Span4Mux_s3_v
    port map (
            O => \N__9911\,
            I => \N__9908\
        );

    \I__2224\ : Span4Mux_v
    port map (
            O => \N__9908\,
            I => \N__9905\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__9905\,
            I => \N_136_i\
        );

    \I__2222\ : CascadeMux
    port map (
            O => \N__9902\,
            I => \N__9898\
        );

    \I__2221\ : InMux
    port map (
            O => \N__9901\,
            I => \N__9895\
        );

    \I__2220\ : InMux
    port map (
            O => \N__9898\,
            I => \N__9891\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__9895\,
            I => \N__9888\
        );

    \I__2218\ : InMux
    port map (
            O => \N__9894\,
            I => \N__9885\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__9891\,
            I => \N__9882\
        );

    \I__2216\ : Span4Mux_v
    port map (
            O => \N__9888\,
            I => \N__9879\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__9885\,
            I => \N__9876\
        );

    \I__2214\ : Span4Mux_v
    port map (
            O => \N__9882\,
            I => \N__9872\
        );

    \I__2213\ : Span4Mux_v
    port map (
            O => \N__9879\,
            I => \N__9867\
        );

    \I__2212\ : Span4Mux_h
    port map (
            O => \N__9876\,
            I => \N__9867\
        );

    \I__2211\ : CascadeMux
    port map (
            O => \N__9875\,
            I => \N__9864\
        );

    \I__2210\ : Span4Mux_v
    port map (
            O => \N__9872\,
            I => \N__9859\
        );

    \I__2209\ : Span4Mux_h
    port map (
            O => \N__9867\,
            I => \N__9859\
        );

    \I__2208\ : InMux
    port map (
            O => \N__9864\,
            I => \N__9854\
        );

    \I__2207\ : Span4Mux_h
    port map (
            O => \N__9859\,
            I => \N__9851\
        );

    \I__2206\ : InMux
    port map (
            O => \N__9858\,
            I => \N__9846\
        );

    \I__2205\ : InMux
    port map (
            O => \N__9857\,
            I => \N__9846\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__9854\,
            I => \N__9843\
        );

    \I__2203\ : Span4Mux_h
    port map (
            O => \N__9851\,
            I => \N__9838\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__9846\,
            I => \N__9838\
        );

    \I__2201\ : Span12Mux_v
    port map (
            O => \N__9843\,
            I => \N__9835\
        );

    \I__2200\ : Span4Mux_h
    port map (
            O => \N__9838\,
            I => \N__9832\
        );

    \I__2199\ : Span12Mux_h
    port map (
            O => \N__9835\,
            I => \N__9829\
        );

    \I__2198\ : Span4Mux_v
    port map (
            O => \N__9832\,
            I => \N__9826\
        );

    \I__2197\ : Odrv12
    port map (
            O => \N__9829\,
            I => \CASUn_c\
        );

    \I__2196\ : Odrv4
    port map (
            O => \N__9826\,
            I => \CASUn_c\
        );

    \I__2195\ : InMux
    port map (
            O => \N__9821\,
            I => \N__9817\
        );

    \I__2194\ : InMux
    port map (
            O => \N__9820\,
            I => \N__9814\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__9817\,
            I => \N__9811\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__9814\,
            I => \N__9805\
        );

    \I__2191\ : Span4Mux_v
    port map (
            O => \N__9811\,
            I => \N__9802\
        );

    \I__2190\ : InMux
    port map (
            O => \N__9810\,
            I => \N__9799\
        );

    \I__2189\ : CascadeMux
    port map (
            O => \N__9809\,
            I => \N__9796\
        );

    \I__2188\ : InMux
    port map (
            O => \N__9808\,
            I => \N__9793\
        );

    \I__2187\ : Span4Mux_v
    port map (
            O => \N__9805\,
            I => \N__9790\
        );

    \I__2186\ : Span4Mux_v
    port map (
            O => \N__9802\,
            I => \N__9785\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__9799\,
            I => \N__9785\
        );

    \I__2184\ : InMux
    port map (
            O => \N__9796\,
            I => \N__9782\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__9793\,
            I => \N__9779\
        );

    \I__2182\ : Sp12to4
    port map (
            O => \N__9790\,
            I => \N__9776\
        );

    \I__2181\ : Span4Mux_v
    port map (
            O => \N__9785\,
            I => \N__9773\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__9782\,
            I => \N__9768\
        );

    \I__2179\ : Sp12to4
    port map (
            O => \N__9779\,
            I => \N__9768\
        );

    \I__2178\ : Span12Mux_h
    port map (
            O => \N__9776\,
            I => \N__9763\
        );

    \I__2177\ : Sp12to4
    port map (
            O => \N__9773\,
            I => \N__9763\
        );

    \I__2176\ : Span12Mux_v
    port map (
            O => \N__9768\,
            I => \N__9760\
        );

    \I__2175\ : Span12Mux_h
    port map (
            O => \N__9763\,
            I => \N__9757\
        );

    \I__2174\ : Span12Mux_h
    port map (
            O => \N__9760\,
            I => \N__9754\
        );

    \I__2173\ : Odrv12
    port map (
            O => \N__9757\,
            I => \RnW_c\
        );

    \I__2172\ : Odrv12
    port map (
            O => \N__9754\,
            I => \RnW_c\
        );

    \I__2171\ : InMux
    port map (
            O => \N__9749\,
            I => \N__9741\
        );

    \I__2170\ : InMux
    port map (
            O => \N__9748\,
            I => \N__9741\
        );

    \I__2169\ : InMux
    port map (
            O => \N__9747\,
            I => \N__9736\
        );

    \I__2168\ : InMux
    port map (
            O => \N__9746\,
            I => \N__9736\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__9741\,
            I => \N__9733\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__9736\,
            I => \N__9730\
        );

    \I__2165\ : Span4Mux_v
    port map (
            O => \N__9733\,
            I => \N__9727\
        );

    \I__2164\ : Span4Mux_v
    port map (
            O => \N__9730\,
            I => \N__9724\
        );

    \I__2163\ : Sp12to4
    port map (
            O => \N__9727\,
            I => \N__9721\
        );

    \I__2162\ : Span4Mux_h
    port map (
            O => \N__9724\,
            I => \N__9718\
        );

    \I__2161\ : Span12Mux_h
    port map (
            O => \N__9721\,
            I => \N__9713\
        );

    \I__2160\ : Sp12to4
    port map (
            O => \N__9718\,
            I => \N__9713\
        );

    \I__2159\ : Odrv12
    port map (
            O => \N__9713\,
            I => \DRA_c_7\
        );

    \I__2158\ : InMux
    port map (
            O => \N__9710\,
            I => \N__9705\
        );

    \I__2157\ : InMux
    port map (
            O => \N__9709\,
            I => \N__9700\
        );

    \I__2156\ : InMux
    port map (
            O => \N__9708\,
            I => \N__9700\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__9705\,
            I => \N__9694\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__9700\,
            I => \N__9694\
        );

    \I__2153\ : InMux
    port map (
            O => \N__9699\,
            I => \N__9691\
        );

    \I__2152\ : Sp12to4
    port map (
            O => \N__9694\,
            I => \N__9686\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__9691\,
            I => \N__9686\
        );

    \I__2150\ : Span12Mux_v
    port map (
            O => \N__9686\,
            I => \N__9683\
        );

    \I__2149\ : Span12Mux_h
    port map (
            O => \N__9683\,
            I => \N__9680\
        );

    \I__2148\ : Odrv12
    port map (
            O => \N__9680\,
            I => \DRA_c_6\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9677\,
            I => \N__9674\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__9674\,
            I => \N__9671\
        );

    \I__2145\ : Odrv4
    port map (
            O => \N__9671\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2144\ : InMux
    port map (
            O => \N__9668\,
            I => \N__9665\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__9665\,
            I => \N__9662\
        );

    \I__2142\ : Span4Mux_h
    port map (
            O => \N__9662\,
            I => \N__9659\
        );

    \I__2141\ : Odrv4
    port map (
            O => \N__9659\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__2140\ : InMux
    port map (
            O => \N__9656\,
            I => \N__9652\
        );

    \I__2139\ : InMux
    port map (
            O => \N__9655\,
            I => \N__9647\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__9652\,
            I => \N__9644\
        );

    \I__2137\ : InMux
    port map (
            O => \N__9651\,
            I => \N__9641\
        );

    \I__2136\ : InMux
    port map (
            O => \N__9650\,
            I => \N__9638\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__9647\,
            I => \N__9635\
        );

    \I__2134\ : Span4Mux_h
    port map (
            O => \N__9644\,
            I => \N__9628\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__9641\,
            I => \N__9628\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__9638\,
            I => \N__9628\
        );

    \I__2131\ : Span4Mux_v
    port map (
            O => \N__9635\,
            I => \N__9625\
        );

    \I__2130\ : Span4Mux_v
    port map (
            O => \N__9628\,
            I => \N__9622\
        );

    \I__2129\ : Sp12to4
    port map (
            O => \N__9625\,
            I => \N__9619\
        );

    \I__2128\ : Span4Mux_v
    port map (
            O => \N__9622\,
            I => \N__9616\
        );

    \I__2127\ : Span12Mux_h
    port map (
            O => \N__9619\,
            I => \N__9613\
        );

    \I__2126\ : Sp12to4
    port map (
            O => \N__9616\,
            I => \N__9610\
        );

    \I__2125\ : Span12Mux_v
    port map (
            O => \N__9613\,
            I => \N__9607\
        );

    \I__2124\ : Span12Mux_h
    port map (
            O => \N__9610\,
            I => \N__9604\
        );

    \I__2123\ : Odrv12
    port map (
            O => \N__9607\,
            I => \DRA_c_4\
        );

    \I__2122\ : Odrv12
    port map (
            O => \N__9604\,
            I => \DRA_c_4\
        );

    \I__2121\ : InMux
    port map (
            O => \N__9599\,
            I => \N__9596\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__9596\,
            I => \N__9590\
        );

    \I__2119\ : InMux
    port map (
            O => \N__9595\,
            I => \N__9587\
        );

    \I__2118\ : InMux
    port map (
            O => \N__9594\,
            I => \N__9584\
        );

    \I__2117\ : InMux
    port map (
            O => \N__9593\,
            I => \N__9581\
        );

    \I__2116\ : Sp12to4
    port map (
            O => \N__9590\,
            I => \N__9572\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__9587\,
            I => \N__9572\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__9584\,
            I => \N__9572\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__9581\,
            I => \N__9572\
        );

    \I__2112\ : Span12Mux_v
    port map (
            O => \N__9572\,
            I => \N__9569\
        );

    \I__2111\ : Span12Mux_h
    port map (
            O => \N__9569\,
            I => \N__9566\
        );

    \I__2110\ : Odrv12
    port map (
            O => \N__9566\,
            I => \DRA_c_3\
        );

    \I__2109\ : InMux
    port map (
            O => \N__9563\,
            I => \N__9560\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__9560\,
            I => \N__9557\
        );

    \I__2107\ : Span4Mux_h
    port map (
            O => \N__9557\,
            I => \N__9554\
        );

    \I__2106\ : Odrv4
    port map (
            O => \N__9554\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2105\ : IoInMux
    port map (
            O => \N__9551\,
            I => \N__9548\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__9548\,
            I => \N__9545\
        );

    \I__2103\ : Span4Mux_s2_h
    port map (
            O => \N__9545\,
            I => \N__9542\
        );

    \I__2102\ : Sp12to4
    port map (
            O => \N__9542\,
            I => \N__9539\
        );

    \I__2101\ : Span12Mux_v
    port map (
            O => \N__9539\,
            I => \N__9536\
        );

    \I__2100\ : Span12Mux_h
    port map (
            O => \N__9536\,
            I => \N__9533\
        );

    \I__2099\ : Odrv12
    port map (
            O => \N__9533\,
            I => \N_146_i\
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__9530\,
            I => \N__9524\
        );

    \I__2097\ : InMux
    port map (
            O => \N__9529\,
            I => \N__9521\
        );

    \I__2096\ : InMux
    port map (
            O => \N__9528\,
            I => \N__9516\
        );

    \I__2095\ : InMux
    port map (
            O => \N__9527\,
            I => \N__9516\
        );

    \I__2094\ : InMux
    port map (
            O => \N__9524\,
            I => \N__9513\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__9521\,
            I => \N__9510\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__9516\,
            I => \N__9505\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__9513\,
            I => \N__9505\
        );

    \I__2090\ : Span4Mux_v
    port map (
            O => \N__9510\,
            I => \N__9502\
        );

    \I__2089\ : Span4Mux_v
    port map (
            O => \N__9505\,
            I => \N__9499\
        );

    \I__2088\ : Sp12to4
    port map (
            O => \N__9502\,
            I => \N__9496\
        );

    \I__2087\ : Span4Mux_h
    port map (
            O => \N__9499\,
            I => \N__9493\
        );

    \I__2086\ : Span12Mux_h
    port map (
            O => \N__9496\,
            I => \N__9488\
        );

    \I__2085\ : Sp12to4
    port map (
            O => \N__9493\,
            I => \N__9488\
        );

    \I__2084\ : Span12Mux_v
    port map (
            O => \N__9488\,
            I => \N__9485\
        );

    \I__2083\ : Odrv12
    port map (
            O => \N__9485\,
            I => \CLK40_PLL_i\
        );

    \I__2082\ : IoInMux
    port map (
            O => \N__9482\,
            I => \N__9478\
        );

    \I__2081\ : IoInMux
    port map (
            O => \N__9481\,
            I => \N__9475\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__9478\,
            I => \N__9472\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__9475\,
            I => \N__9468\
        );

    \I__2078\ : Span4Mux_s2_v
    port map (
            O => \N__9472\,
            I => \N__9465\
        );

    \I__2077\ : IoInMux
    port map (
            O => \N__9471\,
            I => \N__9462\
        );

    \I__2076\ : IoSpan4Mux
    port map (
            O => \N__9468\,
            I => \N__9459\
        );

    \I__2075\ : Sp12to4
    port map (
            O => \N__9465\,
            I => \N__9456\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__9462\,
            I => \N__9453\
        );

    \I__2073\ : Span4Mux_s2_h
    port map (
            O => \N__9459\,
            I => \N__9450\
        );

    \I__2072\ : Span12Mux_h
    port map (
            O => \N__9456\,
            I => \N__9447\
        );

    \I__2071\ : Span12Mux_s2_v
    port map (
            O => \N__9453\,
            I => \N__9444\
        );

    \I__2070\ : Sp12to4
    port map (
            O => \N__9450\,
            I => \N__9441\
        );

    \I__2069\ : Span12Mux_v
    port map (
            O => \N__9447\,
            I => \N__9436\
        );

    \I__2068\ : Span12Mux_v
    port map (
            O => \N__9444\,
            I => \N__9436\
        );

    \I__2067\ : Span12Mux_s8_h
    port map (
            O => \N__9441\,
            I => \N__9433\
        );

    \I__2066\ : Odrv12
    port map (
            O => \N__9436\,
            I => \CLK40_PLL_i_i\
        );

    \I__2065\ : Odrv12
    port map (
            O => \N__9433\,
            I => \CLK40_PLL_i_i\
        );

    \I__2064\ : InMux
    port map (
            O => \N__9428\,
            I => \N__9425\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__9425\,
            I => \U712_BYTE_ENABLE.N_406\
        );

    \I__2062\ : InMux
    port map (
            O => \N__9422\,
            I => \N__9416\
        );

    \I__2061\ : InMux
    port map (
            O => \N__9421\,
            I => \N__9416\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__9416\,
            I => \U712_BYTE_ENABLE.N_284_i\
        );

    \I__2059\ : IoInMux
    port map (
            O => \N__9413\,
            I => \N__9410\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__9410\,
            I => \N__9407\
        );

    \I__2057\ : IoSpan4Mux
    port map (
            O => \N__9407\,
            I => \N__9404\
        );

    \I__2056\ : Span4Mux_s2_v
    port map (
            O => \N__9404\,
            I => \N__9401\
        );

    \I__2055\ : Span4Mux_v
    port map (
            O => \N__9401\,
            I => \N__9398\
        );

    \I__2054\ : Odrv4
    port map (
            O => \N__9398\,
            I => \N_374_i\
        );

    \I__2053\ : CascadeMux
    port map (
            O => \N__9395\,
            I => \N__9392\
        );

    \I__2052\ : InMux
    port map (
            O => \N__9392\,
            I => \N__9388\
        );

    \I__2051\ : InMux
    port map (
            O => \N__9391\,
            I => \N__9385\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__9388\,
            I => \U712_BYTE_ENABLE.N_409\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__9385\,
            I => \U712_BYTE_ENABLE.N_409\
        );

    \I__2048\ : CascadeMux
    port map (
            O => \N__9380\,
            I => \N__9374\
        );

    \I__2047\ : CascadeMux
    port map (
            O => \N__9379\,
            I => \N__9371\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__9378\,
            I => \N__9366\
        );

    \I__2045\ : InMux
    port map (
            O => \N__9377\,
            I => \N__9356\
        );

    \I__2044\ : InMux
    port map (
            O => \N__9374\,
            I => \N__9356\
        );

    \I__2043\ : InMux
    port map (
            O => \N__9371\,
            I => \N__9356\
        );

    \I__2042\ : InMux
    port map (
            O => \N__9370\,
            I => \N__9353\
        );

    \I__2041\ : InMux
    port map (
            O => \N__9369\,
            I => \N__9349\
        );

    \I__2040\ : InMux
    port map (
            O => \N__9366\,
            I => \N__9346\
        );

    \I__2039\ : CascadeMux
    port map (
            O => \N__9365\,
            I => \N__9342\
        );

    \I__2038\ : InMux
    port map (
            O => \N__9364\,
            I => \N__9339\
        );

    \I__2037\ : InMux
    port map (
            O => \N__9363\,
            I => \N__9336\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__9356\,
            I => \N__9331\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__9353\,
            I => \N__9331\
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__9352\,
            I => \N__9328\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__9349\,
            I => \N__9322\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__9346\,
            I => \N__9319\
        );

    \I__2031\ : InMux
    port map (
            O => \N__9345\,
            I => \N__9316\
        );

    \I__2030\ : InMux
    port map (
            O => \N__9342\,
            I => \N__9313\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__9339\,
            I => \N__9310\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__9336\,
            I => \N__9307\
        );

    \I__2027\ : Span4Mux_h
    port map (
            O => \N__9331\,
            I => \N__9304\
        );

    \I__2026\ : InMux
    port map (
            O => \N__9328\,
            I => \N__9301\
        );

    \I__2025\ : InMux
    port map (
            O => \N__9327\,
            I => \N__9298\
        );

    \I__2024\ : InMux
    port map (
            O => \N__9326\,
            I => \N__9295\
        );

    \I__2023\ : InMux
    port map (
            O => \N__9325\,
            I => \N__9292\
        );

    \I__2022\ : Span4Mux_v
    port map (
            O => \N__9322\,
            I => \N__9285\
        );

    \I__2021\ : Span4Mux_v
    port map (
            O => \N__9319\,
            I => \N__9285\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__9316\,
            I => \N__9285\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__9313\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2018\ : Odrv4
    port map (
            O => \N__9310\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2017\ : Odrv12
    port map (
            O => \N__9307\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2016\ : Odrv4
    port map (
            O => \N__9304\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__9301\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__9298\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__9295\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__9292\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2011\ : Odrv4
    port map (
            O => \N__9285\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2010\ : IoInMux
    port map (
            O => \N__9266\,
            I => \N__9263\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__9263\,
            I => \N__9260\
        );

    \I__2008\ : Span12Mux_s4_v
    port map (
            O => \N__9260\,
            I => \N__9257\
        );

    \I__2007\ : Span12Mux_h
    port map (
            O => \N__9257\,
            I => \N__9254\
        );

    \I__2006\ : Odrv12
    port map (
            O => \N__9254\,
            I => \ASn_c\
        );

    \I__2005\ : CEMux
    port map (
            O => \N__9251\,
            I => \N__9248\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__9248\,
            I => \N__9245\
        );

    \I__2003\ : Odrv4
    port map (
            O => \N__9245\,
            I => \U712_REG_SM.N_95_0\
        );

    \I__2002\ : IoInMux
    port map (
            O => \N__9242\,
            I => \N__9239\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__9239\,
            I => \N__9236\
        );

    \I__2000\ : Span4Mux_s2_v
    port map (
            O => \N__9236\,
            I => \N__9233\
        );

    \I__1999\ : Span4Mux_v
    port map (
            O => \N__9233\,
            I => \N__9230\
        );

    \I__1998\ : Odrv4
    port map (
            O => \N__9230\,
            I => \LLBEn_c\
        );

    \I__1997\ : InMux
    port map (
            O => \N__9227\,
            I => \N__9221\
        );

    \I__1996\ : CascadeMux
    port map (
            O => \N__9226\,
            I => \N__9211\
        );

    \I__1995\ : CascadeMux
    port map (
            O => \N__9225\,
            I => \N__9206\
        );

    \I__1994\ : InMux
    port map (
            O => \N__9224\,
            I => \N__9203\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__9221\,
            I => \N__9200\
        );

    \I__1992\ : InMux
    port map (
            O => \N__9220\,
            I => \N__9197\
        );

    \I__1991\ : InMux
    port map (
            O => \N__9219\,
            I => \N__9186\
        );

    \I__1990\ : InMux
    port map (
            O => \N__9218\,
            I => \N__9186\
        );

    \I__1989\ : InMux
    port map (
            O => \N__9217\,
            I => \N__9186\
        );

    \I__1988\ : InMux
    port map (
            O => \N__9216\,
            I => \N__9186\
        );

    \I__1987\ : InMux
    port map (
            O => \N__9215\,
            I => \N__9186\
        );

    \I__1986\ : InMux
    port map (
            O => \N__9214\,
            I => \N__9183\
        );

    \I__1985\ : InMux
    port map (
            O => \N__9211\,
            I => \N__9180\
        );

    \I__1984\ : CascadeMux
    port map (
            O => \N__9210\,
            I => \N__9177\
        );

    \I__1983\ : CascadeMux
    port map (
            O => \N__9209\,
            I => \N__9174\
        );

    \I__1982\ : InMux
    port map (
            O => \N__9206\,
            I => \N__9170\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__9203\,
            I => \N__9153\
        );

    \I__1980\ : Span4Mux_h
    port map (
            O => \N__9200\,
            I => \N__9153\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__9197\,
            I => \N__9153\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__9186\,
            I => \N__9153\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__9183\,
            I => \N__9145\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__9180\,
            I => \N__9145\
        );

    \I__1975\ : InMux
    port map (
            O => \N__9177\,
            I => \N__9138\
        );

    \I__1974\ : InMux
    port map (
            O => \N__9174\,
            I => \N__9138\
        );

    \I__1973\ : InMux
    port map (
            O => \N__9173\,
            I => \N__9138\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__9170\,
            I => \N__9134\
        );

    \I__1971\ : InMux
    port map (
            O => \N__9169\,
            I => \N__9125\
        );

    \I__1970\ : InMux
    port map (
            O => \N__9168\,
            I => \N__9125\
        );

    \I__1969\ : InMux
    port map (
            O => \N__9167\,
            I => \N__9125\
        );

    \I__1968\ : InMux
    port map (
            O => \N__9166\,
            I => \N__9125\
        );

    \I__1967\ : InMux
    port map (
            O => \N__9165\,
            I => \N__9116\
        );

    \I__1966\ : InMux
    port map (
            O => \N__9164\,
            I => \N__9116\
        );

    \I__1965\ : InMux
    port map (
            O => \N__9163\,
            I => \N__9116\
        );

    \I__1964\ : InMux
    port map (
            O => \N__9162\,
            I => \N__9116\
        );

    \I__1963\ : Span4Mux_h
    port map (
            O => \N__9153\,
            I => \N__9113\
        );

    \I__1962\ : InMux
    port map (
            O => \N__9152\,
            I => \N__9106\
        );

    \I__1961\ : InMux
    port map (
            O => \N__9151\,
            I => \N__9106\
        );

    \I__1960\ : InMux
    port map (
            O => \N__9150\,
            I => \N__9106\
        );

    \I__1959\ : Span4Mux_h
    port map (
            O => \N__9145\,
            I => \N__9101\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__9138\,
            I => \N__9101\
        );

    \I__1957\ : InMux
    port map (
            O => \N__9137\,
            I => \N__9098\
        );

    \I__1956\ : Odrv4
    port map (
            O => \N__9134\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__9125\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__9116\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1953\ : Odrv4
    port map (
            O => \N__9113\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__9106\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__9101\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__9098\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1949\ : IoInMux
    port map (
            O => \N__9083\,
            I => \N__9080\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__9080\,
            I => \N__9077\
        );

    \I__1947\ : Span4Mux_s3_v
    port map (
            O => \N__9077\,
            I => \N__9074\
        );

    \I__1946\ : Sp12to4
    port map (
            O => \N__9074\,
            I => \N__9071\
        );

    \I__1945\ : Span12Mux_h
    port map (
            O => \N__9071\,
            I => \N__9068\
        );

    \I__1944\ : Odrv12
    port map (
            O => \N__9068\,
            I => \CASn_c\
        );

    \I__1943\ : InMux
    port map (
            O => \N__9065\,
            I => \N__9059\
        );

    \I__1942\ : InMux
    port map (
            O => \N__9064\,
            I => \N__9056\
        );

    \I__1941\ : InMux
    port map (
            O => \N__9063\,
            I => \N__9051\
        );

    \I__1940\ : InMux
    port map (
            O => \N__9062\,
            I => \N__9051\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__9059\,
            I => \N__9044\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__9056\,
            I => \N__9044\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__9051\,
            I => \N__9044\
        );

    \I__1936\ : Sp12to4
    port map (
            O => \N__9044\,
            I => \N__9041\
        );

    \I__1935\ : Span12Mux_v
    port map (
            O => \N__9041\,
            I => \N__9038\
        );

    \I__1934\ : Span12Mux_h
    port map (
            O => \N__9038\,
            I => \N__9035\
        );

    \I__1933\ : Odrv12
    port map (
            O => \N__9035\,
            I => \DRA_c_5\
        );

    \I__1932\ : InMux
    port map (
            O => \N__9032\,
            I => \N__9029\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__9029\,
            I => \N__9026\
        );

    \I__1930\ : Odrv12
    port map (
            O => \N__9026\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__1929\ : InMux
    port map (
            O => \N__9023\,
            I => \N__9017\
        );

    \I__1928\ : InMux
    port map (
            O => \N__9022\,
            I => \N__9017\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__9017\,
            I => \N__9013\
        );

    \I__1926\ : InMux
    port map (
            O => \N__9016\,
            I => \N__9010\
        );

    \I__1925\ : Span4Mux_h
    port map (
            O => \N__9013\,
            I => \N__9004\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__9010\,
            I => \N__9004\
        );

    \I__1923\ : InMux
    port map (
            O => \N__9009\,
            I => \N__9001\
        );

    \I__1922\ : Span4Mux_h
    port map (
            O => \N__9004\,
            I => \N__8996\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__9001\,
            I => \N__8996\
        );

    \I__1920\ : Sp12to4
    port map (
            O => \N__8996\,
            I => \N__8993\
        );

    \I__1919\ : Span12Mux_v
    port map (
            O => \N__8993\,
            I => \N__8990\
        );

    \I__1918\ : Span12Mux_h
    port map (
            O => \N__8990\,
            I => \N__8987\
        );

    \I__1917\ : Odrv12
    port map (
            O => \N__8987\,
            I => \DRA_c_2\
        );

    \I__1916\ : CascadeMux
    port map (
            O => \N__8984\,
            I => \N__8981\
        );

    \I__1915\ : InMux
    port map (
            O => \N__8981\,
            I => \N__8978\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__8978\,
            I => \N__8975\
        );

    \I__1913\ : Span4Mux_v
    port map (
            O => \N__8975\,
            I => \N__8972\
        );

    \I__1912\ : Odrv4
    port map (
            O => \N__8972\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__1911\ : CascadeMux
    port map (
            O => \N__8969\,
            I => \N__8964\
        );

    \I__1910\ : InMux
    port map (
            O => \N__8968\,
            I => \N__8959\
        );

    \I__1909\ : InMux
    port map (
            O => \N__8967\,
            I => \N__8959\
        );

    \I__1908\ : InMux
    port map (
            O => \N__8964\,
            I => \N__8956\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__8959\,
            I => \N__8952\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__8956\,
            I => \N__8949\
        );

    \I__1905\ : InMux
    port map (
            O => \N__8955\,
            I => \N__8946\
        );

    \I__1904\ : Span4Mux_h
    port map (
            O => \N__8952\,
            I => \N__8939\
        );

    \I__1903\ : Span4Mux_v
    port map (
            O => \N__8949\,
            I => \N__8939\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__8946\,
            I => \N__8939\
        );

    \I__1901\ : Span4Mux_h
    port map (
            O => \N__8939\,
            I => \N__8936\
        );

    \I__1900\ : Sp12to4
    port map (
            O => \N__8936\,
            I => \N__8933\
        );

    \I__1899\ : Span12Mux_v
    port map (
            O => \N__8933\,
            I => \N__8930\
        );

    \I__1898\ : Odrv12
    port map (
            O => \N__8930\,
            I => \DRA_c_1\
        );

    \I__1897\ : InMux
    port map (
            O => \N__8927\,
            I => \N__8923\
        );

    \I__1896\ : InMux
    port map (
            O => \N__8926\,
            I => \N__8920\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__8923\,
            I => \N__8917\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__8920\,
            I => \N__8914\
        );

    \I__1893\ : Span4Mux_v
    port map (
            O => \N__8917\,
            I => \N__8911\
        );

    \I__1892\ : Span4Mux_v
    port map (
            O => \N__8914\,
            I => \N__8908\
        );

    \I__1891\ : Sp12to4
    port map (
            O => \N__8911\,
            I => \N__8905\
        );

    \I__1890\ : Sp12to4
    port map (
            O => \N__8908\,
            I => \N__8902\
        );

    \I__1889\ : Span12Mux_h
    port map (
            O => \N__8905\,
            I => \N__8899\
        );

    \I__1888\ : Span12Mux_h
    port map (
            O => \N__8902\,
            I => \N__8896\
        );

    \I__1887\ : Span12Mux_v
    port map (
            O => \N__8899\,
            I => \N__8893\
        );

    \I__1886\ : Span12Mux_v
    port map (
            O => \N__8896\,
            I => \N__8890\
        );

    \I__1885\ : Odrv12
    port map (
            O => \N__8893\,
            I => \DRA_c_0\
        );

    \I__1884\ : Odrv12
    port map (
            O => \N__8890\,
            I => \DRA_c_0\
        );

    \I__1883\ : InMux
    port map (
            O => \N__8885\,
            I => \N__8882\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__8882\,
            I => \N__8879\
        );

    \I__1881\ : Span4Mux_v
    port map (
            O => \N__8879\,
            I => \N__8876\
        );

    \I__1880\ : Odrv4
    port map (
            O => \N__8876\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__1879\ : InMux
    port map (
            O => \N__8873\,
            I => \N__8868\
        );

    \I__1878\ : InMux
    port map (
            O => \N__8872\,
            I => \N__8865\
        );

    \I__1877\ : InMux
    port map (
            O => \N__8871\,
            I => \N__8862\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__8868\,
            I => \N__8857\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__8865\,
            I => \N__8857\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__8862\,
            I => \N__8854\
        );

    \I__1873\ : Span4Mux_v
    port map (
            O => \N__8857\,
            I => \N__8850\
        );

    \I__1872\ : Span4Mux_v
    port map (
            O => \N__8854\,
            I => \N__8847\
        );

    \I__1871\ : InMux
    port map (
            O => \N__8853\,
            I => \N__8844\
        );

    \I__1870\ : Sp12to4
    port map (
            O => \N__8850\,
            I => \N__8837\
        );

    \I__1869\ : Sp12to4
    port map (
            O => \N__8847\,
            I => \N__8837\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__8844\,
            I => \N__8837\
        );

    \I__1867\ : Span12Mux_h
    port map (
            O => \N__8837\,
            I => \N__8834\
        );

    \I__1866\ : Odrv12
    port map (
            O => \N__8834\,
            I => \DRA_c_8\
        );

    \I__1865\ : InMux
    port map (
            O => \N__8831\,
            I => \N__8828\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__8828\,
            I => \N__8825\
        );

    \I__1863\ : Odrv12
    port map (
            O => \N__8825\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__1862\ : InMux
    port map (
            O => \N__8822\,
            I => \N__8819\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__8819\,
            I => \N__8816\
        );

    \I__1860\ : Span4Mux_h
    port map (
            O => \N__8816\,
            I => \N__8813\
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__8813\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__1858\ : InMux
    port map (
            O => \N__8810\,
            I => \N__8807\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__8807\,
            I => \N__8804\
        );

    \I__1856\ : Odrv4
    port map (
            O => \N__8804\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__1855\ : InMux
    port map (
            O => \N__8801\,
            I => \N__8798\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__8798\,
            I => \N__8795\
        );

    \I__1853\ : Odrv4
    port map (
            O => \N__8795\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__1852\ : InMux
    port map (
            O => \N__8792\,
            I => \N__8789\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__8789\,
            I => \N__8786\
        );

    \I__1850\ : Span4Mux_h
    port map (
            O => \N__8786\,
            I => \N__8783\
        );

    \I__1849\ : Odrv4
    port map (
            O => \N__8783\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__1848\ : InMux
    port map (
            O => \N__8780\,
            I => \N__8777\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__8777\,
            I => \N__8774\
        );

    \I__1846\ : Span4Mux_h
    port map (
            O => \N__8774\,
            I => \N__8771\
        );

    \I__1845\ : Odrv4
    port map (
            O => \N__8771\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1844\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8762\
        );

    \I__1843\ : InMux
    port map (
            O => \N__8767\,
            I => \N__8762\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__8762\,
            I => \N__8759\
        );

    \I__1841\ : Span4Mux_h
    port map (
            O => \N__8759\,
            I => \N__8756\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__8756\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8753\,
            I => \N__8750\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__8750\,
            I => \N__8747\
        );

    \I__1837\ : Span4Mux_v
    port map (
            O => \N__8747\,
            I => \N__8744\
        );

    \I__1836\ : Odrv4
    port map (
            O => \N__8744\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8741\,
            I => \N__8738\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__8738\,
            I => \N__8735\
        );

    \I__1833\ : Span4Mux_h
    port map (
            O => \N__8735\,
            I => \N__8732\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__8732\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__1831\ : InMux
    port map (
            O => \N__8729\,
            I => \N__8726\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8726\,
            I => \N__8722\
        );

    \I__1829\ : InMux
    port map (
            O => \N__8725\,
            I => \N__8719\
        );

    \I__1828\ : Span4Mux_h
    port map (
            O => \N__8722\,
            I => \N__8716\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8719\,
            I => \N__8713\
        );

    \I__1826\ : Span4Mux_v
    port map (
            O => \N__8716\,
            I => \N__8710\
        );

    \I__1825\ : Span4Mux_v
    port map (
            O => \N__8713\,
            I => \N__8707\
        );

    \I__1824\ : Odrv4
    port map (
            O => \N__8710\,
            I => \DBRn_c_i\
        );

    \I__1823\ : Odrv4
    port map (
            O => \N__8707\,
            I => \DBRn_c_i\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8702\,
            I => \N__8699\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__8699\,
            I => \N__8695\
        );

    \I__1820\ : InMux
    port map (
            O => \N__8698\,
            I => \N__8692\
        );

    \I__1819\ : Span4Mux_h
    port map (
            O => \N__8695\,
            I => \N__8689\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__8692\,
            I => \N__8684\
        );

    \I__1817\ : Span4Mux_v
    port map (
            O => \N__8689\,
            I => \N__8684\
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__8684\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8681\,
            I => \N__8675\
        );

    \I__1814\ : InMux
    port map (
            O => \N__8680\,
            I => \N__8675\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__8675\,
            I => \U712_REG_SM.N_95\
        );

    \I__1812\ : IoInMux
    port map (
            O => \N__8672\,
            I => \N__8669\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__8669\,
            I => \N__8666\
        );

    \I__1810\ : Span4Mux_s3_v
    port map (
            O => \N__8666\,
            I => \N__8663\
        );

    \I__1809\ : Span4Mux_v
    port map (
            O => \N__8663\,
            I => \N__8660\
        );

    \I__1808\ : Span4Mux_v
    port map (
            O => \N__8660\,
            I => \N__8656\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__8659\,
            I => \N__8653\
        );

    \I__1806\ : Sp12to4
    port map (
            O => \N__8656\,
            I => \N__8650\
        );

    \I__1805\ : InMux
    port map (
            O => \N__8653\,
            I => \N__8647\
        );

    \I__1804\ : Odrv12
    port map (
            O => \N__8650\,
            I => \UDSn_c\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__8647\,
            I => \UDSn_c\
        );

    \I__1802\ : InMux
    port map (
            O => \N__8642\,
            I => \N__8639\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__8639\,
            I => \U712_REG_SM.N_433\
        );

    \I__1800\ : IoInMux
    port map (
            O => \N__8636\,
            I => \N__8633\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__8633\,
            I => \N__8630\
        );

    \I__1798\ : Odrv12
    port map (
            O => \N__8630\,
            I => \RESETn_c_i\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__8627\,
            I => \N__8624\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8624\,
            I => \N__8621\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__8621\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1794\ : IoInMux
    port map (
            O => \N__8618\,
            I => \N__8615\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__8615\,
            I => \N__8612\
        );

    \I__1792\ : Span12Mux_s3_h
    port map (
            O => \N__8612\,
            I => \N__8609\
        );

    \I__1791\ : Span12Mux_h
    port map (
            O => \N__8609\,
            I => \N__8606\
        );

    \I__1790\ : Odrv12
    port map (
            O => \N__8606\,
            I => \CMA_c_3\
        );

    \I__1789\ : InMux
    port map (
            O => \N__8603\,
            I => \N__8600\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__8600\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__1787\ : IoInMux
    port map (
            O => \N__8597\,
            I => \N__8594\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__8594\,
            I => \N__8591\
        );

    \I__1785\ : Span12Mux_s3_h
    port map (
            O => \N__8591\,
            I => \N__8588\
        );

    \I__1784\ : Span12Mux_h
    port map (
            O => \N__8588\,
            I => \N__8585\
        );

    \I__1783\ : Odrv12
    port map (
            O => \N__8585\,
            I => \CMA_c_4\
        );

    \I__1782\ : InMux
    port map (
            O => \N__8582\,
            I => \N__8577\
        );

    \I__1781\ : InMux
    port map (
            O => \N__8581\,
            I => \N__8572\
        );

    \I__1780\ : InMux
    port map (
            O => \N__8580\,
            I => \N__8572\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__8577\,
            I => \N__8564\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__8572\,
            I => \N__8564\
        );

    \I__1777\ : InMux
    port map (
            O => \N__8571\,
            I => \N__8557\
        );

    \I__1776\ : InMux
    port map (
            O => \N__8570\,
            I => \N__8557\
        );

    \I__1775\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8557\
        );

    \I__1774\ : Span4Mux_h
    port map (
            O => \N__8564\,
            I => \N__8552\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__8557\,
            I => \N__8552\
        );

    \I__1772\ : Span4Mux_h
    port map (
            O => \N__8552\,
            I => \N__8545\
        );

    \I__1771\ : InMux
    port map (
            O => \N__8551\,
            I => \N__8542\
        );

    \I__1770\ : InMux
    port map (
            O => \N__8550\,
            I => \N__8539\
        );

    \I__1769\ : InMux
    port map (
            O => \N__8549\,
            I => \N__8536\
        );

    \I__1768\ : InMux
    port map (
            O => \N__8548\,
            I => \N__8533\
        );

    \I__1767\ : Odrv4
    port map (
            O => \N__8545\,
            I => \U712_CHIP_RAM.N_297\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__8542\,
            I => \U712_CHIP_RAM.N_297\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__8539\,
            I => \U712_CHIP_RAM.N_297\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8536\,
            I => \U712_CHIP_RAM.N_297\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__8533\,
            I => \U712_CHIP_RAM.N_297\
        );

    \I__1762\ : CascadeMux
    port map (
            O => \N__8522\,
            I => \N__8516\
        );

    \I__1761\ : CascadeMux
    port map (
            O => \N__8521\,
            I => \N__8513\
        );

    \I__1760\ : CascadeMux
    port map (
            O => \N__8520\,
            I => \N__8508\
        );

    \I__1759\ : CascadeMux
    port map (
            O => \N__8519\,
            I => \N__8505\
        );

    \I__1758\ : InMux
    port map (
            O => \N__8516\,
            I => \N__8501\
        );

    \I__1757\ : InMux
    port map (
            O => \N__8513\,
            I => \N__8498\
        );

    \I__1756\ : InMux
    port map (
            O => \N__8512\,
            I => \N__8493\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8511\,
            I => \N__8493\
        );

    \I__1754\ : InMux
    port map (
            O => \N__8508\,
            I => \N__8490\
        );

    \I__1753\ : InMux
    port map (
            O => \N__8505\,
            I => \N__8485\
        );

    \I__1752\ : InMux
    port map (
            O => \N__8504\,
            I => \N__8485\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__8501\,
            I => \N__8480\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__8498\,
            I => \N__8480\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__8493\,
            I => \N__8473\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__8490\,
            I => \N__8473\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__8485\,
            I => \N__8473\
        );

    \I__1746\ : Span4Mux_h
    port map (
            O => \N__8480\,
            I => \N__8470\
        );

    \I__1745\ : Odrv4
    port map (
            O => \N__8473\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__1744\ : Odrv4
    port map (
            O => \N__8470\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__1743\ : InMux
    port map (
            O => \N__8465\,
            I => \N__8462\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__8462\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__1741\ : IoInMux
    port map (
            O => \N__8459\,
            I => \N__8456\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__8456\,
            I => \N__8453\
        );

    \I__1739\ : IoSpan4Mux
    port map (
            O => \N__8453\,
            I => \N__8450\
        );

    \I__1738\ : Span4Mux_s1_h
    port map (
            O => \N__8450\,
            I => \N__8447\
        );

    \I__1737\ : Sp12to4
    port map (
            O => \N__8447\,
            I => \N__8444\
        );

    \I__1736\ : Span12Mux_h
    port map (
            O => \N__8444\,
            I => \N__8441\
        );

    \I__1735\ : Odrv12
    port map (
            O => \N__8441\,
            I => \CMA_c_6\
        );

    \I__1734\ : InMux
    port map (
            O => \N__8438\,
            I => \N__8435\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__8435\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__1732\ : InMux
    port map (
            O => \N__8432\,
            I => \N__8429\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__8429\,
            I => \N__8426\
        );

    \I__1730\ : Odrv4
    port map (
            O => \N__8426\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__1729\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8420\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__8420\,
            I => \N__8417\
        );

    \I__1727\ : Span4Mux_v
    port map (
            O => \N__8417\,
            I => \N__8414\
        );

    \I__1726\ : Odrv4
    port map (
            O => \N__8414\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1725\ : InMux
    port map (
            O => \N__8411\,
            I => \N__8408\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__8408\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__1723\ : InMux
    port map (
            O => \N__8405\,
            I => \N__8402\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__8402\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8399\,
            I => \N__8396\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__8396\,
            I => \U712_BYTE_ENABLE.N_451\
        );

    \I__1719\ : IoInMux
    port map (
            O => \N__8393\,
            I => \N__8390\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__8390\,
            I => \N__8387\
        );

    \I__1717\ : Span4Mux_s3_v
    port map (
            O => \N__8387\,
            I => \N__8384\
        );

    \I__1716\ : Span4Mux_h
    port map (
            O => \N__8384\,
            I => \N__8381\
        );

    \I__1715\ : Sp12to4
    port map (
            O => \N__8381\,
            I => \N__8378\
        );

    \I__1714\ : Span12Mux_s10_v
    port map (
            O => \N__8378\,
            I => \N__8375\
        );

    \I__1713\ : Odrv12
    port map (
            O => \N__8375\,
            I => \N_211_i\
        );

    \I__1712\ : CascadeMux
    port map (
            O => \N__8372\,
            I => \U712_BYTE_ENABLE.N_410_cascade_\
        );

    \I__1711\ : IoInMux
    port map (
            O => \N__8369\,
            I => \N__8366\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__8366\,
            I => \N__8363\
        );

    \I__1709\ : Span12Mux_s4_h
    port map (
            O => \N__8363\,
            I => \N__8360\
        );

    \I__1708\ : Span12Mux_h
    port map (
            O => \N__8360\,
            I => \N__8357\
        );

    \I__1707\ : Span12Mux_v
    port map (
            O => \N__8357\,
            I => \N__8354\
        );

    \I__1706\ : Odrv12
    port map (
            O => \N__8354\,
            I => \N_148_i\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8351\,
            I => \N__8345\
        );

    \I__1704\ : InMux
    port map (
            O => \N__8350\,
            I => \N__8345\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__8345\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_a2Z0Z_0\
        );

    \I__1702\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8339\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__8339\,
            I => \N__8333\
        );

    \I__1700\ : InMux
    port map (
            O => \N__8338\,
            I => \N__8330\
        );

    \I__1699\ : InMux
    port map (
            O => \N__8337\,
            I => \N__8326\
        );

    \I__1698\ : InMux
    port map (
            O => \N__8336\,
            I => \N__8323\
        );

    \I__1697\ : Span4Mux_h
    port map (
            O => \N__8333\,
            I => \N__8320\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__8330\,
            I => \N__8317\
        );

    \I__1695\ : InMux
    port map (
            O => \N__8329\,
            I => \N__8314\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__8326\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__8323\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1692\ : Odrv4
    port map (
            O => \N__8320\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1691\ : Odrv4
    port map (
            O => \N__8317\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__8314\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1689\ : InMux
    port map (
            O => \N__8303\,
            I => \N__8300\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__8300\,
            I => \N__8291\
        );

    \I__1687\ : InMux
    port map (
            O => \N__8299\,
            I => \N__8288\
        );

    \I__1686\ : CascadeMux
    port map (
            O => \N__8298\,
            I => \N__8285\
        );

    \I__1685\ : CascadeMux
    port map (
            O => \N__8297\,
            I => \N__8281\
        );

    \I__1684\ : CascadeMux
    port map (
            O => \N__8296\,
            I => \N__8277\
        );

    \I__1683\ : InMux
    port map (
            O => \N__8295\,
            I => \N__8270\
        );

    \I__1682\ : InMux
    port map (
            O => \N__8294\,
            I => \N__8270\
        );

    \I__1681\ : Span4Mux_h
    port map (
            O => \N__8291\,
            I => \N__8267\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__8288\,
            I => \N__8264\
        );

    \I__1679\ : InMux
    port map (
            O => \N__8285\,
            I => \N__8261\
        );

    \I__1678\ : InMux
    port map (
            O => \N__8284\,
            I => \N__8258\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8281\,
            I => \N__8253\
        );

    \I__1676\ : InMux
    port map (
            O => \N__8280\,
            I => \N__8253\
        );

    \I__1675\ : InMux
    port map (
            O => \N__8277\,
            I => \N__8250\
        );

    \I__1674\ : InMux
    port map (
            O => \N__8276\,
            I => \N__8245\
        );

    \I__1673\ : InMux
    port map (
            O => \N__8275\,
            I => \N__8245\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__8270\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1671\ : Odrv4
    port map (
            O => \N__8267\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1670\ : Odrv4
    port map (
            O => \N__8264\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__8261\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__8258\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__8253\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__8250\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__8245\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1664\ : InMux
    port map (
            O => \N__8228\,
            I => \N__8222\
        );

    \I__1663\ : CascadeMux
    port map (
            O => \N__8227\,
            I => \N__8217\
        );

    \I__1662\ : CascadeMux
    port map (
            O => \N__8226\,
            I => \N__8214\
        );

    \I__1661\ : InMux
    port map (
            O => \N__8225\,
            I => \N__8210\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__8222\,
            I => \N__8207\
        );

    \I__1659\ : InMux
    port map (
            O => \N__8221\,
            I => \N__8202\
        );

    \I__1658\ : InMux
    port map (
            O => \N__8220\,
            I => \N__8202\
        );

    \I__1657\ : InMux
    port map (
            O => \N__8217\,
            I => \N__8197\
        );

    \I__1656\ : InMux
    port map (
            O => \N__8214\,
            I => \N__8197\
        );

    \I__1655\ : InMux
    port map (
            O => \N__8213\,
            I => \N__8194\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__8210\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__1653\ : Odrv4
    port map (
            O => \N__8207\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__8202\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__8197\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__8194\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__1649\ : CascadeMux
    port map (
            O => \N__8183\,
            I => \U712_REG_SM.N_95_cascade_\
        );

    \I__1648\ : InMux
    port map (
            O => \N__8180\,
            I => \N__8177\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__8177\,
            I => \U712_REG_SM.N_432\
        );

    \I__1646\ : IoInMux
    port map (
            O => \N__8174\,
            I => \N__8171\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__8171\,
            I => \N__8168\
        );

    \I__1644\ : Span12Mux_s0_v
    port map (
            O => \N__8168\,
            I => \N__8165\
        );

    \I__1643\ : Span12Mux_h
    port map (
            O => \N__8165\,
            I => \N__8161\
        );

    \I__1642\ : InMux
    port map (
            O => \N__8164\,
            I => \N__8158\
        );

    \I__1641\ : Odrv12
    port map (
            O => \N__8161\,
            I => \LDSn_c\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__8158\,
            I => \LDSn_c\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__8153\,
            I => \N__8146\
        );

    \I__1638\ : CascadeMux
    port map (
            O => \N__8152\,
            I => \N__8143\
        );

    \I__1637\ : CascadeMux
    port map (
            O => \N__8151\,
            I => \N__8140\
        );

    \I__1636\ : InMux
    port map (
            O => \N__8150\,
            I => \N__8134\
        );

    \I__1635\ : InMux
    port map (
            O => \N__8149\,
            I => \N__8134\
        );

    \I__1634\ : InMux
    port map (
            O => \N__8146\,
            I => \N__8131\
        );

    \I__1633\ : InMux
    port map (
            O => \N__8143\,
            I => \N__8126\
        );

    \I__1632\ : InMux
    port map (
            O => \N__8140\,
            I => \N__8126\
        );

    \I__1631\ : InMux
    port map (
            O => \N__8139\,
            I => \N__8121\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__8134\,
            I => \N__8106\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__8131\,
            I => \N__8106\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__8126\,
            I => \N__8106\
        );

    \I__1627\ : InMux
    port map (
            O => \N__8125\,
            I => \N__8101\
        );

    \I__1626\ : InMux
    port map (
            O => \N__8124\,
            I => \N__8101\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__8121\,
            I => \N__8098\
        );

    \I__1624\ : InMux
    port map (
            O => \N__8120\,
            I => \N__8095\
        );

    \I__1623\ : InMux
    port map (
            O => \N__8119\,
            I => \N__8092\
        );

    \I__1622\ : InMux
    port map (
            O => \N__8118\,
            I => \N__8089\
        );

    \I__1621\ : InMux
    port map (
            O => \N__8117\,
            I => \N__8082\
        );

    \I__1620\ : InMux
    port map (
            O => \N__8116\,
            I => \N__8082\
        );

    \I__1619\ : InMux
    port map (
            O => \N__8115\,
            I => \N__8082\
        );

    \I__1618\ : InMux
    port map (
            O => \N__8114\,
            I => \N__8077\
        );

    \I__1617\ : InMux
    port map (
            O => \N__8113\,
            I => \N__8077\
        );

    \I__1616\ : Span4Mux_v
    port map (
            O => \N__8106\,
            I => \N__8074\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__8101\,
            I => \N__8071\
        );

    \I__1614\ : Odrv12
    port map (
            O => \N__8098\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__8095\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__8092\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__8089\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__8082\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__8077\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1608\ : Odrv4
    port map (
            O => \N__8074\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1607\ : Odrv4
    port map (
            O => \N__8071\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1606\ : InMux
    port map (
            O => \N__8054\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__1605\ : CascadeMux
    port map (
            O => \N__8051\,
            I => \N__8047\
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__8050\,
            I => \N__8044\
        );

    \I__1603\ : InMux
    port map (
            O => \N__8047\,
            I => \N__8035\
        );

    \I__1602\ : InMux
    port map (
            O => \N__8044\,
            I => \N__8031\
        );

    \I__1601\ : InMux
    port map (
            O => \N__8043\,
            I => \N__8026\
        );

    \I__1600\ : InMux
    port map (
            O => \N__8042\,
            I => \N__8026\
        );

    \I__1599\ : InMux
    port map (
            O => \N__8041\,
            I => \N__8023\
        );

    \I__1598\ : InMux
    port map (
            O => \N__8040\,
            I => \N__8017\
        );

    \I__1597\ : InMux
    port map (
            O => \N__8039\,
            I => \N__8011\
        );

    \I__1596\ : InMux
    port map (
            O => \N__8038\,
            I => \N__8011\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__8035\,
            I => \N__8008\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__8034\,
            I => \N__8001\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__8031\,
            I => \N__7997\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__8026\,
            I => \N__7992\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__8023\,
            I => \N__7992\
        );

    \I__1590\ : InMux
    port map (
            O => \N__8022\,
            I => \N__7985\
        );

    \I__1589\ : InMux
    port map (
            O => \N__8021\,
            I => \N__7985\
        );

    \I__1588\ : InMux
    port map (
            O => \N__8020\,
            I => \N__7985\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__8017\,
            I => \N__7977\
        );

    \I__1586\ : InMux
    port map (
            O => \N__8016\,
            I => \N__7974\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__8011\,
            I => \N__7969\
        );

    \I__1584\ : Span4Mux_v
    port map (
            O => \N__8008\,
            I => \N__7969\
        );

    \I__1583\ : InMux
    port map (
            O => \N__8007\,
            I => \N__7960\
        );

    \I__1582\ : InMux
    port map (
            O => \N__8006\,
            I => \N__7960\
        );

    \I__1581\ : InMux
    port map (
            O => \N__8005\,
            I => \N__7960\
        );

    \I__1580\ : InMux
    port map (
            O => \N__8004\,
            I => \N__7960\
        );

    \I__1579\ : InMux
    port map (
            O => \N__8001\,
            I => \N__7955\
        );

    \I__1578\ : InMux
    port map (
            O => \N__8000\,
            I => \N__7955\
        );

    \I__1577\ : Span4Mux_h
    port map (
            O => \N__7997\,
            I => \N__7948\
        );

    \I__1576\ : Span4Mux_v
    port map (
            O => \N__7992\,
            I => \N__7948\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__7985\,
            I => \N__7948\
        );

    \I__1574\ : InMux
    port map (
            O => \N__7984\,
            I => \N__7941\
        );

    \I__1573\ : InMux
    port map (
            O => \N__7983\,
            I => \N__7941\
        );

    \I__1572\ : InMux
    port map (
            O => \N__7982\,
            I => \N__7941\
        );

    \I__1571\ : InMux
    port map (
            O => \N__7981\,
            I => \N__7936\
        );

    \I__1570\ : InMux
    port map (
            O => \N__7980\,
            I => \N__7936\
        );

    \I__1569\ : Odrv4
    port map (
            O => \N__7977\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__7974\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1567\ : Odrv4
    port map (
            O => \N__7969\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__7960\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__7955\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1564\ : Odrv4
    port map (
            O => \N__7948\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__7941\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__7936\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1561\ : CascadeMux
    port map (
            O => \N__7919\,
            I => \N__7916\
        );

    \I__1560\ : InMux
    port map (
            O => \N__7916\,
            I => \N__7913\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__7913\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__1558\ : InMux
    port map (
            O => \N__7910\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__7907\,
            I => \N__7902\
        );

    \I__1556\ : InMux
    port map (
            O => \N__7906\,
            I => \N__7898\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__7905\,
            I => \N__7894\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7902\,
            I => \N__7889\
        );

    \I__1553\ : InMux
    port map (
            O => \N__7901\,
            I => \N__7889\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__7898\,
            I => \N__7885\
        );

    \I__1551\ : InMux
    port map (
            O => \N__7897\,
            I => \N__7880\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7894\,
            I => \N__7880\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__7889\,
            I => \N__7877\
        );

    \I__1548\ : InMux
    port map (
            O => \N__7888\,
            I => \N__7869\
        );

    \I__1547\ : Span4Mux_h
    port map (
            O => \N__7885\,
            I => \N__7866\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__7880\,
            I => \N__7863\
        );

    \I__1545\ : Span4Mux_h
    port map (
            O => \N__7877\,
            I => \N__7860\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7853\
        );

    \I__1543\ : InMux
    port map (
            O => \N__7875\,
            I => \N__7853\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7874\,
            I => \N__7853\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7873\,
            I => \N__7848\
        );

    \I__1540\ : InMux
    port map (
            O => \N__7872\,
            I => \N__7848\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__7869\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1538\ : Odrv4
    port map (
            O => \N__7866\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1537\ : Odrv4
    port map (
            O => \N__7863\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1536\ : Odrv4
    port map (
            O => \N__7860\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__7853\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__7848\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1533\ : InMux
    port map (
            O => \N__7835\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__1532\ : InMux
    port map (
            O => \N__7832\,
            I => \N__7828\
        );

    \I__1531\ : InMux
    port map (
            O => \N__7831\,
            I => \N__7825\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__7828\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__7825\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7820\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__1527\ : InMux
    port map (
            O => \N__7817\,
            I => \N__7813\
        );

    \I__1526\ : InMux
    port map (
            O => \N__7816\,
            I => \N__7810\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__7813\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__7810\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1523\ : InMux
    port map (
            O => \N__7805\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__1522\ : InMux
    port map (
            O => \N__7802\,
            I => \N__7798\
        );

    \I__1521\ : InMux
    port map (
            O => \N__7801\,
            I => \N__7795\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__7798\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__7795\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1518\ : InMux
    port map (
            O => \N__7790\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__1517\ : InMux
    port map (
            O => \N__7787\,
            I => \N__7772\
        );

    \I__1516\ : InMux
    port map (
            O => \N__7786\,
            I => \N__7772\
        );

    \I__1515\ : InMux
    port map (
            O => \N__7785\,
            I => \N__7772\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7784\,
            I => \N__7772\
        );

    \I__1513\ : InMux
    port map (
            O => \N__7783\,
            I => \N__7769\
        );

    \I__1512\ : InMux
    port map (
            O => \N__7782\,
            I => \N__7764\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7781\,
            I => \N__7764\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__7772\,
            I => \U712_CHIP_RAM.N_200\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__7769\,
            I => \U712_CHIP_RAM.N_200\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7764\,
            I => \U712_CHIP_RAM.N_200\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7757\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__7754\,
            I => \N__7750\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7753\,
            I => \N__7747\
        );

    \I__1504\ : InMux
    port map (
            O => \N__7750\,
            I => \N__7744\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7747\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__7744\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1501\ : CEMux
    port map (
            O => \N__7739\,
            I => \N__7736\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__7736\,
            I => \N__7733\
        );

    \I__1499\ : Span4Mux_v
    port map (
            O => \N__7733\,
            I => \N__7729\
        );

    \I__1498\ : CEMux
    port map (
            O => \N__7732\,
            I => \N__7726\
        );

    \I__1497\ : Span4Mux_v
    port map (
            O => \N__7729\,
            I => \N__7721\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__7726\,
            I => \N__7721\
        );

    \I__1495\ : Span4Mux_h
    port map (
            O => \N__7721\,
            I => \N__7718\
        );

    \I__1494\ : Odrv4
    port map (
            O => \N__7718\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7715\,
            I => \N__7712\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__7712\,
            I => \N__7709\
        );

    \I__1491\ : Odrv12
    port map (
            O => \N__7709\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\
        );

    \I__1490\ : CascadeMux
    port map (
            O => \N__7706\,
            I => \U712_CHIP_RAM.N_294_cascade_\
        );

    \I__1489\ : CascadeMux
    port map (
            O => \N__7703\,
            I => \N__7700\
        );

    \I__1488\ : InMux
    port map (
            O => \N__7700\,
            I => \N__7696\
        );

    \I__1487\ : InMux
    port map (
            O => \N__7699\,
            I => \N__7693\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__7696\,
            I => \N__7687\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__7693\,
            I => \N__7687\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7692\,
            I => \N__7679\
        );

    \I__1483\ : Span4Mux_h
    port map (
            O => \N__7687\,
            I => \N__7672\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7686\,
            I => \N__7669\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7685\,
            I => \N__7664\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7684\,
            I => \N__7664\
        );

    \I__1479\ : InMux
    port map (
            O => \N__7683\,
            I => \N__7659\
        );

    \I__1478\ : InMux
    port map (
            O => \N__7682\,
            I => \N__7659\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__7679\,
            I => \N__7656\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7678\,
            I => \N__7651\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7677\,
            I => \N__7651\
        );

    \I__1474\ : InMux
    port map (
            O => \N__7676\,
            I => \N__7646\
        );

    \I__1473\ : InMux
    port map (
            O => \N__7675\,
            I => \N__7646\
        );

    \I__1472\ : Odrv4
    port map (
            O => \N__7672\,
            I => \U712_CHIP_RAM.N_288\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__7669\,
            I => \U712_CHIP_RAM.N_288\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__7664\,
            I => \U712_CHIP_RAM.N_288\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__7659\,
            I => \U712_CHIP_RAM.N_288\
        );

    \I__1468\ : Odrv4
    port map (
            O => \N__7656\,
            I => \U712_CHIP_RAM.N_288\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__7651\,
            I => \U712_CHIP_RAM.N_288\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7646\,
            I => \U712_CHIP_RAM.N_288\
        );

    \I__1465\ : CascadeMux
    port map (
            O => \N__7631\,
            I => \U712_CHIP_RAM.N_469_cascade_\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7628\,
            I => \N__7624\
        );

    \I__1463\ : InMux
    port map (
            O => \N__7627\,
            I => \N__7619\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__7624\,
            I => \N__7616\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7623\,
            I => \N__7613\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7622\,
            I => \N__7610\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__7619\,
            I => \U712_CHIP_RAM.N_557\
        );

    \I__1458\ : Odrv4
    port map (
            O => \N__7616\,
            I => \U712_CHIP_RAM.N_557\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__7613\,
            I => \U712_CHIP_RAM.N_557\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__7610\,
            I => \U712_CHIP_RAM.N_557\
        );

    \I__1455\ : InMux
    port map (
            O => \N__7601\,
            I => \N__7593\
        );

    \I__1454\ : InMux
    port map (
            O => \N__7600\,
            I => \N__7593\
        );

    \I__1453\ : InMux
    port map (
            O => \N__7599\,
            I => \N__7582\
        );

    \I__1452\ : InMux
    port map (
            O => \N__7598\,
            I => \N__7582\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__7593\,
            I => \N__7577\
        );

    \I__1450\ : CascadeMux
    port map (
            O => \N__7592\,
            I => \N__7571\
        );

    \I__1449\ : InMux
    port map (
            O => \N__7591\,
            I => \N__7564\
        );

    \I__1448\ : InMux
    port map (
            O => \N__7590\,
            I => \N__7564\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7589\,
            I => \N__7559\
        );

    \I__1446\ : InMux
    port map (
            O => \N__7588\,
            I => \N__7559\
        );

    \I__1445\ : InMux
    port map (
            O => \N__7587\,
            I => \N__7556\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__7582\,
            I => \N__7553\
        );

    \I__1443\ : InMux
    port map (
            O => \N__7581\,
            I => \N__7548\
        );

    \I__1442\ : InMux
    port map (
            O => \N__7580\,
            I => \N__7548\
        );

    \I__1441\ : Span4Mux_h
    port map (
            O => \N__7577\,
            I => \N__7545\
        );

    \I__1440\ : InMux
    port map (
            O => \N__7576\,
            I => \N__7538\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7575\,
            I => \N__7538\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7574\,
            I => \N__7538\
        );

    \I__1437\ : InMux
    port map (
            O => \N__7571\,
            I => \N__7531\
        );

    \I__1436\ : InMux
    port map (
            O => \N__7570\,
            I => \N__7531\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7569\,
            I => \N__7531\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__7564\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__7559\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__7556\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1431\ : Odrv4
    port map (
            O => \N__7553\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__7548\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1429\ : Odrv4
    port map (
            O => \N__7545\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__7538\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__7531\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1426\ : InMux
    port map (
            O => \N__7514\,
            I => \N__7511\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__7511\,
            I => \U712_CHIP_RAM.N_555\
        );

    \I__1424\ : CascadeMux
    port map (
            O => \N__7508\,
            I => \U712_CHIP_RAM.N_309_cascade_\
        );

    \I__1423\ : InMux
    port map (
            O => \N__7505\,
            I => \N__7502\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__7502\,
            I => \U712_CHIP_RAM.N_387\
        );

    \I__1421\ : CascadeMux
    port map (
            O => \N__7499\,
            I => \U712_CHIP_RAM.N_200_cascade_\
        );

    \I__1420\ : InMux
    port map (
            O => \N__7496\,
            I => \N__7493\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__7493\,
            I => \U712_CHIP_RAM.N_309\
        );

    \I__1418\ : InMux
    port map (
            O => \N__7490\,
            I => \N__7486\
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__7489\,
            I => \N__7482\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__7486\,
            I => \N__7479\
        );

    \I__1415\ : InMux
    port map (
            O => \N__7485\,
            I => \N__7474\
        );

    \I__1414\ : InMux
    port map (
            O => \N__7482\,
            I => \N__7474\
        );

    \I__1413\ : Odrv4
    port map (
            O => \N__7479\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__7474\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7469\,
            I => \N__7463\
        );

    \I__1410\ : InMux
    port map (
            O => \N__7468\,
            I => \N__7460\
        );

    \I__1409\ : InMux
    port map (
            O => \N__7467\,
            I => \N__7457\
        );

    \I__1408\ : InMux
    port map (
            O => \N__7466\,
            I => \N__7454\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__7463\,
            I => \N__7451\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__7460\,
            I => \N__7448\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__7457\,
            I => \N__7443\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__7454\,
            I => \N__7443\
        );

    \I__1403\ : Span4Mux_h
    port map (
            O => \N__7451\,
            I => \N__7439\
        );

    \I__1402\ : Span4Mux_h
    port map (
            O => \N__7448\,
            I => \N__7436\
        );

    \I__1401\ : Span4Mux_v
    port map (
            O => \N__7443\,
            I => \N__7433\
        );

    \I__1400\ : InMux
    port map (
            O => \N__7442\,
            I => \N__7430\
        );

    \I__1399\ : Odrv4
    port map (
            O => \N__7439\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1398\ : Odrv4
    port map (
            O => \N__7436\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1397\ : Odrv4
    port map (
            O => \N__7433\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__7430\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1395\ : InMux
    port map (
            O => \N__7421\,
            I => \N__7416\
        );

    \I__1394\ : InMux
    port map (
            O => \N__7420\,
            I => \N__7413\
        );

    \I__1393\ : InMux
    port map (
            O => \N__7419\,
            I => \N__7410\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__7416\,
            I => \N__7407\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__7413\,
            I => \N__7404\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__7410\,
            I => \N__7401\
        );

    \I__1389\ : Span4Mux_h
    port map (
            O => \N__7407\,
            I => \N__7398\
        );

    \I__1388\ : Span4Mux_h
    port map (
            O => \N__7404\,
            I => \N__7395\
        );

    \I__1387\ : Odrv4
    port map (
            O => \N__7401\,
            I => \U712_CHIP_RAM.N_285\
        );

    \I__1386\ : Odrv4
    port map (
            O => \N__7398\,
            I => \U712_CHIP_RAM.N_285\
        );

    \I__1385\ : Odrv4
    port map (
            O => \N__7395\,
            I => \U712_CHIP_RAM.N_285\
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__7388\,
            I => \U712_CHIP_RAM.N_285_cascade_\
        );

    \I__1383\ : InMux
    port map (
            O => \N__7385\,
            I => \N__7382\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__7382\,
            I => \N__7379\
        );

    \I__1381\ : Span4Mux_h
    port map (
            O => \N__7379\,
            I => \N__7371\
        );

    \I__1380\ : InMux
    port map (
            O => \N__7378\,
            I => \N__7366\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7377\,
            I => \N__7366\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7376\,
            I => \N__7363\
        );

    \I__1377\ : InMux
    port map (
            O => \N__7375\,
            I => \N__7358\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7374\,
            I => \N__7358\
        );

    \I__1375\ : Odrv4
    port map (
            O => \N__7371\,
            I => \U712_CHIP_RAM.N_293\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__7366\,
            I => \U712_CHIP_RAM.N_293\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__7363\,
            I => \U712_CHIP_RAM.N_293\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__7358\,
            I => \U712_CHIP_RAM.N_293\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__7349\,
            I => \N__7346\
        );

    \I__1370\ : InMux
    port map (
            O => \N__7346\,
            I => \N__7343\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__7343\,
            I => \N__7340\
        );

    \I__1368\ : Span4Mux_h
    port map (
            O => \N__7340\,
            I => \N__7337\
        );

    \I__1367\ : Odrv4
    port map (
            O => \N__7337\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_a2_0_2\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__7334\,
            I => \N__7330\
        );

    \I__1365\ : CascadeMux
    port map (
            O => \N__7333\,
            I => \N__7325\
        );

    \I__1364\ : InMux
    port map (
            O => \N__7330\,
            I => \N__7320\
        );

    \I__1363\ : InMux
    port map (
            O => \N__7329\,
            I => \N__7317\
        );

    \I__1362\ : InMux
    port map (
            O => \N__7328\,
            I => \N__7314\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7325\,
            I => \N__7309\
        );

    \I__1360\ : InMux
    port map (
            O => \N__7324\,
            I => \N__7309\
        );

    \I__1359\ : InMux
    port map (
            O => \N__7323\,
            I => \N__7304\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__7320\,
            I => \N__7299\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7317\,
            I => \N__7299\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__7314\,
            I => \N__7294\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__7309\,
            I => \N__7294\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__7308\,
            I => \N__7287\
        );

    \I__1353\ : InMux
    port map (
            O => \N__7307\,
            I => \N__7282\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__7304\,
            I => \N__7277\
        );

    \I__1351\ : Span4Mux_v
    port map (
            O => \N__7299\,
            I => \N__7277\
        );

    \I__1350\ : Span4Mux_v
    port map (
            O => \N__7294\,
            I => \N__7274\
        );

    \I__1349\ : InMux
    port map (
            O => \N__7293\,
            I => \N__7265\
        );

    \I__1348\ : InMux
    port map (
            O => \N__7292\,
            I => \N__7265\
        );

    \I__1347\ : InMux
    port map (
            O => \N__7291\,
            I => \N__7265\
        );

    \I__1346\ : InMux
    port map (
            O => \N__7290\,
            I => \N__7265\
        );

    \I__1345\ : InMux
    port map (
            O => \N__7287\,
            I => \N__7258\
        );

    \I__1344\ : InMux
    port map (
            O => \N__7286\,
            I => \N__7258\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7285\,
            I => \N__7258\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__7282\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1341\ : Odrv4
    port map (
            O => \N__7277\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1340\ : Odrv4
    port map (
            O => \N__7274\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__7265\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__7258\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1337\ : InMux
    port map (
            O => \N__7247\,
            I => \N__7244\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__7244\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__1335\ : InMux
    port map (
            O => \N__7241\,
            I => \bfn_12_9_0_\
        );

    \I__1334\ : InMux
    port map (
            O => \N__7238\,
            I => \N__7235\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__7235\,
            I => \N__7232\
        );

    \I__1332\ : Span4Mux_v
    port map (
            O => \N__7232\,
            I => \N__7229\
        );

    \I__1331\ : Span4Mux_h
    port map (
            O => \N__7229\,
            I => \N__7226\
        );

    \I__1330\ : Sp12to4
    port map (
            O => \N__7226\,
            I => \N__7223\
        );

    \I__1329\ : Span12Mux_h
    port map (
            O => \N__7223\,
            I => \N__7220\
        );

    \I__1328\ : Span12Mux_v
    port map (
            O => \N__7220\,
            I => \N__7217\
        );

    \I__1327\ : Odrv12
    port map (
            O => \N__7217\,
            I => \A_c_3\
        );

    \I__1326\ : InMux
    port map (
            O => \N__7214\,
            I => \N__7211\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__7211\,
            I => \N__7208\
        );

    \I__1324\ : Span4Mux_h
    port map (
            O => \N__7208\,
            I => \N__7205\
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__7205\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\
        );

    \I__1322\ : InMux
    port map (
            O => \N__7202\,
            I => \N__7199\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__7199\,
            I => \N__7196\
        );

    \I__1320\ : Span4Mux_h
    port map (
            O => \N__7196\,
            I => \N__7193\
        );

    \I__1319\ : Sp12to4
    port map (
            O => \N__7193\,
            I => \N__7190\
        );

    \I__1318\ : Span12Mux_v
    port map (
            O => \N__7190\,
            I => \N__7187\
        );

    \I__1317\ : Span12Mux_h
    port map (
            O => \N__7187\,
            I => \N__7184\
        );

    \I__1316\ : Odrv12
    port map (
            O => \N__7184\,
            I => \A_c_4\
        );

    \I__1315\ : InMux
    port map (
            O => \N__7181\,
            I => \N__7178\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__7178\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\
        );

    \I__1313\ : InMux
    port map (
            O => \N__7175\,
            I => \N__7172\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__7172\,
            I => \N__7169\
        );

    \I__1311\ : Span4Mux_v
    port map (
            O => \N__7169\,
            I => \N__7166\
        );

    \I__1310\ : Span4Mux_v
    port map (
            O => \N__7166\,
            I => \N__7163\
        );

    \I__1309\ : Sp12to4
    port map (
            O => \N__7163\,
            I => \N__7160\
        );

    \I__1308\ : Span12Mux_h
    port map (
            O => \N__7160\,
            I => \N__7157\
        );

    \I__1307\ : Odrv12
    port map (
            O => \N__7157\,
            I => \A_c_7\
        );

    \I__1306\ : InMux
    port map (
            O => \N__7154\,
            I => \N__7151\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__7151\,
            I => \N__7148\
        );

    \I__1304\ : Odrv4
    port map (
            O => \N__7148\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\
        );

    \I__1303\ : InMux
    port map (
            O => \N__7145\,
            I => \N__7142\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__7142\,
            I => \N__7139\
        );

    \I__1301\ : Span4Mux_v
    port map (
            O => \N__7139\,
            I => \N__7136\
        );

    \I__1300\ : Span4Mux_v
    port map (
            O => \N__7136\,
            I => \N__7133\
        );

    \I__1299\ : Sp12to4
    port map (
            O => \N__7133\,
            I => \N__7130\
        );

    \I__1298\ : Span12Mux_h
    port map (
            O => \N__7130\,
            I => \N__7127\
        );

    \I__1297\ : Odrv12
    port map (
            O => \N__7127\,
            I => \A_c_8\
        );

    \I__1296\ : InMux
    port map (
            O => \N__7124\,
            I => \N__7121\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__7121\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\
        );

    \I__1294\ : InMux
    port map (
            O => \N__7118\,
            I => \N__7115\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__7115\,
            I => \N__7112\
        );

    \I__1292\ : Span4Mux_v
    port map (
            O => \N__7112\,
            I => \N__7109\
        );

    \I__1291\ : Span4Mux_v
    port map (
            O => \N__7109\,
            I => \N__7106\
        );

    \I__1290\ : Sp12to4
    port map (
            O => \N__7106\,
            I => \N__7103\
        );

    \I__1289\ : Span12Mux_h
    port map (
            O => \N__7103\,
            I => \N__7100\
        );

    \I__1288\ : Odrv12
    port map (
            O => \N__7100\,
            I => \A_c_18\
        );

    \I__1287\ : InMux
    port map (
            O => \N__7097\,
            I => \N__7094\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__7094\,
            I => \N__7091\
        );

    \I__1285\ : Span4Mux_h
    port map (
            O => \N__7091\,
            I => \N__7088\
        );

    \I__1284\ : Odrv4
    port map (
            O => \N__7088\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\
        );

    \I__1283\ : InMux
    port map (
            O => \N__7085\,
            I => \N__7082\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__7082\,
            I => \N__7079\
        );

    \I__1281\ : Span12Mux_v
    port map (
            O => \N__7079\,
            I => \N__7076\
        );

    \I__1280\ : Span12Mux_h
    port map (
            O => \N__7076\,
            I => \N__7073\
        );

    \I__1279\ : Odrv12
    port map (
            O => \N__7073\,
            I => \A_c_5\
        );

    \I__1278\ : InMux
    port map (
            O => \N__7070\,
            I => \N__7067\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__7067\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\
        );

    \I__1276\ : CEMux
    port map (
            O => \N__7064\,
            I => \N__7061\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__7061\,
            I => \N__7057\
        );

    \I__1274\ : CEMux
    port map (
            O => \N__7060\,
            I => \N__7054\
        );

    \I__1273\ : Span4Mux_v
    port map (
            O => \N__7057\,
            I => \N__7051\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__7054\,
            I => \N__7048\
        );

    \I__1271\ : Span4Mux_h
    port map (
            O => \N__7051\,
            I => \N__7045\
        );

    \I__1270\ : Odrv4
    port map (
            O => \N__7048\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0\
        );

    \I__1269\ : Odrv4
    port map (
            O => \N__7045\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0\
        );

    \I__1268\ : InMux
    port map (
            O => \N__7040\,
            I => \N__7037\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__7037\,
            I => \N__7033\
        );

    \I__1266\ : InMux
    port map (
            O => \N__7036\,
            I => \N__7029\
        );

    \I__1265\ : Span4Mux_v
    port map (
            O => \N__7033\,
            I => \N__7026\
        );

    \I__1264\ : InMux
    port map (
            O => \N__7032\,
            I => \N__7023\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__7029\,
            I => \N__7020\
        );

    \I__1262\ : Sp12to4
    port map (
            O => \N__7026\,
            I => \N__7015\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__7023\,
            I => \N__7015\
        );

    \I__1260\ : Span12Mux_h
    port map (
            O => \N__7020\,
            I => \N__7012\
        );

    \I__1259\ : Span12Mux_h
    port map (
            O => \N__7015\,
            I => \N__7009\
        );

    \I__1258\ : Span12Mux_v
    port map (
            O => \N__7012\,
            I => \N__7006\
        );

    \I__1257\ : Span12Mux_v
    port map (
            O => \N__7009\,
            I => \N__7003\
        );

    \I__1256\ : Odrv12
    port map (
            O => \N__7006\,
            I => \AWEn_c\
        );

    \I__1255\ : Odrv12
    port map (
            O => \N__7003\,
            I => \AWEn_c\
        );

    \I__1254\ : InMux
    port map (
            O => \N__6998\,
            I => \N__6993\
        );

    \I__1253\ : InMux
    port map (
            O => \N__6997\,
            I => \N__6990\
        );

    \I__1252\ : InMux
    port map (
            O => \N__6996\,
            I => \N__6987\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__6993\,
            I => \N__6981\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__6990\,
            I => \N__6978\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__6987\,
            I => \N__6975\
        );

    \I__1248\ : InMux
    port map (
            O => \N__6986\,
            I => \N__6972\
        );

    \I__1247\ : InMux
    port map (
            O => \N__6985\,
            I => \N__6969\
        );

    \I__1246\ : InMux
    port map (
            O => \N__6984\,
            I => \N__6963\
        );

    \I__1245\ : Span4Mux_h
    port map (
            O => \N__6981\,
            I => \N__6960\
        );

    \I__1244\ : Span4Mux_v
    port map (
            O => \N__6978\,
            I => \N__6953\
        );

    \I__1243\ : Span4Mux_v
    port map (
            O => \N__6975\,
            I => \N__6953\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__6972\,
            I => \N__6953\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__6969\,
            I => \N__6950\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6968\,
            I => \N__6945\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6967\,
            I => \N__6945\
        );

    \I__1238\ : InMux
    port map (
            O => \N__6966\,
            I => \N__6942\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__6963\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1236\ : Odrv4
    port map (
            O => \N__6960\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1235\ : Odrv4
    port map (
            O => \N__6953\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1234\ : Odrv4
    port map (
            O => \N__6950\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__6945\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__6942\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1231\ : CEMux
    port map (
            O => \N__6929\,
            I => \N__6926\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__6926\,
            I => \N__6923\
        );

    \I__1229\ : Span4Mux_h
    port map (
            O => \N__6923\,
            I => \N__6920\
        );

    \I__1228\ : Odrv4
    port map (
            O => \N__6920\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0\
        );

    \I__1227\ : IoInMux
    port map (
            O => \N__6917\,
            I => \N__6914\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__6914\,
            I => \N__6911\
        );

    \I__1225\ : Span4Mux_s3_v
    port map (
            O => \N__6911\,
            I => \N__6908\
        );

    \I__1224\ : Span4Mux_h
    port map (
            O => \N__6908\,
            I => \N__6905\
        );

    \I__1223\ : Odrv4
    port map (
            O => \N__6905\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1222\ : InMux
    port map (
            O => \N__6902\,
            I => \N__6898\
        );

    \I__1221\ : CascadeMux
    port map (
            O => \N__6901\,
            I => \N__6894\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6898\,
            I => \N__6891\
        );

    \I__1219\ : CascadeMux
    port map (
            O => \N__6897\,
            I => \N__6886\
        );

    \I__1218\ : InMux
    port map (
            O => \N__6894\,
            I => \N__6883\
        );

    \I__1217\ : Span4Mux_h
    port map (
            O => \N__6891\,
            I => \N__6880\
        );

    \I__1216\ : InMux
    port map (
            O => \N__6890\,
            I => \N__6877\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6889\,
            I => \N__6874\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6886\,
            I => \N__6871\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__6883\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1212\ : Odrv4
    port map (
            O => \N__6880\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__6877\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__6874\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__6871\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1208\ : IoInMux
    port map (
            O => \N__6860\,
            I => \N__6857\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__6857\,
            I => \N__6854\
        );

    \I__1206\ : Span4Mux_s2_h
    port map (
            O => \N__6854\,
            I => \N__6851\
        );

    \I__1205\ : Span4Mux_v
    port map (
            O => \N__6851\,
            I => \N__6848\
        );

    \I__1204\ : Sp12to4
    port map (
            O => \N__6848\,
            I => \N__6845\
        );

    \I__1203\ : Span12Mux_h
    port map (
            O => \N__6845\,
            I => \N__6842\
        );

    \I__1202\ : Odrv12
    port map (
            O => \N__6842\,
            I => \WEn_c\
        );

    \I__1201\ : CascadeMux
    port map (
            O => \N__6839\,
            I => \N__6836\
        );

    \I__1200\ : InMux
    port map (
            O => \N__6836\,
            I => \N__6833\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__6833\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\
        );

    \I__1198\ : InMux
    port map (
            O => \N__6830\,
            I => \N__6827\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6827\,
            I => \N__6824\
        );

    \I__1196\ : Span12Mux_h
    port map (
            O => \N__6824\,
            I => \N__6821\
        );

    \I__1195\ : Odrv12
    port map (
            O => \N__6821\,
            I => \A_c_13\
        );

    \I__1194\ : CascadeMux
    port map (
            O => \N__6818\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\
        );

    \I__1193\ : InMux
    port map (
            O => \N__6815\,
            I => \N__6812\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__6812\,
            I => \N__6809\
        );

    \I__1191\ : Span12Mux_v
    port map (
            O => \N__6809\,
            I => \N__6806\
        );

    \I__1190\ : Span12Mux_h
    port map (
            O => \N__6806\,
            I => \N__6803\
        );

    \I__1189\ : Odrv12
    port map (
            O => \N__6803\,
            I => \A_c_15\
        );

    \I__1188\ : CascadeMux
    port map (
            O => \N__6800\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6797\,
            I => \N__6794\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__6794\,
            I => \N__6791\
        );

    \I__1185\ : Span4Mux_v
    port map (
            O => \N__6791\,
            I => \N__6788\
        );

    \I__1184\ : Span4Mux_v
    port map (
            O => \N__6788\,
            I => \N__6785\
        );

    \I__1183\ : Sp12to4
    port map (
            O => \N__6785\,
            I => \N__6782\
        );

    \I__1182\ : Span12Mux_h
    port map (
            O => \N__6782\,
            I => \N__6779\
        );

    \I__1181\ : Odrv12
    port map (
            O => \N__6779\,
            I => \A_c_6\
        );

    \I__1180\ : InMux
    port map (
            O => \N__6776\,
            I => \N__6773\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__6773\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6770\,
            I => \N__6767\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__6767\,
            I => \N__6764\
        );

    \I__1176\ : Span12Mux_v
    port map (
            O => \N__6764\,
            I => \N__6761\
        );

    \I__1175\ : Span12Mux_h
    port map (
            O => \N__6761\,
            I => \N__6758\
        );

    \I__1174\ : Span12Mux_v
    port map (
            O => \N__6758\,
            I => \N__6755\
        );

    \I__1173\ : Odrv12
    port map (
            O => \N__6755\,
            I => \A_c_2\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6752\,
            I => \N__6749\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__6749\,
            I => \N__6746\
        );

    \I__1170\ : Odrv4
    port map (
            O => \N__6746\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\
        );

    \I__1169\ : InMux
    port map (
            O => \N__6743\,
            I => \N__6740\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__6740\,
            I => \U712_REG_SM.STATE_COUNTsr_0\
        );

    \I__1167\ : InMux
    port map (
            O => \N__6737\,
            I => \N__6734\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6734\,
            I => \N__6731\
        );

    \I__1165\ : Span4Mux_h
    port map (
            O => \N__6731\,
            I => \N__6725\
        );

    \I__1164\ : InMux
    port map (
            O => \N__6730\,
            I => \N__6722\
        );

    \I__1163\ : InMux
    port map (
            O => \N__6729\,
            I => \N__6719\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6728\,
            I => \N__6716\
        );

    \I__1161\ : Odrv4
    port map (
            O => \N__6725\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__6722\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__6719\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__6716\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1157\ : InMux
    port map (
            O => \N__6707\,
            I => \N__6704\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__6704\,
            I => \U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6701\,
            I => \N__6698\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__6698\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_7\
        );

    \I__1153\ : InMux
    port map (
            O => \N__6695\,
            I => \N__6690\
        );

    \I__1152\ : InMux
    port map (
            O => \N__6694\,
            I => \N__6685\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6693\,
            I => \N__6685\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__6690\,
            I => \U712_REG_SM.N_307\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__6685\,
            I => \U712_REG_SM.N_307\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6680\,
            I => \N__6676\
        );

    \I__1147\ : InMux
    port map (
            O => \N__6679\,
            I => \N__6673\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__6676\,
            I => \U712_REG_SM.N_553\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__6673\,
            I => \U712_REG_SM.N_553\
        );

    \I__1144\ : InMux
    port map (
            O => \N__6668\,
            I => \N__6665\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__6665\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_4\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6662\,
            I => \N__6656\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6661\,
            I => \N__6656\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__6656\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_5\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6653\,
            I => \N__6650\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__6650\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_6\
        );

    \I__1137\ : IoInMux
    port map (
            O => \N__6647\,
            I => \N__6644\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6644\,
            I => \N__6641\
        );

    \I__1135\ : IoSpan4Mux
    port map (
            O => \N__6641\,
            I => \N__6638\
        );

    \I__1134\ : Span4Mux_s3_v
    port map (
            O => \N__6638\,
            I => \N__6635\
        );

    \I__1133\ : Span4Mux_v
    port map (
            O => \N__6635\,
            I => \N__6632\
        );

    \I__1132\ : Odrv4
    port map (
            O => \N__6632\,
            I => \N_130_i\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6629\,
            I => \N__6626\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__6626\,
            I => \N__6623\
        );

    \I__1129\ : Odrv4
    port map (
            O => \N__6623\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6620\,
            I => \N__6615\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6619\,
            I => \N__6612\
        );

    \I__1126\ : InMux
    port map (
            O => \N__6618\,
            I => \N__6609\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6615\,
            I => \N__6606\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__6612\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6609\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__1122\ : Odrv4
    port map (
            O => \N__6606\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__1121\ : CascadeMux
    port map (
            O => \N__6599\,
            I => \U712_REG_SM.N_306_cascade_\
        );

    \I__1120\ : CascadeMux
    port map (
            O => \N__6596\,
            I => \U712_REG_SM.N_399_cascade_\
        );

    \I__1119\ : InMux
    port map (
            O => \N__6593\,
            I => \N__6590\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6590\,
            I => \U712_REG_SM.REG_CYCLE_5_iv_0_0\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6587\,
            I => \N__6581\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6586\,
            I => \N__6581\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__6581\,
            I => \U712_REG_SM.N_311\
        );

    \I__1114\ : CascadeMux
    port map (
            O => \N__6578\,
            I => \U712_REG_SM.N_353_cascade_\
        );

    \I__1113\ : InMux
    port map (
            O => \N__6575\,
            I => \N__6570\
        );

    \I__1112\ : InMux
    port map (
            O => \N__6574\,
            I => \N__6565\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6573\,
            I => \N__6565\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6570\,
            I => \N__6562\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__6565\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1108\ : Odrv4
    port map (
            O => \N__6562\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6557\,
            I => \N__6554\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__6554\,
            I => \N__6551\
        );

    \I__1105\ : Odrv4
    port map (
            O => \N__6551\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1104\ : InMux
    port map (
            O => \N__6548\,
            I => \N__6545\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__6545\,
            I => \U712_REG_SM.N_322\
        );

    \I__1102\ : InMux
    port map (
            O => \N__6542\,
            I => \N__6535\
        );

    \I__1101\ : InMux
    port map (
            O => \N__6541\,
            I => \N__6535\
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__6540\,
            I => \N__6532\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__6535\,
            I => \N__6528\
        );

    \I__1098\ : InMux
    port map (
            O => \N__6532\,
            I => \N__6525\
        );

    \I__1097\ : InMux
    port map (
            O => \N__6531\,
            I => \N__6522\
        );

    \I__1096\ : Span4Mux_h
    port map (
            O => \N__6528\,
            I => \N__6519\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__6525\,
            I => \REG_TACK\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6522\,
            I => \REG_TACK\
        );

    \I__1093\ : Odrv4
    port map (
            O => \N__6519\,
            I => \REG_TACK\
        );

    \I__1092\ : CascadeMux
    port map (
            O => \N__6512\,
            I => \U712_CHIP_RAM.N_356_cascade_\
        );

    \I__1091\ : InMux
    port map (
            O => \N__6509\,
            I => \N__6506\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__6506\,
            I => \U712_CHIP_RAM.N_448\
        );

    \I__1089\ : CascadeMux
    port map (
            O => \N__6503\,
            I => \U712_CHIP_RAM.N_288_cascade_\
        );

    \I__1088\ : InMux
    port map (
            O => \N__6500\,
            I => \N__6496\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6499\,
            I => \N__6493\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__6496\,
            I => \U712_CHIP_RAM.N_473\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__6493\,
            I => \U712_CHIP_RAM.N_473\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__6488\,
            I => \U712_CHIP_RAM.N_473_cascade_\
        );

    \I__1083\ : InMux
    port map (
            O => \N__6485\,
            I => \N__6482\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__6482\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_i_1_0\
        );

    \I__1081\ : InMux
    port map (
            O => \N__6479\,
            I => \N__6476\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__6476\,
            I => \N__6471\
        );

    \I__1079\ : InMux
    port map (
            O => \N__6475\,
            I => \N__6466\
        );

    \I__1078\ : InMux
    port map (
            O => \N__6474\,
            I => \N__6466\
        );

    \I__1077\ : Odrv4
    port map (
            O => \N__6471\,
            I => \U712_CHIP_RAM.N_362\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__6466\,
            I => \U712_CHIP_RAM.N_362\
        );

    \I__1075\ : InMux
    port map (
            O => \N__6461\,
            I => \N__6458\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__6458\,
            I => \N__6451\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6457\,
            I => \N__6446\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6456\,
            I => \N__6446\
        );

    \I__1071\ : InMux
    port map (
            O => \N__6455\,
            I => \N__6443\
        );

    \I__1070\ : InMux
    port map (
            O => \N__6454\,
            I => \N__6440\
        );

    \I__1069\ : Odrv4
    port map (
            O => \N__6451\,
            I => \U712_CHIP_RAM.N_463\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__6446\,
            I => \U712_CHIP_RAM.N_463\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__6443\,
            I => \U712_CHIP_RAM.N_463\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__6440\,
            I => \U712_CHIP_RAM.N_463\
        );

    \I__1065\ : CEMux
    port map (
            O => \N__6431\,
            I => \N__6428\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__6428\,
            I => \N__6425\
        );

    \I__1063\ : Odrv4
    port map (
            O => \N__6425\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_0\
        );

    \I__1062\ : InMux
    port map (
            O => \N__6422\,
            I => \N__6418\
        );

    \I__1061\ : InMux
    port map (
            O => \N__6421\,
            I => \N__6415\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__6418\,
            I => \N__6410\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__6415\,
            I => \N__6410\
        );

    \I__1058\ : Odrv4
    port map (
            O => \N__6410\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__1057\ : IoInMux
    port map (
            O => \N__6407\,
            I => \N__6404\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__6404\,
            I => \N__6401\
        );

    \I__1055\ : IoSpan4Mux
    port map (
            O => \N__6401\,
            I => \N__6398\
        );

    \I__1054\ : Span4Mux_s2_v
    port map (
            O => \N__6398\,
            I => \N__6395\
        );

    \I__1053\ : Sp12to4
    port map (
            O => \N__6395\,
            I => \N__6392\
        );

    \I__1052\ : Span12Mux_v
    port map (
            O => \N__6392\,
            I => \N__6388\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6391\,
            I => \N__6385\
        );

    \I__1050\ : Odrv12
    port map (
            O => \N__6388\,
            I => \DBDIR_c\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__6385\,
            I => \DBDIR_c\
        );

    \I__1048\ : CascadeMux
    port map (
            O => \N__6380\,
            I => \N__6377\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6377\,
            I => \N__6374\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__6374\,
            I => \N__6371\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__6371\,
            I => \U712_CHIP_RAM.N_556\
        );

    \I__1044\ : InMux
    port map (
            O => \N__6368\,
            I => \N__6365\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__6365\,
            I => \N__6360\
        );

    \I__1042\ : InMux
    port map (
            O => \N__6364\,
            I => \N__6357\
        );

    \I__1041\ : InMux
    port map (
            O => \N__6363\,
            I => \N__6354\
        );

    \I__1040\ : Odrv4
    port map (
            O => \N__6360\,
            I => \U712_CHIP_RAM.N_302\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__6357\,
            I => \U712_CHIP_RAM.N_302\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__6354\,
            I => \U712_CHIP_RAM.N_302\
        );

    \I__1037\ : InMux
    port map (
            O => \N__6347\,
            I => \N__6344\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__6344\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER19\
        );

    \I__1035\ : CascadeMux
    port map (
            O => \N__6341\,
            I => \U712_CHIP_RAM.N_355_cascade_\
        );

    \I__1034\ : CascadeMux
    port map (
            O => \N__6338\,
            I => \N__6335\
        );

    \I__1033\ : InMux
    port map (
            O => \N__6335\,
            I => \N__6332\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__6332\,
            I => \N__6329\
        );

    \I__1031\ : Odrv4
    port map (
            O => \N__6329\,
            I => \U712_CHIP_RAM.N_389\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6326\,
            I => \N__6320\
        );

    \I__1029\ : InMux
    port map (
            O => \N__6325\,
            I => \N__6320\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__6320\,
            I => \U712_CHIP_RAM.N_301\
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__6317\,
            I => \N__6313\
        );

    \I__1026\ : CascadeMux
    port map (
            O => \N__6316\,
            I => \N__6309\
        );

    \I__1025\ : InMux
    port map (
            O => \N__6313\,
            I => \N__6305\
        );

    \I__1024\ : CascadeMux
    port map (
            O => \N__6312\,
            I => \N__6302\
        );

    \I__1023\ : InMux
    port map (
            O => \N__6309\,
            I => \N__6298\
        );

    \I__1022\ : InMux
    port map (
            O => \N__6308\,
            I => \N__6295\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__6305\,
            I => \N__6292\
        );

    \I__1020\ : InMux
    port map (
            O => \N__6302\,
            I => \N__6287\
        );

    \I__1019\ : InMux
    port map (
            O => \N__6301\,
            I => \N__6287\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__6298\,
            I => \U712_CHIP_RAM.N_289\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__6295\,
            I => \U712_CHIP_RAM.N_289\
        );

    \I__1016\ : Odrv4
    port map (
            O => \N__6292\,
            I => \U712_CHIP_RAM.N_289\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__6287\,
            I => \U712_CHIP_RAM.N_289\
        );

    \I__1014\ : InMux
    port map (
            O => \N__6278\,
            I => \N__6275\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__6275\,
            I => \N__6272\
        );

    \I__1012\ : Odrv4
    port map (
            O => \N__6272\,
            I => \U712_CHIP_RAM.N_356\
        );

    \I__1011\ : CascadeMux
    port map (
            O => \N__6269\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6266\,
            I => \N__6263\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__6263\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__1008\ : InMux
    port map (
            O => \N__6260\,
            I => \N__6257\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__6257\,
            I => \N__6254\
        );

    \I__1006\ : Span4Mux_h
    port map (
            O => \N__6254\,
            I => \N__6250\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6253\,
            I => \N__6247\
        );

    \I__1004\ : Odrv4
    port map (
            O => \N__6250\,
            I => \U712_CHIP_RAM.N_551\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__6247\,
            I => \U712_CHIP_RAM.N_551\
        );

    \I__1002\ : CEMux
    port map (
            O => \N__6242\,
            I => \N__6239\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__6239\,
            I => \N__6236\
        );

    \I__1000\ : Span4Mux_v
    port map (
            O => \N__6236\,
            I => \N__6233\
        );

    \I__999\ : Odrv4
    port map (
            O => \N__6233\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_10_0_0\
        );

    \I__998\ : InMux
    port map (
            O => \N__6230\,
            I => \N__6226\
        );

    \I__997\ : InMux
    port map (
            O => \N__6229\,
            I => \N__6223\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__6226\,
            I => \N__6218\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__6223\,
            I => \N__6218\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__6218\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0\
        );

    \I__993\ : InMux
    port map (
            O => \N__6215\,
            I => \N__6212\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__6212\,
            I => \N__6209\
        );

    \I__991\ : Span4Mux_v
    port map (
            O => \N__6209\,
            I => \N__6206\
        );

    \I__990\ : Sp12to4
    port map (
            O => \N__6206\,
            I => \N__6203\
        );

    \I__989\ : Span12Mux_h
    port map (
            O => \N__6203\,
            I => \N__6200\
        );

    \I__988\ : Span12Mux_v
    port map (
            O => \N__6200\,
            I => \N__6197\
        );

    \I__987\ : Odrv12
    port map (
            O => \N__6197\,
            I => \A_c_20\
        );

    \I__986\ : InMux
    port map (
            O => \N__6194\,
            I => \N__6190\
        );

    \I__985\ : InMux
    port map (
            O => \N__6193\,
            I => \N__6187\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__6190\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__6187\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__982\ : CascadeMux
    port map (
            O => \N__6182\,
            I => \U712_CHIP_RAM.N_555_cascade_\
        );

    \I__981\ : InMux
    port map (
            O => \N__6179\,
            I => \N__6176\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__6176\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER16\
        );

    \I__979\ : InMux
    port map (
            O => \N__6173\,
            I => \N__6170\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__6170\,
            I => \N__6167\
        );

    \I__977\ : Odrv4
    port map (
            O => \N__6167\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__6164\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER16_cascade_\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__6161\,
            I => \U712_REG_SM.N_307_cascade_\
        );

    \I__974\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6153\
        );

    \I__973\ : InMux
    port map (
            O => \N__6157\,
            I => \N__6150\
        );

    \I__972\ : InMux
    port map (
            O => \N__6156\,
            I => \N__6147\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__6153\,
            I => \N__6142\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__6150\,
            I => \N__6142\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__6147\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_3\
        );

    \I__968\ : Odrv4
    port map (
            O => \N__6142\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_3\
        );

    \I__967\ : IoInMux
    port map (
            O => \N__6137\,
            I => \N__6134\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__6134\,
            I => \N__6131\
        );

    \I__965\ : Span4Mux_s2_v
    port map (
            O => \N__6131\,
            I => \N__6128\
        );

    \I__964\ : Sp12to4
    port map (
            O => \N__6128\,
            I => \N__6125\
        );

    \I__963\ : Span12Mux_h
    port map (
            O => \N__6125\,
            I => \N__6120\
        );

    \I__962\ : InMux
    port map (
            O => \N__6124\,
            I => \N__6117\
        );

    \I__961\ : InMux
    port map (
            O => \N__6123\,
            I => \N__6114\
        );

    \I__960\ : Odrv12
    port map (
            O => \N__6120\,
            I => \REGENn_c\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__6117\,
            I => \REGENn_c\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__6114\,
            I => \REGENn_c\
        );

    \I__957\ : InMux
    port map (
            O => \N__6107\,
            I => \N__6104\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__6104\,
            I => \U712_REG_SM.REGENn_e_1\
        );

    \I__955\ : InMux
    port map (
            O => \N__6101\,
            I => \N__6095\
        );

    \I__954\ : InMux
    port map (
            O => \N__6100\,
            I => \N__6095\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__6095\,
            I => \N__6090\
        );

    \I__952\ : InMux
    port map (
            O => \N__6094\,
            I => \N__6087\
        );

    \I__951\ : InMux
    port map (
            O => \N__6093\,
            I => \N__6084\
        );

    \I__950\ : Odrv4
    port map (
            O => \N__6090\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__6087\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__6084\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__947\ : InMux
    port map (
            O => \N__6077\,
            I => \N__6070\
        );

    \I__946\ : InMux
    port map (
            O => \N__6076\,
            I => \N__6070\
        );

    \I__945\ : InMux
    port map (
            O => \N__6075\,
            I => \N__6067\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__6070\,
            I => \N__6064\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__6067\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__942\ : Odrv4
    port map (
            O => \N__6064\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__941\ : InMux
    port map (
            O => \N__6059\,
            I => \N__6056\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__6056\,
            I => \N__6053\
        );

    \I__939\ : Span12Mux_h
    port map (
            O => \N__6053\,
            I => \N__6050\
        );

    \I__938\ : Odrv12
    port map (
            O => \N__6050\,
            I => \A_c_12\
        );

    \I__937\ : IoInMux
    port map (
            O => \N__6047\,
            I => \N__6044\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__6044\,
            I => \N__6041\
        );

    \I__935\ : IoSpan4Mux
    port map (
            O => \N__6041\,
            I => \N__6038\
        );

    \I__934\ : Span4Mux_s2_v
    port map (
            O => \N__6038\,
            I => \N__6034\
        );

    \I__933\ : InMux
    port map (
            O => \N__6037\,
            I => \N__6031\
        );

    \I__932\ : Sp12to4
    port map (
            O => \N__6034\,
            I => \N__6028\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__6031\,
            I => \N__6025\
        );

    \I__930\ : Span12Mux_s8_v
    port map (
            O => \N__6028\,
            I => \N__6022\
        );

    \I__929\ : Span4Mux_v
    port map (
            O => \N__6025\,
            I => \N__6019\
        );

    \I__928\ : Span12Mux_v
    port map (
            O => \N__6022\,
            I => \N__6016\
        );

    \I__927\ : Sp12to4
    port map (
            O => \N__6019\,
            I => \N__6013\
        );

    \I__926\ : Span12Mux_h
    port map (
            O => \N__6016\,
            I => \N__6010\
        );

    \I__925\ : Span12Mux_h
    port map (
            O => \N__6013\,
            I => \N__6007\
        );

    \I__924\ : Odrv12
    port map (
            O => \N__6010\,
            I => \A_c_11\
        );

    \I__923\ : Odrv12
    port map (
            O => \N__6007\,
            I => \A_c_11\
        );

    \I__922\ : InMux
    port map (
            O => \N__6002\,
            I => \N__5998\
        );

    \I__921\ : InMux
    port map (
            O => \N__6001\,
            I => \N__5995\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__5998\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__5995\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\
        );

    \I__918\ : CascadeMux
    port map (
            O => \N__5990\,
            I => \N__5987\
        );

    \I__917\ : InMux
    port map (
            O => \N__5987\,
            I => \N__5984\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__5984\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\
        );

    \I__915\ : InMux
    port map (
            O => \N__5981\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\
        );

    \I__914\ : InMux
    port map (
            O => \N__5978\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__5975\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3_cascade_\
        );

    \I__912\ : InMux
    port map (
            O => \N__5972\,
            I => \N__5968\
        );

    \I__911\ : InMux
    port map (
            O => \N__5971\,
            I => \N__5965\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__5968\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5965\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\
        );

    \I__908\ : InMux
    port map (
            O => \N__5960\,
            I => \N__5957\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__5957\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\
        );

    \I__906\ : InMux
    port map (
            O => \N__5954\,
            I => \N__5950\
        );

    \I__905\ : InMux
    port map (
            O => \N__5953\,
            I => \N__5947\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__5950\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ0Z_1\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5947\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ0Z_1\
        );

    \I__902\ : InMux
    port map (
            O => \N__5942\,
            I => \N__5931\
        );

    \I__901\ : InMux
    port map (
            O => \N__5941\,
            I => \N__5931\
        );

    \I__900\ : InMux
    port map (
            O => \N__5940\,
            I => \N__5924\
        );

    \I__899\ : InMux
    port map (
            O => \N__5939\,
            I => \N__5924\
        );

    \I__898\ : InMux
    port map (
            O => \N__5938\,
            I => \N__5924\
        );

    \I__897\ : InMux
    port map (
            O => \N__5937\,
            I => \N__5919\
        );

    \I__896\ : InMux
    port map (
            O => \N__5936\,
            I => \N__5919\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__5931\,
            I => \N__5916\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__5924\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__5919\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__892\ : Odrv4
    port map (
            O => \N__5916\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__5909\,
            I => \N__5906\
        );

    \I__890\ : InMux
    port map (
            O => \N__5906\,
            I => \N__5903\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__5903\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\
        );

    \I__888\ : CascadeMux
    port map (
            O => \N__5900\,
            I => \N__5897\
        );

    \I__887\ : InMux
    port map (
            O => \N__5897\,
            I => \N__5893\
        );

    \I__886\ : InMux
    port map (
            O => \N__5896\,
            I => \N__5890\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5893\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__5890\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\
        );

    \I__883\ : CascadeMux
    port map (
            O => \N__5885\,
            I => \N__5882\
        );

    \I__882\ : InMux
    port map (
            O => \N__5882\,
            I => \N__5875\
        );

    \I__881\ : InMux
    port map (
            O => \N__5881\,
            I => \N__5875\
        );

    \I__880\ : InMux
    port map (
            O => \N__5880\,
            I => \N__5872\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__5875\,
            I => \N__5866\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__5872\,
            I => \N__5866\
        );

    \I__877\ : InMux
    port map (
            O => \N__5871\,
            I => \N__5863\
        );

    \I__876\ : Span4Mux_v
    port map (
            O => \N__5866\,
            I => \N__5860\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5863\,
            I => \CPU_TACKm\
        );

    \I__874\ : Odrv4
    port map (
            O => \N__5860\,
            I => \CPU_TACKm\
        );

    \I__873\ : InMux
    port map (
            O => \N__5855\,
            I => \N__5852\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__5852\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__871\ : CascadeMux
    port map (
            O => \N__5849\,
            I => \N__5842\
        );

    \I__870\ : CascadeMux
    port map (
            O => \N__5848\,
            I => \N__5838\
        );

    \I__869\ : InMux
    port map (
            O => \N__5847\,
            I => \N__5834\
        );

    \I__868\ : InMux
    port map (
            O => \N__5846\,
            I => \N__5827\
        );

    \I__867\ : InMux
    port map (
            O => \N__5845\,
            I => \N__5827\
        );

    \I__866\ : InMux
    port map (
            O => \N__5842\,
            I => \N__5827\
        );

    \I__865\ : InMux
    port map (
            O => \N__5841\,
            I => \N__5820\
        );

    \I__864\ : InMux
    port map (
            O => \N__5838\,
            I => \N__5820\
        );

    \I__863\ : InMux
    port map (
            O => \N__5837\,
            I => \N__5820\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__5834\,
            I => \N__5815\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__5827\,
            I => \N__5810\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__5820\,
            I => \N__5810\
        );

    \I__859\ : InMux
    port map (
            O => \N__5819\,
            I => \N__5805\
        );

    \I__858\ : InMux
    port map (
            O => \N__5818\,
            I => \N__5805\
        );

    \I__857\ : Odrv12
    port map (
            O => \N__5815\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__856\ : Odrv4
    port map (
            O => \N__5810\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__5805\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__854\ : CascadeMux
    port map (
            O => \N__5798\,
            I => \N__5794\
        );

    \I__853\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5791\
        );

    \I__852\ : InMux
    port map (
            O => \N__5794\,
            I => \N__5788\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__5791\,
            I => \DBR_SYNC_i_1\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__5788\,
            I => \DBR_SYNC_i_1\
        );

    \I__849\ : InMux
    port map (
            O => \N__5783\,
            I => \N__5780\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__5780\,
            I => \U712_CHIP_RAM.N_360\
        );

    \I__847\ : InMux
    port map (
            O => \N__5777\,
            I => \N__5773\
        );

    \I__846\ : InMux
    port map (
            O => \N__5776\,
            I => \N__5770\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__5773\,
            I => \U712_CHIP_RAM.N_418\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__5770\,
            I => \U712_CHIP_RAM.N_418\
        );

    \I__843\ : InMux
    port map (
            O => \N__5765\,
            I => \N__5762\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__5762\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_5_0\
        );

    \I__841\ : CascadeMux
    port map (
            O => \N__5759\,
            I => \U712_REG_SM.N_400_cascade_\
        );

    \I__840\ : CascadeMux
    port map (
            O => \N__5756\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3_cascade_\
        );

    \I__839\ : CascadeMux
    port map (
            O => \N__5753\,
            I => \N__5750\
        );

    \I__838\ : InMux
    port map (
            O => \N__5750\,
            I => \N__5747\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__5747\,
            I => \U712_CHIP_RAM.N_405\
        );

    \I__836\ : InMux
    port map (
            O => \N__5744\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\
        );

    \I__835\ : CascadeMux
    port map (
            O => \N__5741\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_cascade_\
        );

    \I__834\ : InMux
    port map (
            O => \N__5738\,
            I => \N__5735\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__5735\,
            I => \N__5732\
        );

    \I__832\ : Odrv4
    port map (
            O => \N__5732\,
            I => \U712_CHIP_RAM.N_439\
        );

    \I__831\ : InMux
    port map (
            O => \N__5729\,
            I => \N__5726\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__5726\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_0_a2_1_0\
        );

    \I__829\ : CascadeMux
    port map (
            O => \N__5723\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\
        );

    \I__828\ : CascadeMux
    port map (
            O => \N__5720\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_cascade_\
        );

    \I__827\ : IoInMux
    port map (
            O => \N__5717\,
            I => \N__5714\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__5714\,
            I => \N__5711\
        );

    \I__825\ : Span4Mux_s2_h
    port map (
            O => \N__5711\,
            I => \N__5708\
        );

    \I__824\ : Span4Mux_h
    port map (
            O => \N__5708\,
            I => \N__5705\
        );

    \I__823\ : Sp12to4
    port map (
            O => \N__5705\,
            I => \N__5702\
        );

    \I__822\ : Span12Mux_s11_v
    port map (
            O => \N__5702\,
            I => \N__5699\
        );

    \I__821\ : Span12Mux_h
    port map (
            O => \N__5699\,
            I => \N__5696\
        );

    \I__820\ : Odrv12
    port map (
            O => \N__5696\,
            I => \CLK_EN_c\
        );

    \I__819\ : CEMux
    port map (
            O => \N__5693\,
            I => \N__5690\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__5690\,
            I => \N__5687\
        );

    \I__817\ : Span4Mux_h
    port map (
            O => \N__5687\,
            I => \N__5684\
        );

    \I__816\ : Odrv4
    port map (
            O => \N__5684\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0\
        );

    \I__815\ : CascadeMux
    port map (
            O => \N__5681\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_10_0_cascade_\
        );

    \I__814\ : InMux
    port map (
            O => \N__5678\,
            I => \N__5675\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5675\,
            I => \N__5672\
        );

    \I__812\ : Span4Mux_v
    port map (
            O => \N__5672\,
            I => \N__5664\
        );

    \I__811\ : InMux
    port map (
            O => \N__5671\,
            I => \N__5661\
        );

    \I__810\ : InMux
    port map (
            O => \N__5670\,
            I => \N__5656\
        );

    \I__809\ : InMux
    port map (
            O => \N__5669\,
            I => \N__5656\
        );

    \I__808\ : InMux
    port map (
            O => \N__5668\,
            I => \N__5653\
        );

    \I__807\ : InMux
    port map (
            O => \N__5667\,
            I => \N__5650\
        );

    \I__806\ : Odrv4
    port map (
            O => \N__5664\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__5661\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__5656\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5653\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__5650\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__801\ : InMux
    port map (
            O => \N__5639\,
            I => \N__5633\
        );

    \I__800\ : InMux
    port map (
            O => \N__5638\,
            I => \N__5626\
        );

    \I__799\ : InMux
    port map (
            O => \N__5637\,
            I => \N__5626\
        );

    \I__798\ : InMux
    port map (
            O => \N__5636\,
            I => \N__5626\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5633\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__5626\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__5621\,
            I => \N__5618\
        );

    \I__794\ : InMux
    port map (
            O => \N__5618\,
            I => \N__5615\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__5615\,
            I => \U712_CHIP_RAM.N_445\
        );

    \I__792\ : CascadeMux
    port map (
            O => \N__5612\,
            I => \N__5609\
        );

    \I__791\ : InMux
    port map (
            O => \N__5609\,
            I => \N__5606\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__5606\,
            I => \U712_CHIP_RAM.N_208\
        );

    \I__789\ : InMux
    port map (
            O => \N__5603\,
            I => \N__5599\
        );

    \I__788\ : InMux
    port map (
            O => \N__5602\,
            I => \N__5596\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5599\,
            I => \U712_CHIP_RAM.N_303\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__5596\,
            I => \U712_CHIP_RAM.N_303\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__5591\,
            I => \U712_CHIP_RAM.N_443_cascade_\
        );

    \I__784\ : InMux
    port map (
            O => \N__5588\,
            I => \N__5585\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__5585\,
            I => \U712_CHIP_RAM.N_204\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__5582\,
            I => \U712_CHIP_RAM.N_463_cascade_\
        );

    \I__781\ : CascadeMux
    port map (
            O => \N__5579\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\
        );

    \I__780\ : CascadeMux
    port map (
            O => \N__5576\,
            I => \N__5573\
        );

    \I__779\ : InMux
    port map (
            O => \N__5573\,
            I => \N__5570\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__5570\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__777\ : InMux
    port map (
            O => \N__5567\,
            I => \N__5564\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__5564\,
            I => \N__5561\
        );

    \I__775\ : Span4Mux_v
    port map (
            O => \N__5561\,
            I => \N__5558\
        );

    \I__774\ : Span4Mux_v
    port map (
            O => \N__5558\,
            I => \N__5555\
        );

    \I__773\ : Sp12to4
    port map (
            O => \N__5555\,
            I => \N__5552\
        );

    \I__772\ : Span12Mux_h
    port map (
            O => \N__5552\,
            I => \N__5549\
        );

    \I__771\ : Odrv12
    port map (
            O => \N__5549\,
            I => \A_c_17\
        );

    \I__770\ : CascadeMux
    port map (
            O => \N__5546\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_\
        );

    \I__769\ : InMux
    port map (
            O => \N__5543\,
            I => \N__5540\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__5540\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\
        );

    \I__767\ : InMux
    port map (
            O => \N__5537\,
            I => \N__5534\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__5534\,
            I => \N__5531\
        );

    \I__765\ : Span4Mux_v
    port map (
            O => \N__5531\,
            I => \N__5528\
        );

    \I__764\ : Odrv4
    port map (
            O => \N__5528\,
            I => \U712_CHIP_RAM.N_346\
        );

    \I__763\ : InMux
    port map (
            O => \N__5525\,
            I => \N__5520\
        );

    \I__762\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5515\
        );

    \I__761\ : InMux
    port map (
            O => \N__5523\,
            I => \N__5515\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__5520\,
            I => \U712_CHIP_RAM.N_388\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__5515\,
            I => \U712_CHIP_RAM.N_388\
        );

    \I__758\ : InMux
    port map (
            O => \N__5510\,
            I => \N__5505\
        );

    \I__757\ : CascadeMux
    port map (
            O => \N__5509\,
            I => \N__5501\
        );

    \I__756\ : InMux
    port map (
            O => \N__5508\,
            I => \N__5498\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__5505\,
            I => \N__5495\
        );

    \I__754\ : CascadeMux
    port map (
            O => \N__5504\,
            I => \N__5492\
        );

    \I__753\ : InMux
    port map (
            O => \N__5501\,
            I => \N__5488\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__5498\,
            I => \N__5483\
        );

    \I__751\ : Span4Mux_v
    port map (
            O => \N__5495\,
            I => \N__5483\
        );

    \I__750\ : InMux
    port map (
            O => \N__5492\,
            I => \N__5480\
        );

    \I__749\ : InMux
    port map (
            O => \N__5491\,
            I => \N__5477\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__5488\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__747\ : Odrv4
    port map (
            O => \N__5483\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__5480\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__5477\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__744\ : SRMux
    port map (
            O => \N__5468\,
            I => \N__5465\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__5465\,
            I => \N__5461\
        );

    \I__742\ : InMux
    port map (
            O => \N__5464\,
            I => \N__5458\
        );

    \I__741\ : Span4Mux_h
    port map (
            O => \N__5461\,
            I => \N__5455\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__5458\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__739\ : Odrv4
    port map (
            O => \N__5455\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__738\ : CascadeMux
    port map (
            O => \N__5450\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_cascade_\
        );

    \I__737\ : InMux
    port map (
            O => \N__5447\,
            I => \N__5443\
        );

    \I__736\ : InMux
    port map (
            O => \N__5446\,
            I => \N__5440\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__5443\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__5440\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__733\ : InMux
    port map (
            O => \N__5435\,
            I => \N__5431\
        );

    \I__732\ : IoInMux
    port map (
            O => \N__5434\,
            I => \N__5428\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__5431\,
            I => \N__5425\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__5428\,
            I => \N__5422\
        );

    \I__729\ : Span4Mux_v
    port map (
            O => \N__5425\,
            I => \N__5419\
        );

    \I__728\ : IoSpan4Mux
    port map (
            O => \N__5422\,
            I => \N__5416\
        );

    \I__727\ : Sp12to4
    port map (
            O => \N__5419\,
            I => \N__5413\
        );

    \I__726\ : IoSpan4Mux
    port map (
            O => \N__5416\,
            I => \N__5410\
        );

    \I__725\ : Span12Mux_h
    port map (
            O => \N__5413\,
            I => \N__5407\
        );

    \I__724\ : IoSpan4Mux
    port map (
            O => \N__5410\,
            I => \N__5404\
        );

    \I__723\ : Odrv12
    port map (
            O => \N__5407\,
            I => \C1_c\
        );

    \I__722\ : Odrv4
    port map (
            O => \N__5404\,
            I => \C1_c\
        );

    \I__721\ : InMux
    port map (
            O => \N__5399\,
            I => \N__5396\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__5396\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__719\ : IoInMux
    port map (
            O => \N__5393\,
            I => \N__5390\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__5390\,
            I => \N__5387\
        );

    \I__717\ : IoSpan4Mux
    port map (
            O => \N__5387\,
            I => \N__5384\
        );

    \I__716\ : Span4Mux_s2_v
    port map (
            O => \N__5384\,
            I => \N__5381\
        );

    \I__715\ : Span4Mux_v
    port map (
            O => \N__5381\,
            I => \N__5378\
        );

    \I__714\ : Span4Mux_h
    port map (
            O => \N__5378\,
            I => \N__5375\
        );

    \I__713\ : Odrv4
    port map (
            O => \N__5375\,
            I => \CRCSn_c\
        );

    \I__712\ : IoInMux
    port map (
            O => \N__5372\,
            I => \N__5369\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__5369\,
            I => \N__5366\
        );

    \I__710\ : IoSpan4Mux
    port map (
            O => \N__5366\,
            I => \N__5363\
        );

    \I__709\ : Sp12to4
    port map (
            O => \N__5363\,
            I => \N__5360\
        );

    \I__708\ : Span12Mux_s9_v
    port map (
            O => \N__5360\,
            I => \N__5357\
        );

    \I__707\ : Odrv12
    port map (
            O => \N__5357\,
            I => \RASn_c\
        );

    \I__706\ : IoInMux
    port map (
            O => \N__5354\,
            I => \N__5351\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__5351\,
            I => \N__5348\
        );

    \I__704\ : Span12Mux_s10_v
    port map (
            O => \N__5348\,
            I => \N__5345\
        );

    \I__703\ : Odrv12
    port map (
            O => \N__5345\,
            I => \CMA_c_0\
        );

    \I__702\ : IoInMux
    port map (
            O => \N__5342\,
            I => \N__5339\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__5339\,
            I => \N__5336\
        );

    \I__700\ : Span12Mux_s10_v
    port map (
            O => \N__5336\,
            I => \N__5333\
        );

    \I__699\ : Odrv12
    port map (
            O => \N__5333\,
            I => \CMA_c_10\
        );

    \I__698\ : IoInMux
    port map (
            O => \N__5330\,
            I => \N__5327\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__5327\,
            I => \N__5324\
        );

    \I__696\ : Span12Mux_s10_v
    port map (
            O => \N__5324\,
            I => \N__5321\
        );

    \I__695\ : Odrv12
    port map (
            O => \N__5321\,
            I => \CMA_c_2\
        );

    \I__694\ : IoInMux
    port map (
            O => \N__5318\,
            I => \N__5314\
        );

    \I__693\ : InMux
    port map (
            O => \N__5317\,
            I => \N__5311\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__5314\,
            I => \N__5308\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__5311\,
            I => \N__5305\
        );

    \I__690\ : Span12Mux_s4_v
    port map (
            O => \N__5308\,
            I => \N__5302\
        );

    \I__689\ : Span4Mux_h
    port map (
            O => \N__5305\,
            I => \N__5299\
        );

    \I__688\ : Span12Mux_v
    port map (
            O => \N__5302\,
            I => \N__5296\
        );

    \I__687\ : Span4Mux_v
    port map (
            O => \N__5299\,
            I => \N__5293\
        );

    \I__686\ : Span12Mux_h
    port map (
            O => \N__5296\,
            I => \N__5290\
        );

    \I__685\ : Sp12to4
    port map (
            O => \N__5293\,
            I => \N__5287\
        );

    \I__684\ : Odrv12
    port map (
            O => \N__5290\,
            I => \A_c_9\
        );

    \I__683\ : Odrv12
    port map (
            O => \N__5287\,
            I => \A_c_9\
        );

    \I__682\ : InMux
    port map (
            O => \N__5282\,
            I => \N__5279\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__5279\,
            I => \U712_CYCLE_TERM.N_312\
        );

    \I__680\ : InMux
    port map (
            O => \N__5276\,
            I => \N__5270\
        );

    \I__679\ : InMux
    port map (
            O => \N__5275\,
            I => \N__5270\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__5270\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__677\ : InMux
    port map (
            O => \N__5267\,
            I => \N__5262\
        );

    \I__676\ : InMux
    port map (
            O => \N__5266\,
            I => \N__5257\
        );

    \I__675\ : InMux
    port map (
            O => \N__5265\,
            I => \N__5257\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__5262\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__5257\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__672\ : IoInMux
    port map (
            O => \N__5252\,
            I => \N__5249\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__5249\,
            I => \N__5245\
        );

    \I__670\ : IoInMux
    port map (
            O => \N__5248\,
            I => \N__5242\
        );

    \I__669\ : IoSpan4Mux
    port map (
            O => \N__5245\,
            I => \N__5238\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__5242\,
            I => \N__5235\
        );

    \I__667\ : IoInMux
    port map (
            O => \N__5241\,
            I => \N__5232\
        );

    \I__666\ : Sp12to4
    port map (
            O => \N__5238\,
            I => \N__5229\
        );

    \I__665\ : Span4Mux_s3_v
    port map (
            O => \N__5235\,
            I => \N__5226\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__5232\,
            I => \N__5223\
        );

    \I__663\ : Span12Mux_s7_h
    port map (
            O => \N__5229\,
            I => \N__5220\
        );

    \I__662\ : Sp12to4
    port map (
            O => \N__5226\,
            I => \N__5217\
        );

    \I__661\ : IoSpan4Mux
    port map (
            O => \N__5223\,
            I => \N__5214\
        );

    \I__660\ : Span12Mux_h
    port map (
            O => \N__5220\,
            I => \N__5209\
        );

    \I__659\ : Span12Mux_h
    port map (
            O => \N__5217\,
            I => \N__5209\
        );

    \I__658\ : Sp12to4
    port map (
            O => \N__5214\,
            I => \N__5206\
        );

    \I__657\ : Span12Mux_v
    port map (
            O => \N__5209\,
            I => \N__5200\
        );

    \I__656\ : Span12Mux_h
    port map (
            O => \N__5206\,
            I => \N__5200\
        );

    \I__655\ : InMux
    port map (
            O => \N__5205\,
            I => \N__5197\
        );

    \I__654\ : Odrv12
    port map (
            O => \N__5200\,
            I => \TACK_OUTn\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__5197\,
            I => \TACK_OUTn\
        );

    \I__652\ : InMux
    port map (
            O => \N__5192\,
            I => \N__5189\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__5189\,
            I => \N__5185\
        );

    \I__650\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5182\
        );

    \I__649\ : Span4Mux_v
    port map (
            O => \N__5185\,
            I => \N__5179\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__5182\,
            I => \N__5176\
        );

    \I__647\ : Span4Mux_h
    port map (
            O => \N__5179\,
            I => \N__5171\
        );

    \I__646\ : Span4Mux_v
    port map (
            O => \N__5176\,
            I => \N__5171\
        );

    \I__645\ : Span4Mux_h
    port map (
            O => \N__5171\,
            I => \N__5168\
        );

    \I__644\ : Sp12to4
    port map (
            O => \N__5168\,
            I => \N__5165\
        );

    \I__643\ : Odrv12
    port map (
            O => \N__5165\,
            I => \DBRn_c\
        );

    \I__642\ : InMux
    port map (
            O => \N__5162\,
            I => \N__5159\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__5159\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__640\ : InMux
    port map (
            O => \N__5156\,
            I => \N__5152\
        );

    \I__639\ : InMux
    port map (
            O => \N__5155\,
            I => \N__5149\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__5152\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__5149\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__636\ : InMux
    port map (
            O => \N__5144\,
            I => \N__5136\
        );

    \I__635\ : InMux
    port map (
            O => \N__5143\,
            I => \N__5136\
        );

    \I__634\ : InMux
    port map (
            O => \N__5142\,
            I => \N__5131\
        );

    \I__633\ : InMux
    port map (
            O => \N__5141\,
            I => \N__5131\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__5136\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__5131\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__630\ : CascadeMux
    port map (
            O => \N__5126\,
            I => \N__5123\
        );

    \I__629\ : InMux
    port map (
            O => \N__5123\,
            I => \N__5120\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__5120\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\
        );

    \I__627\ : InMux
    port map (
            O => \N__5117\,
            I => \N__5108\
        );

    \I__626\ : InMux
    port map (
            O => \N__5116\,
            I => \N__5108\
        );

    \I__625\ : InMux
    port map (
            O => \N__5115\,
            I => \N__5108\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__5108\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__623\ : IoInMux
    port map (
            O => \N__5105\,
            I => \N__5102\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__5102\,
            I => \N__5099\
        );

    \I__621\ : IoSpan4Mux
    port map (
            O => \N__5099\,
            I => \N__5096\
        );

    \I__620\ : Span4Mux_s3_h
    port map (
            O => \N__5096\,
            I => \N__5093\
        );

    \I__619\ : Span4Mux_v
    port map (
            O => \N__5093\,
            I => \N__5089\
        );

    \I__618\ : InMux
    port map (
            O => \N__5092\,
            I => \N__5086\
        );

    \I__617\ : Span4Mux_h
    port map (
            O => \N__5089\,
            I => \N__5083\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__5086\,
            I => \N__5080\
        );

    \I__615\ : Sp12to4
    port map (
            O => \N__5083\,
            I => \N__5077\
        );

    \I__614\ : Span4Mux_v
    port map (
            O => \N__5080\,
            I => \N__5074\
        );

    \I__613\ : Span12Mux_h
    port map (
            O => \N__5077\,
            I => \N__5069\
        );

    \I__612\ : Sp12to4
    port map (
            O => \N__5074\,
            I => \N__5069\
        );

    \I__611\ : Span12Mux_h
    port map (
            O => \N__5069\,
            I => \N__5066\
        );

    \I__610\ : Odrv12
    port map (
            O => \N__5066\,
            I => \C3_c\
        );

    \I__609\ : InMux
    port map (
            O => \N__5063\,
            I => \N__5060\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__5060\,
            I => \N__5056\
        );

    \I__607\ : InMux
    port map (
            O => \N__5059\,
            I => \N__5053\
        );

    \I__606\ : Odrv12
    port map (
            O => \N__5056\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__5053\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\
        );

    \I__604\ : IoInMux
    port map (
            O => \N__5048\,
            I => \N__5045\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__5045\,
            I => \N__5042\
        );

    \I__602\ : Span4Mux_s3_v
    port map (
            O => \N__5042\,
            I => \N__5039\
        );

    \I__601\ : Span4Mux_h
    port map (
            O => \N__5039\,
            I => \N__5036\
        );

    \I__600\ : Span4Mux_v
    port map (
            O => \N__5036\,
            I => \N__5033\
        );

    \I__599\ : Span4Mux_v
    port map (
            O => \N__5033\,
            I => \N__5030\
        );

    \I__598\ : Span4Mux_v
    port map (
            O => \N__5030\,
            I => \N__5026\
        );

    \I__597\ : InMux
    port map (
            O => \N__5029\,
            I => \N__5023\
        );

    \I__596\ : Odrv4
    port map (
            O => \N__5026\,
            I => \LATCH_CLK_c\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__5023\,
            I => \LATCH_CLK_c\
        );

    \I__594\ : InMux
    port map (
            O => \N__5018\,
            I => \N__5015\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__5015\,
            I => \N__5012\
        );

    \I__592\ : Span4Mux_h
    port map (
            O => \N__5012\,
            I => \N__5008\
        );

    \I__591\ : InMux
    port map (
            O => \N__5011\,
            I => \N__5005\
        );

    \I__590\ : Span4Mux_h
    port map (
            O => \N__5008\,
            I => \N__5000\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__5005\,
            I => \N__5000\
        );

    \I__588\ : Span4Mux_v
    port map (
            O => \N__5000\,
            I => \N__4997\
        );

    \I__587\ : Sp12to4
    port map (
            O => \N__4997\,
            I => \N__4994\
        );

    \I__586\ : Span12Mux_h
    port map (
            O => \N__4994\,
            I => \N__4991\
        );

    \I__585\ : Span12Mux_v
    port map (
            O => \N__4991\,
            I => \N__4988\
        );

    \I__584\ : Odrv12
    port map (
            O => \N__4988\,
            I => \TSn_c\
        );

    \I__583\ : CascadeMux
    port map (
            O => \N__4985\,
            I => \N__4982\
        );

    \I__582\ : InMux
    port map (
            O => \N__4982\,
            I => \N__4979\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__4979\,
            I => \N__4976\
        );

    \I__580\ : Span4Mux_v
    port map (
            O => \N__4976\,
            I => \N__4973\
        );

    \I__579\ : Sp12to4
    port map (
            O => \N__4973\,
            I => \N__4970\
        );

    \I__578\ : Span12Mux_h
    port map (
            O => \N__4970\,
            I => \N__4967\
        );

    \I__577\ : Span12Mux_v
    port map (
            O => \N__4967\,
            I => \N__4964\
        );

    \I__576\ : Odrv12
    port map (
            O => \N__4964\,
            I => \REGSPACEn_c\
        );

    \I__575\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4958\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__4958\,
            I => \U712_REG_SM.N_414\
        );

    \I__573\ : CascadeMux
    port map (
            O => \N__4955\,
            I => \U712_CYCLE_TERM.N_452_cascade_\
        );

    \I__572\ : InMux
    port map (
            O => \N__4952\,
            I => \N__4949\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__4949\,
            I => \N__4946\
        );

    \I__570\ : Span12Mux_h
    port map (
            O => \N__4946\,
            I => \N__4943\
        );

    \I__569\ : Span12Mux_v
    port map (
            O => \N__4943\,
            I => \N__4940\
        );

    \I__568\ : Odrv12
    port map (
            O => \N__4940\,
            I => \RAMSPACEn_c\
        );

    \I__567\ : CascadeMux
    port map (
            O => \N__4937\,
            I => \U712_CHIP_RAM.N_417_cascade_\
        );

    \I__566\ : InMux
    port map (
            O => \N__4934\,
            I => \N__4929\
        );

    \I__565\ : InMux
    port map (
            O => \N__4933\,
            I => \N__4924\
        );

    \I__564\ : InMux
    port map (
            O => \N__4932\,
            I => \N__4924\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__4929\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__4924\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__561\ : CascadeMux
    port map (
            O => \N__4919\,
            I => \N__4916\
        );

    \I__560\ : InMux
    port map (
            O => \N__4916\,
            I => \N__4913\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__4913\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_1\
        );

    \I__558\ : InMux
    port map (
            O => \N__4910\,
            I => \N__4907\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__4907\,
            I => \U712_CHIP_RAM.N_206\
        );

    \I__556\ : InMux
    port map (
            O => \N__4904\,
            I => \N__4901\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__4901\,
            I => \U712_CHIP_RAM.N_457\
        );

    \I__554\ : InMux
    port map (
            O => \N__4898\,
            I => \N__4895\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__4895\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_5\
        );

    \I__552\ : InMux
    port map (
            O => \N__4892\,
            I => \N__4886\
        );

    \I__551\ : InMux
    port map (
            O => \N__4891\,
            I => \N__4886\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__4886\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\
        );

    \I__549\ : InMux
    port map (
            O => \N__4883\,
            I => \N__4880\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__4880\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_i_1\
        );

    \I__547\ : InMux
    port map (
            O => \N__4877\,
            I => \N__4874\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__4874\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_95_i_a2_i_0\
        );

    \I__545\ : CascadeMux
    port map (
            O => \N__4871\,
            I => \U712_CHIP_RAM.N_556_cascade_\
        );

    \I__544\ : InMux
    port map (
            O => \N__4868\,
            I => \N__4865\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4865\,
            I => \U712_CHIP_RAM.N_202\
        );

    \I__542\ : CascadeMux
    port map (
            O => \N__4862\,
            I => \U712_CHIP_RAM.N_388_cascade_\
        );

    \I__541\ : InMux
    port map (
            O => \N__4859\,
            I => \N__4856\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__4856\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_i_0\
        );

    \I__539\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4849\
        );

    \I__538\ : InMux
    port map (
            O => \N__4852\,
            I => \N__4846\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__4849\,
            I => \N__4843\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4846\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__535\ : Odrv12
    port map (
            O => \N__4843\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__534\ : InMux
    port map (
            O => \N__4838\,
            I => \N__4835\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__4835\,
            I => \N__4832\
        );

    \I__532\ : Odrv4
    port map (
            O => \N__4832\,
            I => \U712_CHIP_RAM.REFRESH5lto7_0\
        );

    \I__531\ : InMux
    port map (
            O => \N__4829\,
            I => \N__4826\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__4826\,
            I => \N__4823\
        );

    \I__529\ : Odrv12
    port map (
            O => \N__4823\,
            I => \U712_CHIP_RAM.REFRESH5lt7\
        );

    \I__528\ : CascadeMux
    port map (
            O => \N__4820\,
            I => \N__4816\
        );

    \I__527\ : InMux
    port map (
            O => \N__4819\,
            I => \N__4810\
        );

    \I__526\ : InMux
    port map (
            O => \N__4816\,
            I => \N__4810\
        );

    \I__525\ : InMux
    port map (
            O => \N__4815\,
            I => \N__4807\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__4810\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4807\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__522\ : CascadeMux
    port map (
            O => \N__4802\,
            I => \N__4798\
        );

    \I__521\ : InMux
    port map (
            O => \N__4801\,
            I => \N__4795\
        );

    \I__520\ : InMux
    port map (
            O => \N__4798\,
            I => \N__4792\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__4795\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__4792\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__517\ : InMux
    port map (
            O => \N__4787\,
            I => \N__4783\
        );

    \I__516\ : InMux
    port map (
            O => \N__4786\,
            I => \N__4780\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__4783\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__4780\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__513\ : InMux
    port map (
            O => \N__4775\,
            I => \N__4772\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__4772\,
            I => \N__4769\
        );

    \I__511\ : Sp12to4
    port map (
            O => \N__4769\,
            I => \N__4766\
        );

    \I__510\ : Span12Mux_v
    port map (
            O => \N__4766\,
            I => \N__4763\
        );

    \I__509\ : Span12Mux_h
    port map (
            O => \N__4763\,
            I => \N__4760\
        );

    \I__508\ : Odrv12
    port map (
            O => \N__4760\,
            I => \A_c_16\
        );

    \I__507\ : CascadeMux
    port map (
            O => \N__4757\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_\
        );

    \I__506\ : InMux
    port map (
            O => \N__4754\,
            I => \N__4750\
        );

    \I__505\ : InMux
    port map (
            O => \N__4753\,
            I => \N__4747\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__4750\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4747\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__502\ : InMux
    port map (
            O => \N__4742\,
            I => \N__4738\
        );

    \I__501\ : InMux
    port map (
            O => \N__4741\,
            I => \N__4735\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4738\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4735\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__498\ : IoInMux
    port map (
            O => \N__4730\,
            I => \N__4727\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__4727\,
            I => \N__4724\
        );

    \I__496\ : IoSpan4Mux
    port map (
            O => \N__4724\,
            I => \N__4721\
        );

    \I__495\ : IoSpan4Mux
    port map (
            O => \N__4721\,
            I => \N__4718\
        );

    \I__494\ : Span4Mux_s2_v
    port map (
            O => \N__4718\,
            I => \N__4714\
        );

    \I__493\ : InMux
    port map (
            O => \N__4717\,
            I => \N__4711\
        );

    \I__492\ : Sp12to4
    port map (
            O => \N__4714\,
            I => \N__4708\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__4711\,
            I => \N__4705\
        );

    \I__490\ : Span12Mux_s8_v
    port map (
            O => \N__4708\,
            I => \N__4702\
        );

    \I__489\ : Span4Mux_h
    port map (
            O => \N__4705\,
            I => \N__4699\
        );

    \I__488\ : Span12Mux_v
    port map (
            O => \N__4702\,
            I => \N__4694\
        );

    \I__487\ : Sp12to4
    port map (
            O => \N__4699\,
            I => \N__4694\
        );

    \I__486\ : Odrv12
    port map (
            O => \N__4694\,
            I => \A_c_10\
        );

    \I__485\ : CascadeMux
    port map (
            O => \N__4691\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\
        );

    \I__484\ : InMux
    port map (
            O => \N__4688\,
            I => \N__4685\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__4685\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\
        );

    \I__482\ : InMux
    port map (
            O => \N__4682\,
            I => \N__4679\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__4679\,
            I => \N__4676\
        );

    \I__480\ : Odrv4
    port map (
            O => \N__4676\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__479\ : IoInMux
    port map (
            O => \N__4673\,
            I => \N__4670\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__4670\,
            I => \N__4667\
        );

    \I__477\ : IoSpan4Mux
    port map (
            O => \N__4667\,
            I => \N__4664\
        );

    \I__476\ : Sp12to4
    port map (
            O => \N__4664\,
            I => \N__4661\
        );

    \I__475\ : Span12Mux_s7_h
    port map (
            O => \N__4661\,
            I => \N__4658\
        );

    \I__474\ : Span12Mux_h
    port map (
            O => \N__4658\,
            I => \N__4655\
        );

    \I__473\ : Odrv12
    port map (
            O => \N__4655\,
            I => \CMA_c_7\
        );

    \I__472\ : IoInMux
    port map (
            O => \N__4652\,
            I => \N__4649\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__4649\,
            I => \N__4646\
        );

    \I__470\ : IoSpan4Mux
    port map (
            O => \N__4646\,
            I => \N__4643\
        );

    \I__469\ : Sp12to4
    port map (
            O => \N__4643\,
            I => \N__4640\
        );

    \I__468\ : Span12Mux_s7_h
    port map (
            O => \N__4640\,
            I => \N__4637\
        );

    \I__467\ : Span12Mux_h
    port map (
            O => \N__4637\,
            I => \N__4634\
        );

    \I__466\ : Odrv12
    port map (
            O => \N__4634\,
            I => \CMA_c_8\
        );

    \I__465\ : InMux
    port map (
            O => \N__4631\,
            I => \N__4628\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__4628\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__463\ : InMux
    port map (
            O => \N__4625\,
            I => \bfn_9_5_0_\
        );

    \I__462\ : InMux
    port map (
            O => \N__4622\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__461\ : InMux
    port map (
            O => \N__4619\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__460\ : InMux
    port map (
            O => \N__4616\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__459\ : InMux
    port map (
            O => \N__4613\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__458\ : InMux
    port map (
            O => \N__4610\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__457\ : InMux
    port map (
            O => \N__4607\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__456\ : InMux
    port map (
            O => \N__4604\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__455\ : ClkMux
    port map (
            O => \N__4601\,
            I => \N__4586\
        );

    \I__454\ : ClkMux
    port map (
            O => \N__4600\,
            I => \N__4586\
        );

    \I__453\ : ClkMux
    port map (
            O => \N__4599\,
            I => \N__4586\
        );

    \I__452\ : ClkMux
    port map (
            O => \N__4598\,
            I => \N__4586\
        );

    \I__451\ : ClkMux
    port map (
            O => \N__4597\,
            I => \N__4586\
        );

    \I__450\ : GlobalMux
    port map (
            O => \N__4586\,
            I => \N__4583\
        );

    \I__449\ : gio2CtrlBuf
    port map (
            O => \N__4583\,
            I => \C1_c_g\
        );

    \I__448\ : InMux
    port map (
            O => \N__4580\,
            I => \N__4576\
        );

    \I__447\ : InMux
    port map (
            O => \N__4579\,
            I => \N__4573\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__4576\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__4573\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__444\ : InMux
    port map (
            O => \N__4568\,
            I => \N__4564\
        );

    \I__443\ : InMux
    port map (
            O => \N__4567\,
            I => \N__4561\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__4564\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__4561\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__440\ : IoInMux
    port map (
            O => \N__4556\,
            I => \N__4553\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__4553\,
            I => \N__4550\
        );

    \I__438\ : Span4Mux_s0_v
    port map (
            O => \N__4550\,
            I => \N__4547\
        );

    \I__437\ : Span4Mux_v
    port map (
            O => \N__4547\,
            I => \N__4544\
        );

    \I__436\ : Span4Mux_v
    port map (
            O => \N__4544\,
            I => \N__4541\
        );

    \I__435\ : Span4Mux_v
    port map (
            O => \N__4541\,
            I => \N__4538\
        );

    \I__434\ : Odrv4
    port map (
            O => \N__4538\,
            I => \CMA_c_1\
        );

    \I__433\ : InMux
    port map (
            O => \N__4535\,
            I => \N__4532\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__4532\,
            I => \U712_CHIP_RAM.N_340\
        );

    \I__431\ : IoInMux
    port map (
            O => \N__4529\,
            I => \N__4526\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__4526\,
            I => \N__4523\
        );

    \I__429\ : IoSpan4Mux
    port map (
            O => \N__4523\,
            I => \N__4520\
        );

    \I__428\ : Span4Mux_s3_h
    port map (
            O => \N__4520\,
            I => \N__4517\
        );

    \I__427\ : Sp12to4
    port map (
            O => \N__4517\,
            I => \N__4514\
        );

    \I__426\ : Span12Mux_s8_h
    port map (
            O => \N__4514\,
            I => \N__4511\
        );

    \I__425\ : Span12Mux_h
    port map (
            O => \N__4511\,
            I => \N__4508\
        );

    \I__424\ : Odrv12
    port map (
            O => \N__4508\,
            I => \CMA_c_5\
        );

    \I__423\ : InMux
    port map (
            O => \N__4505\,
            I => \N__4502\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__4502\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__421\ : CascadeMux
    port map (
            O => \N__4499\,
            I => \U712_CHIP_RAM.N_297_cascade_\
        );

    \I__420\ : InMux
    port map (
            O => \N__4496\,
            I => \N__4493\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__4493\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__418\ : CascadeMux
    port map (
            O => \N__4490\,
            I => \U712_CHIP_RAM.N_196_cascade_\
        );

    \I__417\ : IoInMux
    port map (
            O => \N__4487\,
            I => \N__4483\
        );

    \I__416\ : IoInMux
    port map (
            O => \N__4486\,
            I => \N__4480\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__4483\,
            I => \N__4477\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__4480\,
            I => \N__4474\
        );

    \I__413\ : Span4Mux_s2_v
    port map (
            O => \N__4477\,
            I => \N__4471\
        );

    \I__412\ : IoSpan4Mux
    port map (
            O => \N__4474\,
            I => \N__4468\
        );

    \I__411\ : Span4Mux_h
    port map (
            O => \N__4471\,
            I => \N__4465\
        );

    \I__410\ : Span4Mux_s2_v
    port map (
            O => \N__4468\,
            I => \N__4462\
        );

    \I__409\ : Sp12to4
    port map (
            O => \N__4465\,
            I => \N__4458\
        );

    \I__408\ : Span4Mux_h
    port map (
            O => \N__4462\,
            I => \N__4455\
        );

    \I__407\ : IoInMux
    port map (
            O => \N__4461\,
            I => \N__4452\
        );

    \I__406\ : Span12Mux_h
    port map (
            O => \N__4458\,
            I => \N__4447\
        );

    \I__405\ : Sp12to4
    port map (
            O => \N__4455\,
            I => \N__4447\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__4452\,
            I => \N__4444\
        );

    \I__403\ : Span12Mux_v
    port map (
            O => \N__4447\,
            I => \N__4438\
        );

    \I__402\ : Span12Mux_s11_h
    port map (
            O => \N__4444\,
            I => \N__4438\
        );

    \I__401\ : InMux
    port map (
            O => \N__4443\,
            I => \N__4435\
        );

    \I__400\ : Odrv12
    port map (
            O => \N__4438\,
            I => \TACK_EN\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__4435\,
            I => \TACK_EN\
        );

    \I__398\ : IoInMux
    port map (
            O => \N__4430\,
            I => \N__4427\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__4427\,
            I => \N__4424\
        );

    \I__396\ : Span12Mux_s6_v
    port map (
            O => \N__4424\,
            I => \N__4421\
        );

    \I__395\ : Odrv12
    port map (
            O => \N__4421\,
            I => \CLK80_PLL_i_i\
        );

    \I__394\ : IoInMux
    port map (
            O => \N__4418\,
            I => \N__4415\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__4415\,
            I => \N__4412\
        );

    \I__392\ : Span4Mux_s3_h
    port map (
            O => \N__4412\,
            I => \N__4409\
        );

    \I__391\ : Odrv4
    port map (
            O => \N__4409\,
            I => \DBRn_c_i_0\
        );

    \I__390\ : IoInMux
    port map (
            O => \N__4406\,
            I => \N__4403\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__4403\,
            I => \N__4400\
        );

    \I__388\ : Span12Mux_s3_v
    port map (
            O => \N__4400\,
            I => \N__4397\
        );

    \I__387\ : Odrv12
    port map (
            O => \N__4397\,
            I => \VBENn_c\
        );

    \I__386\ : InMux
    port map (
            O => \N__4394\,
            I => \N__4391\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__4391\,
            I => \N__4388\
        );

    \I__384\ : Span4Mux_h
    port map (
            O => \N__4388\,
            I => \N__4385\
        );

    \I__383\ : Sp12to4
    port map (
            O => \N__4385\,
            I => \N__4382\
        );

    \I__382\ : Span12Mux_v
    port map (
            O => \N__4382\,
            I => \N__4379\
        );

    \I__381\ : Odrv12
    port map (
            O => \N__4379\,
            I => \A_c_14\
        );

    \I__380\ : IoInMux
    port map (
            O => \N__4376\,
            I => \N__4373\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__4373\,
            I => \N__4370\
        );

    \I__378\ : IoSpan4Mux
    port map (
            O => \N__4370\,
            I => \N__4367\
        );

    \I__377\ : Span4Mux_s2_v
    port map (
            O => \N__4367\,
            I => \N__4364\
        );

    \I__376\ : Sp12to4
    port map (
            O => \N__4364\,
            I => \N__4361\
        );

    \I__375\ : Span12Mux_v
    port map (
            O => \N__4361\,
            I => \N__4358\
        );

    \I__374\ : Odrv12
    port map (
            O => \N__4358\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            I => \N__4600\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            I => \N__4597\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__4598\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__4599\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_9_0_\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_10_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_12_0_\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5434\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8636\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4418\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5105\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10274\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10736\,
            in2 => \_gnd_net_\,
            in3 => \N__8725\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBRn_ibuf_RNIBAB_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5188\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_0_a2_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__10042\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10126\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4394\,
            in1 => \N__10041\,
            in2 => \_gnd_net_\,
            in3 => \N__9032\,
            lcout => \U712_CHIP_RAM.N_340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4505\,
            in1 => \N__4496\,
            in2 => \_gnd_net_\,
            in3 => \N__4688\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10246\,
            ce => \N__11217\,
            sr => \N__10700\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__8549\,
            in1 => \N__4535\,
            in2 => \N__9225\,
            in3 => \N__5537\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10246\,
            ce => \N__11217\,
            sr => \N__10700\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100001111"
        )
    port map (
            in0 => \N__10050\,
            in1 => \N__8768\,
            in2 => \N__9226\,
            in3 => \N__8548\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5668\,
            in2 => \_gnd_net_\,
            in3 => \N__6889\,
            lcout => \U712_CHIP_RAM.N_297\,
            ltout => \U712_CHIP_RAM.N_297_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000001111"
        )
    port map (
            in0 => \N__10051\,
            in1 => \N__8767\,
            in2 => \N__4499\,
            in3 => \N__9214\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__4883\,
            in1 => \N__7599\,
            in2 => \N__7703\,
            in3 => \N__4859\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_196_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101111"
        )
    port map (
            in0 => \N__5871\,
            in1 => \N__5738\,
            in2 => \N__4490\,
            in3 => \N__8139\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10253\,
            ce => 'H',
            sr => \N__10687\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110100"
        )
    port map (
            in0 => \N__7468\,
            in1 => \N__7598\,
            in2 => \N__8051\,
            in3 => \N__7329\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4877\,
            in1 => \N__5602\,
            in2 => \_gnd_net_\,
            in3 => \N__6479\,
            lcout => \U712_CHIP_RAM.N_202\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011111111"
        )
    port map (
            in0 => \N__5155\,
            in1 => \N__4443\,
            in2 => \_gnd_net_\,
            in3 => \N__5282\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10267\,
            ce => 'H',
            sr => \N__10667\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4631\,
            in2 => \_gnd_net_\,
            in3 => \N__4625\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_9_5_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__4601\,
            ce => 'H',
            sr => \N__5468\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4568\,
            in2 => \_gnd_net_\,
            in3 => \N__4622\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__4601\,
            ce => 'H',
            sr => \N__5468\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4787\,
            in2 => \_gnd_net_\,
            in3 => \N__4619\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__4601\,
            ce => 'H',
            sr => \N__5468\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4580\,
            in2 => \_gnd_net_\,
            in3 => \N__4616\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__4601\,
            ce => 'H',
            sr => \N__5468\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4801\,
            in2 => \_gnd_net_\,
            in3 => \N__4613\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__4601\,
            ce => 'H',
            sr => \N__5468\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4742\,
            in2 => \_gnd_net_\,
            in3 => \N__4610\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__4601\,
            ce => 'H',
            sr => \N__5468\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4754\,
            in2 => \_gnd_net_\,
            in3 => \N__4607\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__4601\,
            ce => 'H',
            sr => \N__5468\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4852\,
            in2 => \_gnd_net_\,
            in3 => \N__4604\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4601\,
            ce => 'H',
            sr => \N__5468\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__4579\,
            in1 => \N__4567\,
            in2 => \N__4802\,
            in3 => \N__4786\,
            lcout => \U712_CHIP_RAM.REFRESH5lt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4775\,
            in1 => \N__7097\,
            in2 => \_gnd_net_\,
            in3 => \N__9167\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9169\,
            in1 => \N__10029\,
            in2 => \N__4757\,
            in3 => \N__8741\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4753\,
            in2 => \_gnd_net_\,
            in3 => \N__4741\,
            lcout => \U712_CHIP_RAM.REFRESH5lto7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4717\,
            in1 => \N__7214\,
            in2 => \_gnd_net_\,
            in3 => \N__9166\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9168\,
            in1 => \N__10028\,
            in2 => \N__4691\,
            in3 => \N__8822\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__8550\,
            in1 => \N__8831\,
            in2 => \N__8521\,
            in3 => \N__4682\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10240\,
            ce => \N__11195\,
            sr => \N__10695\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__8551\,
            in1 => \N__8753\,
            in2 => \N__8522\,
            in3 => \N__5543\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10240\,
            ce => \N__11195\,
            sr => \N__10695\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5667\,
            in1 => \N__9137\,
            in2 => \N__6897\,
            in3 => \N__5491\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__4910\,
            in1 => \N__5523\,
            in2 => \N__6901\,
            in3 => \N__5637\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011101010"
        )
    port map (
            in0 => \N__8038\,
            in1 => \N__7589\,
            in2 => \N__8153\,
            in3 => \N__7323\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_95_i_a2_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__5588\,
            in1 => \N__5524\,
            in2 => \N__5509\,
            in3 => \N__5638\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000101"
        )
    port map (
            in0 => \N__6967\,
            in1 => \N__5063\,
            in2 => \N__4820\,
            in3 => \N__4934\,
            lcout => \U712_CHIP_RAM.N_556\,
            ltout => \U712_CHIP_RAM.N_556_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_0_2_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__10567\,
            in1 => \N__8039\,
            in2 => \N__4871\,
            in3 => \N__6455\,
            lcout => \U712_CHIP_RAM.N_388\,
            ltout => \U712_CHIP_RAM.N_388_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__5636\,
            in1 => \N__4868\,
            in2 => \N__4862\,
            in3 => \N__5671\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000010"
        )
    port map (
            in0 => \N__7588\,
            in1 => \N__4819\,
            in2 => \N__8050\,
            in3 => \N__6968\,
            lcout => \U712_CHIP_RAM.N_445\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010110010111"
        )
    port map (
            in0 => \N__8150\,
            in1 => \N__7897\,
            in2 => \N__7333\,
            in3 => \N__7469\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__4815\,
            in1 => \N__5059\,
            in2 => \_gnd_net_\,
            in3 => \N__4932\,
            lcout => \U712_CHIP_RAM.N_551\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010110000"
        )
    port map (
            in0 => \N__4853\,
            in1 => \N__4838\,
            in2 => \N__10568\,
            in3 => \N__4829\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10250\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIMM5O1_3_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__7587\,
            in1 => \N__7324\,
            in2 => \N__7905\,
            in3 => \N__8149\,
            lcout => \U712_CHIP_RAM.N_303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000001000"
        )
    port map (
            in0 => \N__6984\,
            in1 => \N__10562\,
            in2 => \N__11174\,
            in3 => \N__4904\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10250\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10052\,
            in2 => \_gnd_net_\,
            in3 => \N__4933\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_417_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000000"
        )
    port map (
            in0 => \N__4952\,
            in1 => \N__5018\,
            in2 => \N__4937\,
            in3 => \N__10561\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10250\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__10563\,
            in1 => \N__6278\,
            in2 => \N__4919\,
            in3 => \N__7699\,
            lcout => \U712_CHIP_RAM.N_206\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__4898\,
            in1 => \N__4891\,
            in2 => \_gnd_net_\,
            in3 => \N__5941\,
            lcout => \U712_CHIP_RAM.N_457\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_5_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10560\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4892\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10254\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_4_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10559\,
            in2 => \_gnd_net_\,
            in3 => \N__7715\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10254\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__10049\,
            in1 => \N__5783\,
            in2 => \_gnd_net_\,
            in3 => \N__7385\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100000000"
        )
    port map (
            in0 => \N__5942\,
            in1 => \N__5847\,
            in2 => \N__5753\,
            in3 => \N__10558\,
            lcout => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10254\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__11168\,
            in1 => \N__5765\,
            in2 => \N__7334\,
            in3 => \N__5029\,
            lcout => \LATCH_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10257\,
            ce => 'H',
            sr => \N__10670\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10549\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6629\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000100"
        )
    port map (
            in0 => \N__5011\,
            in1 => \N__10550\,
            in2 => \N__4985\,
            in3 => \N__4961\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5276\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10553\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__5446\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6093\,
            lcout => \U712_REG_SM.N_414\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010011"
        )
    port map (
            in0 => \N__5116\,
            in1 => \N__5141\,
            in2 => \N__5885\,
            in3 => \N__6542\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_452_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__10551\,
            in1 => \N__9528\,
            in2 => \N__4955\,
            in3 => \N__5117\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__9527\,
            in1 => \N__10552\,
            in2 => \_gnd_net_\,
            in3 => \N__5142\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__6541\,
            in1 => \N__5881\,
            in2 => \_gnd_net_\,
            in3 => \N__5115\,
            lcout => \U712_CYCLE_TERM.N_312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5266\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10554\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5265\,
            in2 => \_gnd_net_\,
            in3 => \N__5275\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111000100"
        )
    port map (
            in0 => \N__5144\,
            in1 => \N__5205\,
            in2 => \N__9530\,
            in3 => \N__5267\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10268\,
            ce => 'H',
            sr => \N__10665\
        );

    \U712_REG_SM.C1_SYNC_1_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5399\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10268\,
            ce => 'H',
            sr => \N__10665\
        );

    \DBR_SYNC_0_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5192\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10268\,
            ce => 'H',
            sr => \N__10665\
        );

    \DBR_SYNC_1_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5162\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10268\,
            ce => 'H',
            sr => \N__10665\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001000100010"
        )
    port map (
            in0 => \N__5156\,
            in1 => \N__5143\,
            in2 => \N__5126\,
            in3 => \N__5855\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10268\,
            ce => 'H',
            sr => \N__10665\
        );

    \U712_REG_SM.C3_SYNC_0_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5092\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10268\,
            ce => 'H',
            sr => \N__10665\
        );

    \U712_REG_SM.START_RST_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__6618\,
            in1 => \N__5447\,
            in2 => \_gnd_net_\,
            in3 => \N__8342\,
            lcout => \U712_REG_SM.START_RSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10268\,
            ce => 'H',
            sr => \N__10665\
        );

    \U712_REG_SM.REGENn_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010011010100010"
        )
    port map (
            in0 => \N__6124\,
            in1 => \N__6107\,
            in2 => \N__9365\,
            in3 => \N__6737\,
            lcout => \REGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10269\,
            ce => 'H',
            sr => \N__10664\
        );

    \U712_REG_SM.C1_SYNC_0_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5435\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10269\,
            ce => 'H',
            sr => \N__10664\
        );

    \U712_CHIP_RAM.CRCSn_LC_10_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5510\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10225\,
            ce => 'H',
            sr => \N__10707\
        );

    \U712_CHIP_RAM.RASn_LC_10_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5678\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10229\,
            ce => 'H',
            sr => \N__10703\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__8511\,
            in1 => \N__8569\,
            in2 => \N__5576\,
            in3 => \N__8885\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10232\,
            ce => \N__11207\,
            sr => \N__10701\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__9224\,
            in1 => \N__5508\,
            in2 => \_gnd_net_\,
            in3 => \N__8570\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10232\,
            ce => \N__11207\,
            sr => \N__10701\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__8571\,
            in1 => \N__8512\,
            in2 => \N__8984\,
            in3 => \N__6266\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10232\,
            ce => \N__11207\,
            sr => \N__10701\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6752\,
            in1 => \N__5317\,
            in2 => \_gnd_net_\,
            in3 => \N__9162\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9164\,
            in1 => \N__10000\,
            in2 => \N__5579\,
            in3 => \N__8423\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5567\,
            in1 => \N__6193\,
            in2 => \_gnd_net_\,
            in3 => \N__9163\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9165\,
            in1 => \N__10001\,
            in2 => \N__5546\,
            in3 => \N__8702\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7154\,
            in1 => \N__9999\,
            in2 => \_gnd_net_\,
            in3 => \N__8792\,
            lcout => \U712_CHIP_RAM.N_346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__9152\,
            in1 => \N__5639\,
            in2 => \N__5612\,
            in3 => \N__5525\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10238\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__5669\,
            in1 => \N__9150\,
            in2 => \N__5504\,
            in3 => \N__5464\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_CMA25_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10734\,
            in1 => \_gnd_net_\,
            in2 => \N__5450\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_CMA25_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10735\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7485\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__6985\,
            in1 => \N__7420\,
            in2 => \N__7489\,
            in3 => \N__7628\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10733\,
            in1 => \_gnd_net_\,
            in2 => \N__5681\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_10_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__5670\,
            in1 => \N__9151\,
            in2 => \_gnd_net_\,
            in3 => \N__6890\,
            lcout => \U712_CHIP_RAM.CMA_5_i_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIEVI78_3_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__10548\,
            in1 => \N__7906\,
            in2 => \N__6338\,
            in3 => \N__6500\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__6325\,
            in1 => \N__6485\,
            in2 => \N__5621\,
            in3 => \N__6474\,
            lcout => \U712_CHIP_RAM.N_208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__7576\,
            in1 => \_gnd_net_\,
            in2 => \N__8152\,
            in3 => \N__8022\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_443_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6326\,
            in1 => \N__5603\,
            in2 => \N__5591\,
            in3 => \N__6475\,
            lcout => \U712_CHIP_RAM.N_204\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_0_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7467\,
            in2 => \_gnd_net_\,
            in3 => \N__8021\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_0_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__7675\,
            in1 => \N__6363\,
            in2 => \N__6312\,
            in3 => \N__7575\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI05TJ3_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__7574\,
            in1 => \N__6301\,
            in2 => \N__8151\,
            in3 => \N__7676\,
            lcout => \U712_CHIP_RAM.N_463\,
            ltout => \U712_CHIP_RAM.N_463_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIU7TF5_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__8020\,
            in1 => \N__6966\,
            in2 => \N__5582\,
            in3 => \N__6253\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__7590\,
            in1 => \N__6509\,
            in2 => \N__7349\,
            in3 => \N__7684\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10730\,
            in1 => \_gnd_net_\,
            in2 => \N__5741\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI9UML3_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__11131\,
            in1 => \N__7376\,
            in2 => \_gnd_net_\,
            in3 => \N__6499\,
            lcout => \U712_CHIP_RAM.N_418\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__7685\,
            in1 => \N__10059\,
            in2 => \N__6316\,
            in3 => \N__8043\,
            lcout => \U712_CHIP_RAM.N_439\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__7591\,
            in1 => \N__6347\,
            in2 => \_gnd_net_\,
            in3 => \N__10545\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10248\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6986\,
            in1 => \N__8042\,
            in2 => \_gnd_net_\,
            in3 => \N__6454\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIMAOKC_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__5729\,
            in1 => \N__5776\,
            in2 => \N__5723\,
            in3 => \N__7623\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10731\,
            in1 => \_gnd_net_\,
            in2 => \N__5720\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__6368\,
            in1 => \_gnd_net_\,
            in2 => \N__7907\,
            in3 => \N__7328\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10251\,
            ce => \N__5693\,
            sr => \N__10671\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110011"
        )
    port map (
            in0 => \N__7466\,
            in1 => \N__8041\,
            in2 => \_gnd_net_\,
            in3 => \N__7901\,
            lcout => \U712_CHIP_RAM.N_360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__7421\,
            in1 => \N__5777\,
            in2 => \_gnd_net_\,
            in3 => \N__7627\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_2_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__5841\,
            in1 => \N__10412\,
            in2 => \N__5990\,
            in3 => \N__5937\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10255\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__6575\,
            in1 => \N__6156\,
            in2 => \N__5848\,
            in3 => \N__8299\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_400_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000010"
        )
    port map (
            in0 => \N__10413\,
            in1 => \N__8303\,
            in2 => \N__5759\,
            in3 => \N__9364\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10255\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5971\,
            in1 => \N__6001\,
            in2 => \N__5900\,
            in3 => \N__5936\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5954\,
            in2 => \N__5756\,
            in3 => \N__5837\,
            lcout => \U712_CHIP_RAM.N_405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5896\,
            in2 => \N__5798\,
            in3 => \N__5797\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_10_12_0_\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5953\,
            in2 => \_gnd_net_\,
            in3 => \N__5744\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6002\,
            in2 => \_gnd_net_\,
            in3 => \N__5981\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5972\,
            in2 => \_gnd_net_\,
            in3 => \N__5978\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_3_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__5939\,
            in1 => \N__10489\,
            in2 => \N__5975\,
            in3 => \N__5846\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10258\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_1_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__10488\,
            in1 => \N__5940\,
            in2 => \N__5849\,
            in3 => \N__5960\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10258\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_0_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__5938\,
            in1 => \N__5845\,
            in2 => \N__5909\,
            in3 => \N__10487\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10258\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIH4AH_1_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8280\,
            in2 => \_gnd_net_\,
            in3 => \N__5819\,
            lcout => \U712_REG_SM.N_311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6728\,
            in1 => \N__6094\,
            in2 => \N__8297\,
            in3 => \N__9326\,
            lcout => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__6531\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5880\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_RNITKK4_1_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5818\,
            lcout => \DBR_SYNC_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9325\,
            in2 => \_gnd_net_\,
            in3 => \N__8275\,
            lcout => \U712_REG_SM.N_307\,
            ltout => \U712_REG_SM.N_307_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_1_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__8220\,
            in1 => \N__10112\,
            in2 => \N__6161\,
            in3 => \N__6077\,
            lcout => \U712_REG_SM.REG_CYCLE_5_iv_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIJUGT_3_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__8276\,
            in1 => \N__9327\,
            in2 => \_gnd_net_\,
            in3 => \N__6158\,
            lcout => \U712_REG_SM.N_553\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6076\,
            in1 => \N__6157\,
            in2 => \_gnd_net_\,
            in3 => \N__8221\,
            lcout => \U712_REG_SM.N_322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_RNO_0_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__6100\,
            in1 => \N__8338\,
            in2 => \N__8298\,
            in3 => \N__6123\,
            lcout => \U712_REG_SM.REGENn_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100000000"
        )
    port map (
            in0 => \N__6101\,
            in1 => \N__8284\,
            in2 => \N__9352\,
            in3 => \N__6729\,
            lcout => \U712_REG_SM.STATE_COUNTsr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.WRITE_CYCLE_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__9808\,
            in1 => \N__6075\,
            in2 => \_gnd_net_\,
            in3 => \N__6620\,
            lcout => \U712_REG_SM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10270\,
            ce => 'H',
            sr => \N__10661\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__6059\,
            in1 => \N__7070\,
            in2 => \N__9209\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__6037\,
            in1 => \N__7181\,
            in2 => \N__9210\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9220\,
            in1 => \N__9993\,
            in2 => \N__6269\,
            in3 => \N__9668\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9992\,
            in2 => \_gnd_net_\,
            in3 => \N__9173\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6997\,
            in1 => \N__6179\,
            in2 => \_gnd_net_\,
            in3 => \N__6260\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10233\,
            ce => \N__6242\,
            sr => \N__10688\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_0_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6229\,
            in2 => \_gnd_net_\,
            in3 => \N__10732\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_1_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7980\,
            in2 => \_gnd_net_\,
            in3 => \N__8124\,
            lcout => \U712_CHIP_RAM.N_302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__6230\,
            in1 => \N__6215\,
            in2 => \N__10997\,
            in3 => \N__6194\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10236\,
            ce => 'H',
            sr => \N__10680\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_1_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__7692\,
            in1 => \N__6308\,
            in2 => \_gnd_net_\,
            in3 => \N__8125\,
            lcout => \U712_CHIP_RAM.N_555\,
            ltout => \U712_CHIP_RAM.N_555_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__7981\,
            in1 => \_gnd_net_\,
            in2 => \N__6182\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER16\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100111011101110"
        )
    port map (
            in0 => \N__6173\,
            in1 => \N__11046\,
            in2 => \N__6164\,
            in3 => \N__8432\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10236\,
            ce => 'H',
            sr => \N__10680\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_2_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__6457\,
            in1 => \N__8005\,
            in2 => \N__6380\,
            in3 => \N__10547\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6364\,
            in1 => \N__7378\,
            in2 => \_gnd_net_\,
            in3 => \N__7683\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOV791_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__7580\,
            in1 => \N__8004\,
            in2 => \_gnd_net_\,
            in3 => \N__8118\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_355_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__10546\,
            in1 => \N__7377\,
            in2 => \N__6341\,
            in3 => \N__7682\,
            lcout => \U712_CHIP_RAM.N_389\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7873\,
            in2 => \_gnd_net_\,
            in3 => \N__7285\,
            lcout => \U712_CHIP_RAM.N_289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8007\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6456\,
            lcout => \U712_CHIP_RAM.N_387\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_0_3_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7872\,
            in2 => \_gnd_net_\,
            in3 => \N__7286\,
            lcout => \U712_CHIP_RAM.N_293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNILL5O1_0_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000001010"
        )
    port map (
            in0 => \N__8006\,
            in1 => \N__8119\,
            in2 => \N__7308\,
            in3 => \N__7581\,
            lcout => \U712_CHIP_RAM.N_301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111110000"
        )
    port map (
            in0 => \N__8116\,
            in1 => \N__8000\,
            in2 => \N__6317\,
            in3 => \N__7570\,
            lcout => \U712_CHIP_RAM.N_356\,
            ltout => \U712_CHIP_RAM.N_356_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_RNO_2_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__7875\,
            in1 => \N__7291\,
            in2 => \N__6512\,
            in3 => \N__7677\,
            lcout => \U712_CHIP_RAM.N_448\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__7801\,
            in1 => \N__7816\,
            in2 => \N__7754\,
            in3 => \N__7831\,
            lcout => \U712_CHIP_RAM.N_288\,
            ltout => \U712_CHIP_RAM.N_288_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__7569\,
            in1 => \_gnd_net_\,
            in2 => \N__6503\,
            in3 => \N__8115\,
            lcout => \U712_CHIP_RAM.N_473\,
            ltout => \U712_CHIP_RAM.N_473_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_3_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__7290\,
            in1 => \_gnd_net_\,
            in2 => \N__6488\,
            in3 => \N__7874\,
            lcout => \U712_CHIP_RAM.N_557\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100010100"
        )
    port map (
            in0 => \N__7876\,
            in1 => \N__7293\,
            in2 => \N__7592\,
            in3 => \N__8117\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001000000000"
        )
    port map (
            in0 => \N__6422\,
            in1 => \N__7040\,
            in2 => \N__11670\,
            in3 => \N__10509\,
            lcout => \DMA_WRITE_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10241\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIS5F93_0_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101011101"
        )
    port map (
            in0 => \N__10510\,
            in1 => \N__7292\,
            in2 => \N__8034\,
            in3 => \N__7678\,
            lcout => \U712_CHIP_RAM.N_362\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6996\,
            in1 => \N__8040\,
            in2 => \_gnd_net_\,
            in3 => \N__6461\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10249\,
            ce => \N__6431\,
            sr => \N__10668\
        );

    \U712_CHIP_RAM.DBDIR_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__7032\,
            in1 => \N__6391\,
            in2 => \_gnd_net_\,
            in3 => \N__6421\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10252\,
            ce => 'H',
            sr => \N__10666\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__11163\,
            in1 => \N__11748\,
            in2 => \_gnd_net_\,
            in3 => \N__11062\,
            lcout => \U712_BYTE_ENABLE.N_451\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__10486\,
            in1 => \N__9901\,
            in2 => \_gnd_net_\,
            in3 => \N__11749\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10256\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9370\,
            in2 => \_gnd_net_\,
            in3 => \N__8294\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_306_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__8337\,
            in1 => \N__6619\,
            in2 => \N__6599\,
            in3 => \N__10491\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10259\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_0_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__8228\,
            in1 => \N__6586\,
            in2 => \N__9380\,
            in3 => \N__6573\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_399_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__10113\,
            in1 => \N__10490\,
            in2 => \N__6596\,
            in3 => \N__6593\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10259\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100011111101"
        )
    port map (
            in0 => \N__8336\,
            in1 => \N__8295\,
            in2 => \N__9379\,
            in3 => \N__6574\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_353_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100000000"
        )
    port map (
            in0 => \N__6587\,
            in1 => \N__9377\,
            in2 => \N__6578\,
            in3 => \N__10492\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10259\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_1_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6557\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10263\,
            ce => 'H',
            sr => \N__10662\
        );

    \U712_REG_SM.REG_TACK_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__6680\,
            in1 => \N__6707\,
            in2 => \N__6540\,
            in3 => \N__6548\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10263\,
            ce => 'H',
            sr => \N__10662\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__6743\,
            in1 => \N__6695\,
            in2 => \_gnd_net_\,
            in3 => \N__8225\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10263\,
            ce => 'H',
            sr => \N__10662\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111110"
        )
    port map (
            in0 => \N__6730\,
            in1 => \N__6661\,
            in2 => \N__8226\,
            in3 => \N__6693\,
            lcout => \U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10505\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6668\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_RNO_0_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__11534\,
            in1 => \N__11375\,
            in2 => \N__9809\,
            in3 => \N__11465\,
            lcout => \U712_REG_SM.N_432\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_7_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10507\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6653\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_8_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__6701\,
            in1 => \N__10508\,
            in2 => \N__8227\,
            in3 => \N__6694\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10504\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6679\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10506\,
            in2 => \_gnd_net_\,
            in3 => \N__6662\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.N_130_i_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__11677\,
            in1 => \N__9894\,
            in2 => \_gnd_net_\,
            in3 => \N__11750\,
            lcout => \N_130_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WEn_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6902\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10226\,
            ce => 'H',
            sr => \N__10694\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__10010\,
            in1 => \N__9217\,
            in2 => \N__6839\,
            in3 => \N__8810\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6830\,
            in1 => \N__6776\,
            in2 => \_gnd_net_\,
            in3 => \N__9216\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9218\,
            in1 => \N__10012\,
            in2 => \N__6818\,
            in3 => \N__8801\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9215\,
            in1 => \N__6815\,
            in2 => \_gnd_net_\,
            in3 => \N__7124\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__10011\,
            in1 => \N__8780\,
            in2 => \N__6800\,
            in3 => \N__9219\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6797\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10227\,
            ce => \N__7060\,
            sr => \N__10686\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6770\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10228\,
            ce => \N__7064\,
            sr => \N__10679\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7238\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10228\,
            ce => \N__7064\,
            sr => \N__10679\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7202\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10228\,
            ce => \N__7064\,
            sr => \N__10679\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7175\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10228\,
            ce => \N__7064\,
            sr => \N__10679\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7145\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10228\,
            ce => \N__7064\,
            sr => \N__10679\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7118\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10228\,
            ce => \N__7064\,
            sr => \N__10679\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7085\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10228\,
            ce => \N__7064\,
            sr => \N__10679\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__7036\,
            in1 => \N__9821\,
            in2 => \_gnd_net_\,
            in3 => \N__6998\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10231\,
            ce => \N__6929\,
            sr => \N__10673\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI324S_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7983\,
            in1 => \N__11153\,
            in2 => \_gnd_net_\,
            in3 => \N__7600\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_294_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI8MK44_1_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__8114\,
            in1 => \N__7374\,
            in2 => \N__7706\,
            in3 => \N__7686\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_469_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVM119_1_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110011"
        )
    port map (
            in0 => \N__7419\,
            in1 => \N__10428\,
            in2 => \N__7631\,
            in3 => \N__7622\,
            lcout => \U712_CHIP_RAM.N_309\,
            ltout => \U712_CHIP_RAM.N_309_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIUJS3D_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111100"
        )
    port map (
            in0 => \N__7601\,
            in1 => \N__7514\,
            in2 => \N__7508\,
            in3 => \N__7984\,
            lcout => \U712_CHIP_RAM.N_200\,
            ltout => \U712_CHIP_RAM.N_200_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000111010"
        )
    port map (
            in0 => \N__7247\,
            in1 => \N__7505\,
            in2 => \N__7499\,
            in3 => \N__7496\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10235\,
            ce => \N__7739\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__10427\,
            in1 => \N__7490\,
            in2 => \N__7919\,
            in3 => \N__7783\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10235\,
            ce => \N__7739\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7982\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7442\,
            lcout => \U712_CHIP_RAM.N_285\,
            ltout => \U712_CHIP_RAM.N_285_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_RNO_3_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8113\,
            in1 => \N__10016\,
            in2 => \N__7388\,
            in3 => \N__7375\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_a2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7307\,
            in2 => \_gnd_net_\,
            in3 => \N__7241\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7784\,
            in1 => \N__8120\,
            in2 => \_gnd_net_\,
            in3 => \N__8054\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__10237\,
            ce => \N__7732\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8016\,
            in2 => \_gnd_net_\,
            in3 => \N__7910\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7785\,
            in1 => \N__7888\,
            in2 => \_gnd_net_\,
            in3 => \N__7835\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__10237\,
            ce => \N__7732\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7781\,
            in1 => \N__7832\,
            in2 => \_gnd_net_\,
            in3 => \N__7820\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__10237\,
            ce => \N__7732\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7786\,
            in1 => \N__7817\,
            in2 => \_gnd_net_\,
            in3 => \N__7805\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__10237\,
            ce => \N__7732\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7782\,
            in1 => \N__7802\,
            in2 => \_gnd_net_\,
            in3 => \N__7790\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__10237\,
            ce => \N__7732\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7787\,
            in1 => \N__7753\,
            in2 => \_gnd_net_\,
            in3 => \N__7757\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10237\,
            ce => \N__7732\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_1_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10424\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10286\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10239\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_3_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10426\,
            in2 => \_gnd_net_\,
            in3 => \N__8405\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10239\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_2_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10425\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8411\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10239\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_211_i_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__8351\,
            in1 => \N__11610\,
            in2 => \N__9395\,
            in3 => \N__8399\,
            lcout => \N_211_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__11744\,
            in1 => \N__11164\,
            in2 => \_gnd_net_\,
            in3 => \N__11078\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_410_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_148_i_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001101"
        )
    port map (
            in0 => \N__8350\,
            in1 => \N__11609\,
            in2 => \N__8372\,
            in3 => \N__9391\,
            lcout => \N_148_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__10069\,
            in1 => \N__11530\,
            in2 => \_gnd_net_\,
            in3 => \N__11379\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_a2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI3HF31_1_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__8329\,
            in1 => \N__9345\,
            in2 => \N__8296\,
            in3 => \N__8213\,
            lcout => \U712_REG_SM.N_95\,
            ltout => \U712_REG_SM.N_95_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_RNO_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10729\,
            in1 => \_gnd_net_\,
            in2 => \N__8183\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.N_95_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__8164\,
            in1 => \N__8681\,
            in2 => \N__9378\,
            in3 => \N__8180\,
            lcout => \LDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10261\,
            ce => 'H',
            sr => \N__10657\
        );

    \U712_REG_SM.UDSn_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__8642\,
            in1 => \N__8680\,
            in2 => \N__8659\,
            in3 => \N__9369\,
            lcout => \UDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10261\,
            ce => 'H',
            sr => \N__10657\
        );

    \U712_REG_SM.UDSn_RNO_0_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__9810\,
            in1 => \N__11506\,
            in2 => \N__11381\,
            in3 => \N__11466\,
            lcout => \U712_REG_SM.N_433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10469\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__8504\,
            in1 => \N__8580\,
            in2 => \N__8627\,
            in3 => \N__9563\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10230\,
            ce => \N__11218\,
            sr => \N__10696\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__8581\,
            in1 => \N__8438\,
            in2 => \N__8520\,
            in3 => \N__8603\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10230\,
            ce => \N__11218\,
            sr => \N__10696\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__8582\,
            in1 => \N__9677\,
            in2 => \N__8519\,
            in3 => \N__8465\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10230\,
            ce => \N__11218\,
            sr => \N__10696\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9655\,
            in1 => \N__10996\,
            in2 => \_gnd_net_\,
            in3 => \N__9065\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10793\,
            ce => \N__10766\,
            sr => \N__10689\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10982\,
            in1 => \N__8967\,
            in2 => \_gnd_net_\,
            in3 => \N__8927\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10764\,
            sr => \N__10681\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8968\,
            in1 => \N__10983\,
            in2 => \_gnd_net_\,
            in3 => \N__9022\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10764\,
            sr => \N__10681\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__9023\,
            in1 => \_gnd_net_\,
            in2 => \N__10998\,
            in3 => \N__9599\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10764\,
            sr => \N__10681\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__9062\,
            in1 => \_gnd_net_\,
            in2 => \N__10999\,
            in3 => \N__9656\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10764\,
            sr => \N__10681\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9708\,
            in1 => \N__10990\,
            in2 => \_gnd_net_\,
            in3 => \N__9063\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10764\,
            sr => \N__10681\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__9748\,
            in1 => \_gnd_net_\,
            in2 => \N__11000\,
            in3 => \N__9709\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10764\,
            sr => \N__10681\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8873\,
            in1 => \N__10994\,
            in2 => \_gnd_net_\,
            in3 => \N__9749\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10764\,
            sr => \N__10681\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__9009\,
            in1 => \_gnd_net_\,
            in2 => \N__8969\,
            in3 => \N__10980\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10790\,
            ce => \N__10762\,
            sr => \N__10674\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10846\,
            in1 => \N__10981\,
            in2 => \_gnd_net_\,
            in3 => \N__8872\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10790\,
            ce => \N__10762\,
            sr => \N__10674\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8853\,
            in1 => \N__10979\,
            in2 => \_gnd_net_\,
            in3 => \N__10845\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__10761\,
            sr => \N__10672\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__8729\,
            in1 => \N__10945\,
            in2 => \N__10847\,
            in3 => \N__8698\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            ce => 'H',
            sr => \N__10669\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__10070\,
            in1 => \N__11380\,
            in2 => \_gnd_net_\,
            in3 => \N__11470\,
            lcout => \U712_BYTE_ENABLE.N_409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9363\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10264\,
            ce => \N__9251\,
            sr => \N__10663\
        );

    \U712_BYTE_ENABLE.LLBE_0_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101010000"
        )
    port map (
            in0 => \N__11611\,
            in1 => \N__11547\,
            in2 => \N__11362\,
            in3 => \N__11440\,
            lcout => \LLBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CASn_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9227\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10234\,
            ce => 'H',
            sr => \N__10702\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10995\,
            in1 => \N__9710\,
            in2 => \_gnd_net_\,
            in3 => \N__9064\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10792\,
            ce => \N__10768\,
            sr => \N__10697\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9016\,
            in1 => \N__10936\,
            in2 => \_gnd_net_\,
            in3 => \N__9595\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10791\,
            ce => \N__10767\,
            sr => \N__10690\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8955\,
            in1 => \N__10935\,
            in2 => \_gnd_net_\,
            in3 => \N__8926\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10791\,
            ce => \N__10767\,
            sr => \N__10690\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9747\,
            in1 => \N__10938\,
            in2 => \_gnd_net_\,
            in3 => \N__8871\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10791\,
            ce => \N__10767\,
            sr => \N__10690\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9746\,
            in1 => \N__10937\,
            in2 => \_gnd_net_\,
            in3 => \N__9699\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10791\,
            ce => \N__10767\,
            sr => \N__10690\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10934\,
            in1 => \N__9651\,
            in2 => \_gnd_net_\,
            in3 => \N__9594\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__10765\,
            sr => \N__10682\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10933\,
            in1 => \N__9650\,
            in2 => \_gnd_net_\,
            in3 => \N__9593\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10789\,
            ce => \N__10763\,
            sr => \N__10675\
        );

    \U712_BYTE_ENABLE.N_146_i_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101010101"
        )
    port map (
            in0 => \N__9428\,
            in1 => \N__11089\,
            in2 => \N__9875\,
            in3 => \N__11172\,
            lcout => \N_146_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_RNI8MQ3_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9529\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110000"
        )
    port map (
            in0 => \N__11621\,
            in1 => \N__9422\,
            in2 => \N__10090\,
            in3 => \N__11549\,
            lcout => \U712_BYTE_ENABLE.N_406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_a2_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110000"
        )
    port map (
            in0 => \N__11620\,
            in1 => \N__9421\,
            in2 => \N__10089\,
            in3 => \N__11548\,
            lcout => \U712_BYTE_ENABLE.N_411\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11471\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11336\,
            lcout => \U712_BYTE_ENABLE.N_284_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_374_i_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111010000"
        )
    port map (
            in0 => \N__11613\,
            in1 => \N__11551\,
            in2 => \N__11463\,
            in3 => \N__11349\,
            lcout => \N_374_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_373_i_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011100000"
        )
    port map (
            in0 => \N__11612\,
            in1 => \N__11550\,
            in2 => \N__11462\,
            in3 => \N__11348\,
            lcout => \N_373_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UMBE_0_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010110000"
        )
    port map (
            in0 => \N__11614\,
            in1 => \N__11552\,
            in2 => \N__11464\,
            in3 => \N__11350\,
            lcout => \UMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__11270\,
            in1 => \N__11261\,
            in2 => \N__10079\,
            in3 => \N__10799\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10242\,
            ce => \N__11222\,
            sr => \N__10698\
        );

    \U712_BYTE_ENABLE.N_150_i_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110001"
        )
    port map (
            in0 => \N__11173\,
            in1 => \N__11099\,
            in2 => \N__9902\,
            in3 => \N__11088\,
            lcout => \N_150_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10309\,
            in1 => \N__10978\,
            in2 => \_gnd_net_\,
            in3 => \N__10832\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10788\,
            ce => \N__10769\,
            sr => \N__10699\
        );

    \U712_CHIP_RAM.RAS_SYNC_0_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__10470\,
            in1 => \N__10325\,
            in2 => \_gnd_net_\,
            in3 => \N__10313\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10260\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.N_136_i_LC_24_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000110000"
        )
    port map (
            in0 => \N__9858\,
            in1 => \N__10133\,
            in2 => \N__10094\,
            in3 => \N__11731\,
            lcout => \N_136_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001111111"
        )
    port map (
            in0 => \N__9857\,
            in1 => \N__9820\,
            in2 => \N__11743\,
            in3 => \N__11687\,
            lcout => \N_357\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

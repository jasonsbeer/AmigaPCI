-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 10 2025 20:32:12

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U400_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U400_TOP
entity U400_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    MA : out std_logic_vector(12 downto 0);
    A : in std_logic_vector(31 downto 0);
    LBENn : out std_logic;
    CS0n : out std_logic;
    UUBEn : out std_logic;
    TAn : out std_logic;
    CLK40 : in std_logic;
    RnW : in std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    WEn : out std_logic;
    LLBEn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    RASn : out std_logic;
    CS1n : out std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic);
end U400_TOP;

-- Architecture of U400_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U400_TOP is

signal \N__7251\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3353\ : std_logic;
signal \N__3350\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3306\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3254\ : std_logic;
signal \N__3251\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3102\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2904\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2862\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2854\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2747\ : std_logic;
signal \N__2744\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2737\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2705\ : std_logic;
signal \N__2702\ : std_logic;
signal \N__2699\ : std_logic;
signal \CLK40_ibuf_gb_io_gb_input\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \INVU400_SDRAM.REFRESH_COUNTER_1C_net\ : std_logic;
signal \A_c_21\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \A_c_22\ : std_logic;
signal \BANK1_c\ : std_logic;
signal \INVU400_SDRAM.BANK0C_net\ : std_logic;
signal \INVU400_SDRAM.CS1_ENC_net\ : std_logic;
signal \U400_SDRAM.un1_SDRAM_COUNTER59_0\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_5_sqmuxa\ : std_logic;
signal \INVU400_SDRAM.RAM_CYCLEC_net\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_0\ : std_logic;
signal \bfn_2_4_0_\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_1\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_2\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_3\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_4\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_5\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_6\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_7\ : std_logic;
signal \INVU400_SDRAM.REFRESH_COUNTER_2C_net\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_RNIV59H2Z0Z_1\ : std_logic;
signal \INVU400_SDRAM.CS0_ENC_net\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_8\ : std_logic;
signal \U400_SDRAM.un1_REFRESH_COUNTERlt7_0_cascade_\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U400_SDRAM.N_337_1_cascade_\ : std_logic;
signal \U400_SDRAM.N_64_cascade_\ : std_logic;
signal \U400_SDRAM.CS1_EN_0\ : std_logic;
signal \U400_SDRAM.N_64\ : std_logic;
signal \U400_SDRAM.N_72_cascade_\ : std_logic;
signal \U400_SDRAM.N_40\ : std_logic;
signal \A_c_23\ : std_logic;
signal \U400_SDRAM.N_40_cascade_\ : std_logic;
signal \U400_SDRAM.CS0_EN_0\ : std_logic;
signal \U400_SDRAM.N_115\ : std_logic;
signal \U400_SDRAM.RAM_CYCLEZ0\ : std_logic;
signal \U400_SDRAM.CS1_ENZ0\ : std_logic;
signal \CS1n_c\ : std_logic;
signal \CASn_c\ : std_logic;
signal \WEn_c\ : std_logic;
signal \INVU400_SDRAM.CS1nC_net\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U400_SDRAM.CS0_ENZ0\ : std_logic;
signal \CS0n_c\ : std_logic;
signal \INVU400_SDRAM.RASnC_net\ : std_logic;
signal \A_c_31\ : std_logic;
signal \A_c_30\ : std_logic;
signal \A_c_29\ : std_logic;
signal \A_c_28\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U400_SDRAM.N_101\ : std_logic;
signal \U400_ADDRESS_DECODE_RAM_SPACE_i_o3_2\ : std_logic;
signal \A_c_27\ : std_logic;
signal \U400_ADDRESS_DECODE_RAM_SPACE_i_o3_1\ : std_logic;
signal \INVU400_SDRAM.SDRAM_COUNTER_1C_net\ : std_logic;
signal \INVU400_SDRAM.SDRAM_CONFIGUREDC_net\ : std_logic;
signal \U400_SDRAM.N_113_cascade_\ : std_logic;
signal \U400_SDRAM.N_39_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_1_sqmuxa_i_0_1\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_a2_1_0_0\ : std_logic;
signal \U400_SDRAM.N_78_cascade_\ : std_logic;
signal \U400_SDRAM.N_337_1\ : std_logic;
signal \U400_SDRAM.N_12_cascade_\ : std_logic;
signal \U400_SDRAM.N_91_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_0_103_i_i_a3_0_0\ : std_logic;
signal \U400_SDRAM.N_89\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_0_103_i_i_0_cascade_\ : std_logic;
signal \INVU400_SDRAM.SDRAM_CMD_1C_net\ : std_logic;
signal \A_c_8\ : std_logic;
signal \A_c_19\ : std_logic;
signal \MA_c_6\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_17\ : std_logic;
signal \MA_c_4\ : std_logic;
signal \A_c_20\ : std_logic;
signal \A_c_9\ : std_logic;
signal \MA_c_7\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_6C_net\ : std_logic;
signal \U400_SDRAM.RAM_CYCLE_STARTZ0\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_4_sqmuxa_0_a3_0\ : std_logic;
signal \RnW_c\ : std_logic;
signal \INVU400_SDRAM.TACKC_net\ : std_logic;
signal \U400_SDRAM.N_113\ : std_logic;
signal \U400_SDRAM.N_63\ : std_logic;
signal \U400_SDRAM.N_20_cascade_\ : std_logic;
signal \U400_SDRAM.N_35\ : std_logic;
signal \U400_SDRAM.N_39\ : std_logic;
signal \U400_SDRAM.N_35_cascade_\ : std_logic;
signal \U400_SDRAM.N_44_cascade_\ : std_logic;
signal \U400_SDRAM.N_108\ : std_logic;
signal \U400_SDRAM.N_108_cascade_\ : std_logic;
signal \U400_SDRAM.N_109\ : std_logic;
signal \U400_SDRAM.N_52\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \U400_SDRAM.N_86\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_1_0_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_3_sqmuxa\ : std_logic;
signal \U400_SDRAM.N_118\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_3_sqmuxa_0_a3_0_a2_0\ : std_logic;
signal \INVU400_SDRAM.SDRAM_COUNTER_0C_net\ : std_logic;
signal \U400_SDRAM.N_46_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_a2_0_0_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_1_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_3\ : std_logic;
signal \U400_SDRAM.N_60\ : std_logic;
signal \U400_SDRAM.N_97_cascade_\ : std_logic;
signal \U400_SDRAM.N_20\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_1_66_i_0_2_cascade_\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U400_SDRAM.N_11\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_1\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_3_cascade_\ : std_logic;
signal \U400_SDRAM.N_38\ : std_logic;
signal \INVU400_SDRAM.SDRAM_CMD_0C_net\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_a2_2_0_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_2\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_16\ : std_logic;
signal \MA_c_3\ : std_logic;
signal \A_c_26\ : std_logic;
signal \MA_c_12\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U400_SDRAM.MA_5_iv_0_5\ : std_logic;
signal \MA_c_5\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_3C_net\ : std_logic;
signal \U400_SDRAM.N_8_cascade_\ : std_logic;
signal \U400_SDRAM.un1_SDRAM_COUNTER59_4_i_1\ : std_logic;
signal \U400_SDRAM.N_15_cascade_\ : std_logic;
signal \U400_SDRAM.N_87\ : std_logic;
signal \U400_SDRAM.N_25\ : std_logic;
signal \U400_SDRAM.N_84\ : std_logic;
signal \U400_SDRAM.N_88\ : std_logic;
signal \U400_SDRAM.N_48\ : std_logic;
signal \bfn_6_6_0_\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_s_1\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_s_3\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U400_SDRAM.N_29\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \INVU400_SDRAM.SDRAM_COUNTER_2C_net\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U400_SDRAM.N_336_1\ : std_logic;
signal \U400_SDRAM.N_56_cascade_\ : std_logic;
signal \U400_SDRAM.TACK_7_iv_i_0\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U400_SDRAM.N_28\ : std_logic;
signal \U400_SDRAM.N_110\ : std_logic;
signal \U400_SDRAM.WRITE_CYCLEZ0\ : std_logic;
signal \U400_SDRAM.N_13\ : std_logic;
signal \U400_SDRAM.N_44\ : std_logic;
signal \U400_SDRAM.N_8\ : std_logic;
signal \U400_SDRAM.N_13_cascade_\ : std_logic;
signal \U400_SDRAM.N_76\ : std_logic;
signal \U400_SDRAM.un1_SDRAM_COUNTER59_1_1_0\ : std_logic;
signal \U400_SDRAM.N_46\ : std_logic;
signal \U400_SDRAM.N_33_cascade_\ : std_logic;
signal \U400_SDRAM.N_67\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_1_66_i_0_1\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U400_SDRAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U400_SDRAM.N_30\ : std_logic;
signal \U400_SDRAM.TA_COUNTER_srsts_0_a4_0_0\ : std_logic;
signal \U400_SDRAM.N_243_0\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U400_SDRAM.TA_COUNTERZ0Z_0\ : std_logic;
signal \U400_SDRAM.N_243_0_cascade_\ : std_logic;
signal \U400_SDRAM.TACKZ0\ : std_logic;
signal \U400_SDRAM.N_241_0_en\ : std_logic;
signal \U400_SDRAM.un1_TA_COUNTER_6_0_0\ : std_logic;
signal \U400_SDRAM.N_244_0\ : std_logic;
signal \TA_OUT\ : std_logic;
signal \N_53\ : std_logic;
signal \U400_SDRAM.TA_COUNTERZ0Z_1\ : std_logic;
signal \U400_SDRAM.TA_OUT_5_0\ : std_logic;
signal \A_c_24\ : std_logic;
signal \MA_c_11\ : std_logic;
signal \A_c_11\ : std_logic;
signal \MA_c_9\ : std_logic;
signal \A_c_25\ : std_logic;
signal \A_c_10\ : std_logic;
signal \MA_c_8\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_11C_net\ : std_logic;
signal \U400_SDRAM.TA_COUNTERZ0Z_4\ : std_logic;
signal \U400_SDRAM.TA_COUNTERZ0Z_5\ : std_logic;
signal \U400_SDRAM.TA_COUNTERZ0Z_2\ : std_logic;
signal \U400_SDRAM.TA_COUNTERZ0Z_3\ : std_logic;
signal \CLK40_c_g\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_1_sqmuxa_1\ : std_logic;
signal \U400_SDRAM.BURSTZ0\ : std_logic;
signal \INVU400_SDRAM.BURSTC_net\ : std_logic;
signal \A_c_12\ : std_logic;
signal \MA_c_10\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_13\ : std_logic;
signal \MA_c_0\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_10C_net\ : std_logic;
signal \N_51\ : std_logic;
signal \N_47\ : std_logic;
signal \TA_EN_i\ : std_logic;
signal \N_542_i\ : std_logic;
signal \U400_BYTE_ENABLE.N_71\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \U400_BYTE_ENABLE.N_54_i\ : std_logic;
signal \A_c_0\ : std_logic;
signal \RAM_SPACE_i_o3dup\ : std_logic;
signal \U400_BYTE_ENABLE.N_54_i_cascade_\ : std_logic;
signal \A_c_1\ : std_logic;
signal \N_49\ : std_logic;
signal \U400_SDRAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U400_SDRAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U400_SDRAM.MA_5_iv_0_1\ : std_logic;
signal \MA_c_1\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U400_SDRAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U400_SDRAM.MA20\ : std_logic;
signal \MA_c_2\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_1C_net\ : std_logic;
signal \U400_SDRAM.un1_MA21_0_i_0\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;

signal \MA_wire\ : std_logic_vector(12 downto 0);
signal \A_wire\ : std_logic_vector(31 downto 0);
signal \CASn_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \UUBEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \LLBEn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \TAn_wire\ : std_logic;
signal \LBENn_wire\ : std_logic;
signal \CS1n_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CS0n_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CLK40_wire\ : std_logic;

begin
    MA <= \MA_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    BANK1 <= \BANK1_wire\;
    UUBEn <= \UUBEn_wire\;
    \SIZ_wire\ <= SIZ;
    LLBEn <= \LLBEn_wire\;
    \TSn_wire\ <= TSn;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    \RESETn_wire\ <= RESETn;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    TAn <= \TAn_wire\;
    LBENn <= \LBENn_wire\;
    CS1n <= \CS1n_wire\;
    WEn <= \WEn_wire\;
    \RnW_wire\ <= RnW;
    CS0n <= \CS0n_wire\;
    LMBEn <= \LMBEn_wire\;
    \CLK40_wire\ <= CLK40;

    \MA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7251\,
            DIN => \N__7250\,
            DOUT => \N__7249\,
            PACKAGEPIN => \MA_wire\(7)
        );

    \MA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7251\,
            PADOUT => \N__7250\,
            PADIN => \N__7249\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3371\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7242\,
            DIN => \N__7241\,
            DOUT => \N__7240\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7242\,
            PADOUT => \N__7241\,
            PADIN => \N__7240\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7233\,
            DIN => \N__7232\,
            DOUT => \N__7231\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7233\,
            PADOUT => \N__7232\,
            PADIN => \N__7231\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3038\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7224\,
            DIN => \N__7223\,
            DOUT => \N__7222\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7224\,
            PADOUT => \N__7223\,
            PADIN => \N__7222\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2753\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7215\,
            DIN => \N__7214\,
            DOUT => \N__7213\,
            PACKAGEPIN => \MA_wire\(8)
        );

    \MA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7215\,
            PADOUT => \N__7214\,
            PADIN => \N__7213\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5564\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7206\,
            DIN => \N__7205\,
            DOUT => \N__7204\,
            PACKAGEPIN => \MA_wire\(10)
        );

    \MA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7206\,
            PADOUT => \N__7205\,
            PADIN => \N__7204\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6284\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7197\,
            DIN => \N__7196\,
            DOUT => \N__7195\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7197\,
            PADOUT => \N__7196\,
            PADIN => \N__7195\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7188\,
            DIN => \N__7187\,
            DOUT => \N__7186\,
            PACKAGEPIN => \MA_wire\(2)
        );

    \MA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7188\,
            PADOUT => \N__7187\,
            PADIN => \N__7186\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6428\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7179\,
            DIN => \N__7178\,
            DOUT => \N__7177\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7179\,
            PADOUT => \N__7178\,
            PADIN => \N__7177\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7170\,
            DIN => \N__7169\,
            DOUT => \N__7168\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7170\,
            PADOUT => \N__7169\,
            PADIN => \N__7168\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7161\,
            DIN => \N__7160\,
            DOUT => \N__7159\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7161\,
            PADOUT => \N__7160\,
            PADIN => \N__7159\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5093\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7152\,
            DIN => \N__7151\,
            DOUT => \N__7150\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7152\,
            PADOUT => \N__7151\,
            PADIN => \N__7150\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7143\,
            DIN => \N__7142\,
            DOUT => \N__7141\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7143\,
            PADOUT => \N__7142\,
            PADIN => \N__7141\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7134\,
            DIN => \N__7133\,
            DOUT => \N__7132\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7134\,
            PADOUT => \N__7133\,
            PADIN => \N__7132\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7125\,
            DIN => \N__7124\,
            DOUT => \N__7123\,
            PACKAGEPIN => \MA_wire\(12)
        );

    \MA_obuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7125\,
            PADOUT => \N__7124\,
            PADIN => \N__7123\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3932\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7116\,
            DIN => \N__7115\,
            DOUT => \N__7114\,
            PACKAGEPIN => \MA_wire\(1)
        );

    \MA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7116\,
            PADOUT => \N__7115\,
            PADIN => \N__7114\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6638\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7107\,
            DIN => \N__7106\,
            DOUT => \N__7105\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7107\,
            PADOUT => \N__7106\,
            PADIN => \N__7105\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7098\,
            DIN => \N__7097\,
            DOUT => \N__7096\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7098\,
            PADOUT => \N__7097\,
            PADIN => \N__7096\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7089\,
            DIN => \N__7088\,
            DOUT => \N__7087\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7089\,
            PADOUT => \N__7088\,
            PADIN => \N__7087\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7080\,
            DIN => \N__7079\,
            DOUT => \N__7078\,
            PACKAGEPIN => \MA_wire\(4)
        );

    \MA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7080\,
            PADOUT => \N__7079\,
            PADIN => \N__7078\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3416\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7071\,
            DIN => \N__7070\,
            DOUT => \N__7069\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7071\,
            PADOUT => \N__7070\,
            PADIN => \N__7069\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7062\,
            DIN => \N__7061\,
            DOUT => \N__7060\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7062\,
            PADOUT => \N__7061\,
            PADIN => \N__7060\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7053\,
            DIN => \N__7052\,
            DOUT => \N__7051\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7053\,
            PADOUT => \N__7052\,
            PADIN => \N__7051\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6236\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7044\,
            DIN => \N__7043\,
            DOUT => \N__7042\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7044\,
            PADOUT => \N__7043\,
            PADIN => \N__7042\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7035\,
            DIN => \N__7034\,
            DOUT => \N__7033\,
            PACKAGEPIN => \MA_wire\(9)
        );

    \MA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7035\,
            PADOUT => \N__7034\,
            PADIN => \N__7033\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5600\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7026\,
            DIN => \N__7025\,
            DOUT => \N__7024\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7026\,
            PADOUT => \N__7025\,
            PADIN => \N__7024\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6245\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7017\,
            DIN => \N__7016\,
            DOUT => \N__7015\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7017\,
            PADOUT => \N__7016\,
            PADIN => \N__7015\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7008\,
            DIN => \N__7007\,
            DOUT => \N__7006\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7008\,
            PADOUT => \N__7007\,
            PADIN => \N__7006\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6999\,
            DIN => \N__6998\,
            DOUT => \N__6997\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6999\,
            PADOUT => \N__6998\,
            PADIN => \N__6997\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2792\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6990\,
            DIN => \N__6989\,
            DOUT => \N__6988\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6990\,
            PADOUT => \N__6989\,
            PADIN => \N__6988\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6981\,
            DIN => \N__6980\,
            DOUT => \N__6979\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6981\,
            PADOUT => \N__6980\,
            PADIN => \N__6979\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6972\,
            DIN => \N__6971\,
            DOUT => \N__6970\,
            PACKAGEPIN => \MA_wire\(3)
        );

    \MA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6972\,
            PADOUT => \N__6971\,
            PADIN => \N__6970\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3965\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6963\,
            DIN => \N__6962\,
            DOUT => \N__6961\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6963\,
            PADOUT => \N__6962\,
            PADIN => \N__6961\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6954\,
            DIN => \N__6953\,
            DOUT => \N__6952\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6954\,
            PADOUT => \N__6953\,
            PADIN => \N__6952\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6945\,
            DIN => \N__6944\,
            DOUT => \N__6943\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6945\,
            PADOUT => \N__6944\,
            PADIN => \N__6943\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6936\,
            DIN => \N__6935\,
            DOUT => \N__6934\,
            PACKAGEPIN => \MA_wire\(6)
        );

    \MA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6936\,
            PADOUT => \N__6935\,
            PADIN => \N__6934\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3449\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6927\,
            DIN => \N__6926\,
            DOUT => \N__6925\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6927\,
            PADOUT => \N__6926\,
            PADIN => \N__6925\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6918\,
            DIN => \N__6917\,
            DOUT => \N__6916\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6918\,
            PADOUT => \N__6917\,
            PADIN => \N__6916\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6909\,
            DIN => \N__6908\,
            DOUT => \N__6907\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6909\,
            PADOUT => \N__6908\,
            PADIN => \N__6907\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6900\,
            DIN => \N__6899\,
            DOUT => \N__6898\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6900\,
            PADOUT => \N__6899\,
            PADIN => \N__6898\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3299\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6891\,
            DIN => \N__6890\,
            DOUT => \N__6889\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6891\,
            PADOUT => \N__6890\,
            PADIN => \N__6889\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6882\,
            DIN => \N__6881\,
            DOUT => \N__6880\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6882\,
            PADOUT => \N__6881\,
            PADIN => \N__6880\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2816\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6873\,
            DIN => \N__6872\,
            DOUT => \N__6871\,
            PACKAGEPIN => \MA_wire\(11)
        );

    \MA_obuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6873\,
            PADOUT => \N__6872\,
            PADIN => \N__6871\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5618\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TAn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6864\,
            DIN => \N__6863\,
            DOUT => \N__6862\,
            PACKAGEPIN => \TAn_wire\
        );

    \TAn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__6864\,
            PADOUT => \N__6863\,
            PADIN => \N__6862\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6212\,
            DIN0 => OPEN,
            DOUT0 => \N__5111\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6855\,
            DIN => \N__6854\,
            DOUT => \N__6853\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6855\,
            PADOUT => \N__6854\,
            PADIN => \N__6853\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6846\,
            DIN => \N__6845\,
            DOUT => \N__6844\,
            PACKAGEPIN => \MA_wire\(5)
        );

    \MA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6846\,
            PADOUT => \N__6845\,
            PADIN => \N__6844\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3896\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6837\,
            DIN => \N__6836\,
            DOUT => \N__6835\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6837\,
            PADOUT => \N__6836\,
            PADIN => \N__6835\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6828\,
            DIN => \N__6827\,
            DOUT => \N__6826\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6828\,
            PADOUT => \N__6827\,
            PADIN => \N__6826\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LBENn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6819\,
            DIN => \N__6818\,
            DOUT => \N__6817\,
            PACKAGEPIN => \LBENn_wire\
        );

    \LBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6819\,
            PADOUT => \N__6818\,
            PADIN => \N__6817\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5984\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6810\,
            DIN => \N__6809\,
            DOUT => \N__6808\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6810\,
            PADOUT => \N__6809\,
            PADIN => \N__6808\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CS1n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6801\,
            DIN => \N__6800\,
            DOUT => \N__6799\,
            PACKAGEPIN => \CS1n_wire\
        );

    \CS1n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6801\,
            PADOUT => \N__6800\,
            PADIN => \N__6799\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3053\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6792\,
            DIN => \N__6791\,
            DOUT => \N__6790\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6792\,
            PADOUT => \N__6791\,
            PADIN => \N__6790\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6783\,
            DIN => \N__6782\,
            DOUT => \N__6781\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6783\,
            PADOUT => \N__6782\,
            PADIN => \N__6781\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6774\,
            DIN => \N__6773\,
            DOUT => \N__6772\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6774\,
            PADOUT => \N__6773\,
            PADIN => \N__6772\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6765\,
            DIN => \N__6764\,
            DOUT => \N__6763\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6765\,
            PADOUT => \N__6764\,
            PADIN => \N__6763\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6756\,
            DIN => \N__6755\,
            DOUT => \N__6754\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6756\,
            PADOUT => \N__6755\,
            PADIN => \N__6754\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3029\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6747\,
            DIN => \N__6746\,
            DOUT => \N__6745\,
            PACKAGEPIN => \MA_wire\(0)
        );

    \MA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6747\,
            PADOUT => \N__6746\,
            PADIN => \N__6745\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6251\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6738\,
            DIN => \N__6737\,
            DOUT => \N__6736\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6738\,
            PADOUT => \N__6737\,
            PADIN => \N__6736\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6729\,
            DIN => \N__6728\,
            DOUT => \N__6727\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6729\,
            PADOUT => \N__6728\,
            PADIN => \N__6727\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6720\,
            DIN => \N__6719\,
            DOUT => \N__6718\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6720\,
            PADOUT => \N__6719\,
            PADIN => \N__6718\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CS0n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6711\,
            DIN => \N__6710\,
            DOUT => \N__6709\,
            PACKAGEPIN => \CS0n_wire\
        );

    \CS0n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6711\,
            PADOUT => \N__6710\,
            PADIN => \N__6709\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3272\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6702\,
            DIN => \N__6701\,
            DOUT => \N__6700\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6702\,
            PADOUT => \N__6701\,
            PADIN => \N__6700\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6693\,
            DIN => \N__6692\,
            DOUT => \N__6691\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6693\,
            PADOUT => \N__6692\,
            PADIN => \N__6691\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5891\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6684\,
            DIN => \N__6683\,
            DOUT => \N__6682\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6684\,
            PADOUT => \N__6683\,
            PADIN => \N__6682\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6675\,
            DIN => \N__6674\,
            DOUT => \N__6673\,
            PACKAGEPIN => \CLK40_wire\
        );

    \CLK40_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6675\,
            PADOUT => \N__6674\,
            PADIN => \N__6673\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_ibuf_gb_io_gb_input\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1565\ : InMux
    port map (
            O => \N__6656\,
            I => \N__6653\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__6653\,
            I => \N__6650\
        );

    \I__1563\ : Span4Mux_h
    port map (
            O => \N__6650\,
            I => \N__6647\
        );

    \I__1562\ : Odrv4
    port map (
            O => \N__6647\,
            I => \A_c_3\
        );

    \I__1561\ : InMux
    port map (
            O => \N__6644\,
            I => \N__6641\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__6641\,
            I => \U400_SDRAM.MA_5_iv_0_1\
        );

    \I__1559\ : IoInMux
    port map (
            O => \N__6638\,
            I => \N__6635\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__6635\,
            I => \MA_c_1\
        );

    \I__1557\ : InMux
    port map (
            O => \N__6632\,
            I => \N__6629\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__6629\,
            I => \N__6626\
        );

    \I__1555\ : Span4Mux_s2_v
    port map (
            O => \N__6626\,
            I => \N__6623\
        );

    \I__1554\ : IoSpan4Mux
    port map (
            O => \N__6623\,
            I => \N__6620\
        );

    \I__1553\ : Odrv4
    port map (
            O => \N__6620\,
            I => \A_c_4\
        );

    \I__1552\ : InMux
    port map (
            O => \N__6617\,
            I => \N__6609\
        );

    \I__1551\ : InMux
    port map (
            O => \N__6616\,
            I => \N__6604\
        );

    \I__1550\ : InMux
    port map (
            O => \N__6615\,
            I => \N__6604\
        );

    \I__1549\ : InMux
    port map (
            O => \N__6614\,
            I => \N__6597\
        );

    \I__1548\ : InMux
    port map (
            O => \N__6613\,
            I => \N__6597\
        );

    \I__1547\ : InMux
    port map (
            O => \N__6612\,
            I => \N__6597\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__6609\,
            I => \N__6585\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__6604\,
            I => \N__6585\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__6597\,
            I => \N__6582\
        );

    \I__1543\ : InMux
    port map (
            O => \N__6596\,
            I => \N__6579\
        );

    \I__1542\ : InMux
    port map (
            O => \N__6595\,
            I => \N__6571\
        );

    \I__1541\ : InMux
    port map (
            O => \N__6594\,
            I => \N__6571\
        );

    \I__1540\ : InMux
    port map (
            O => \N__6593\,
            I => \N__6568\
        );

    \I__1539\ : InMux
    port map (
            O => \N__6592\,
            I => \N__6565\
        );

    \I__1538\ : InMux
    port map (
            O => \N__6591\,
            I => \N__6560\
        );

    \I__1537\ : InMux
    port map (
            O => \N__6590\,
            I => \N__6560\
        );

    \I__1536\ : Span4Mux_s1_v
    port map (
            O => \N__6585\,
            I => \N__6553\
        );

    \I__1535\ : Span4Mux_h
    port map (
            O => \N__6582\,
            I => \N__6553\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__6579\,
            I => \N__6553\
        );

    \I__1533\ : CascadeMux
    port map (
            O => \N__6578\,
            I => \N__6550\
        );

    \I__1532\ : InMux
    port map (
            O => \N__6577\,
            I => \N__6544\
        );

    \I__1531\ : InMux
    port map (
            O => \N__6576\,
            I => \N__6544\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__6571\,
            I => \N__6539\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__6568\,
            I => \N__6539\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__6565\,
            I => \N__6533\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__6560\,
            I => \N__6533\
        );

    \I__1526\ : Span4Mux_v
    port map (
            O => \N__6553\,
            I => \N__6530\
        );

    \I__1525\ : InMux
    port map (
            O => \N__6550\,
            I => \N__6524\
        );

    \I__1524\ : InMux
    port map (
            O => \N__6549\,
            I => \N__6524\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__6544\,
            I => \N__6521\
        );

    \I__1522\ : Span4Mux_v
    port map (
            O => \N__6539\,
            I => \N__6518\
        );

    \I__1521\ : InMux
    port map (
            O => \N__6538\,
            I => \N__6515\
        );

    \I__1520\ : Span4Mux_v
    port map (
            O => \N__6533\,
            I => \N__6510\
        );

    \I__1519\ : Span4Mux_h
    port map (
            O => \N__6530\,
            I => \N__6510\
        );

    \I__1518\ : InMux
    port map (
            O => \N__6529\,
            I => \N__6507\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__6524\,
            I => \N__6502\
        );

    \I__1516\ : Span12Mux_s3_v
    port map (
            O => \N__6521\,
            I => \N__6502\
        );

    \I__1515\ : Odrv4
    port map (
            O => \N__6518\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__6515\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1513\ : Odrv4
    port map (
            O => \N__6510\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__6507\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1511\ : Odrv12
    port map (
            O => \N__6502\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1510\ : CascadeMux
    port map (
            O => \N__6491\,
            I => \N__6488\
        );

    \I__1509\ : InMux
    port map (
            O => \N__6488\,
            I => \N__6485\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__6485\,
            I => \A_c_15\
        );

    \I__1507\ : InMux
    port map (
            O => \N__6482\,
            I => \N__6476\
        );

    \I__1506\ : InMux
    port map (
            O => \N__6481\,
            I => \N__6473\
        );

    \I__1505\ : InMux
    port map (
            O => \N__6480\,
            I => \N__6468\
        );

    \I__1504\ : InMux
    port map (
            O => \N__6479\,
            I => \N__6468\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__6476\,
            I => \N__6463\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__6473\,
            I => \N__6463\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__6468\,
            I => \N__6457\
        );

    \I__1500\ : Span4Mux_s2_v
    port map (
            O => \N__6463\,
            I => \N__6452\
        );

    \I__1499\ : InMux
    port map (
            O => \N__6462\,
            I => \N__6445\
        );

    \I__1498\ : InMux
    port map (
            O => \N__6461\,
            I => \N__6445\
        );

    \I__1497\ : InMux
    port map (
            O => \N__6460\,
            I => \N__6445\
        );

    \I__1496\ : Span4Mux_s2_v
    port map (
            O => \N__6457\,
            I => \N__6442\
        );

    \I__1495\ : InMux
    port map (
            O => \N__6456\,
            I => \N__6437\
        );

    \I__1494\ : InMux
    port map (
            O => \N__6455\,
            I => \N__6437\
        );

    \I__1493\ : Odrv4
    port map (
            O => \N__6452\,
            I => \U400_SDRAM.MA20\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__6445\,
            I => \U400_SDRAM.MA20\
        );

    \I__1491\ : Odrv4
    port map (
            O => \N__6442\,
            I => \U400_SDRAM.MA20\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__6437\,
            I => \U400_SDRAM.MA20\
        );

    \I__1489\ : IoInMux
    port map (
            O => \N__6428\,
            I => \N__6425\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__6425\,
            I => \MA_c_2\
        );

    \I__1487\ : CEMux
    port map (
            O => \N__6422\,
            I => \N__6415\
        );

    \I__1486\ : CEMux
    port map (
            O => \N__6421\,
            I => \N__6412\
        );

    \I__1485\ : CEMux
    port map (
            O => \N__6420\,
            I => \N__6409\
        );

    \I__1484\ : CEMux
    port map (
            O => \N__6419\,
            I => \N__6406\
        );

    \I__1483\ : CEMux
    port map (
            O => \N__6418\,
            I => \N__6403\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__6415\,
            I => \N__6400\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__6412\,
            I => \N__6397\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__6409\,
            I => \N__6392\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__6406\,
            I => \N__6392\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__6403\,
            I => \N__6389\
        );

    \I__1477\ : Span4Mux_h
    port map (
            O => \N__6400\,
            I => \N__6386\
        );

    \I__1476\ : Span4Mux_v
    port map (
            O => \N__6397\,
            I => \N__6383\
        );

    \I__1475\ : Span4Mux_s2_v
    port map (
            O => \N__6392\,
            I => \N__6378\
        );

    \I__1474\ : Span4Mux_v
    port map (
            O => \N__6389\,
            I => \N__6378\
        );

    \I__1473\ : Odrv4
    port map (
            O => \N__6386\,
            I => \U400_SDRAM.un1_MA21_0_i_0\
        );

    \I__1472\ : Odrv4
    port map (
            O => \N__6383\,
            I => \U400_SDRAM.un1_MA21_0_i_0\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__6378\,
            I => \U400_SDRAM.un1_MA21_0_i_0\
        );

    \I__1470\ : CascadeMux
    port map (
            O => \N__6371\,
            I => \N__6368\
        );

    \I__1469\ : InMux
    port map (
            O => \N__6368\,
            I => \N__6365\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__6365\,
            I => \N__6359\
        );

    \I__1467\ : SRMux
    port map (
            O => \N__6364\,
            I => \N__6305\
        );

    \I__1466\ : SRMux
    port map (
            O => \N__6363\,
            I => \N__6305\
        );

    \I__1465\ : SRMux
    port map (
            O => \N__6362\,
            I => \N__6305\
        );

    \I__1464\ : Glb2LocalMux
    port map (
            O => \N__6359\,
            I => \N__6305\
        );

    \I__1463\ : SRMux
    port map (
            O => \N__6358\,
            I => \N__6305\
        );

    \I__1462\ : SRMux
    port map (
            O => \N__6357\,
            I => \N__6305\
        );

    \I__1461\ : SRMux
    port map (
            O => \N__6356\,
            I => \N__6305\
        );

    \I__1460\ : SRMux
    port map (
            O => \N__6355\,
            I => \N__6305\
        );

    \I__1459\ : SRMux
    port map (
            O => \N__6354\,
            I => \N__6305\
        );

    \I__1458\ : SRMux
    port map (
            O => \N__6353\,
            I => \N__6305\
        );

    \I__1457\ : SRMux
    port map (
            O => \N__6352\,
            I => \N__6305\
        );

    \I__1456\ : SRMux
    port map (
            O => \N__6351\,
            I => \N__6305\
        );

    \I__1455\ : SRMux
    port map (
            O => \N__6350\,
            I => \N__6305\
        );

    \I__1454\ : SRMux
    port map (
            O => \N__6349\,
            I => \N__6305\
        );

    \I__1453\ : SRMux
    port map (
            O => \N__6348\,
            I => \N__6305\
        );

    \I__1452\ : SRMux
    port map (
            O => \N__6347\,
            I => \N__6305\
        );

    \I__1451\ : SRMux
    port map (
            O => \N__6346\,
            I => \N__6305\
        );

    \I__1450\ : SRMux
    port map (
            O => \N__6345\,
            I => \N__6305\
        );

    \I__1449\ : SRMux
    port map (
            O => \N__6344\,
            I => \N__6305\
        );

    \I__1448\ : GlobalMux
    port map (
            O => \N__6305\,
            I => \N__6302\
        );

    \I__1447\ : gio2CtrlBuf
    port map (
            O => \N__6302\,
            I => \RESETn_c_i_g\
        );

    \I__1446\ : CascadeMux
    port map (
            O => \N__6299\,
            I => \N__6296\
        );

    \I__1445\ : InMux
    port map (
            O => \N__6296\,
            I => \N__6293\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__6293\,
            I => \N__6290\
        );

    \I__1443\ : Span4Mux_h
    port map (
            O => \N__6290\,
            I => \N__6287\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__6287\,
            I => \A_c_12\
        );

    \I__1441\ : IoInMux
    port map (
            O => \N__6284\,
            I => \N__6281\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__6281\,
            I => \MA_c_10\
        );

    \I__1439\ : InMux
    port map (
            O => \N__6278\,
            I => \N__6275\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__6275\,
            I => \N__6272\
        );

    \I__1437\ : Span4Mux_h
    port map (
            O => \N__6272\,
            I => \N__6269\
        );

    \I__1436\ : Odrv4
    port map (
            O => \N__6269\,
            I => \A_c_2\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__6266\,
            I => \N__6263\
        );

    \I__1434\ : InMux
    port map (
            O => \N__6263\,
            I => \N__6260\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__6260\,
            I => \N__6257\
        );

    \I__1432\ : Span12Mux_s5_v
    port map (
            O => \N__6257\,
            I => \N__6254\
        );

    \I__1431\ : Odrv12
    port map (
            O => \N__6254\,
            I => \A_c_13\
        );

    \I__1430\ : IoInMux
    port map (
            O => \N__6251\,
            I => \N__6248\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__6248\,
            I => \MA_c_0\
        );

    \I__1428\ : IoInMux
    port map (
            O => \N__6245\,
            I => \N__6242\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__6242\,
            I => \N__6239\
        );

    \I__1426\ : Odrv4
    port map (
            O => \N__6239\,
            I => \N_51\
        );

    \I__1425\ : IoInMux
    port map (
            O => \N__6236\,
            I => \N__6233\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__6233\,
            I => \N__6230\
        );

    \I__1423\ : Odrv4
    port map (
            O => \N__6230\,
            I => \N_47\
        );

    \I__1422\ : InMux
    port map (
            O => \N__6227\,
            I => \N__6224\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__6224\,
            I => \N__6220\
        );

    \I__1420\ : InMux
    port map (
            O => \N__6223\,
            I => \N__6217\
        );

    \I__1419\ : Odrv4
    port map (
            O => \N__6220\,
            I => \TA_EN_i\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__6217\,
            I => \TA_EN_i\
        );

    \I__1417\ : IoInMux
    port map (
            O => \N__6212\,
            I => \N__6209\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__6209\,
            I => \N__6206\
        );

    \I__1415\ : IoSpan4Mux
    port map (
            O => \N__6206\,
            I => \N__6203\
        );

    \I__1414\ : Odrv4
    port map (
            O => \N__6203\,
            I => \N_542_i\
        );

    \I__1413\ : InMux
    port map (
            O => \N__6200\,
            I => \N__6194\
        );

    \I__1412\ : InMux
    port map (
            O => \N__6199\,
            I => \N__6194\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__6194\,
            I => \U400_BYTE_ENABLE.N_71\
        );

    \I__1410\ : InMux
    port map (
            O => \N__6191\,
            I => \N__6187\
        );

    \I__1409\ : InMux
    port map (
            O => \N__6190\,
            I => \N__6182\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__6187\,
            I => \N__6179\
        );

    \I__1407\ : InMux
    port map (
            O => \N__6186\,
            I => \N__6174\
        );

    \I__1406\ : InMux
    port map (
            O => \N__6185\,
            I => \N__6174\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__6182\,
            I => \N__6167\
        );

    \I__1404\ : Span4Mux_h
    port map (
            O => \N__6179\,
            I => \N__6162\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__6174\,
            I => \N__6162\
        );

    \I__1402\ : InMux
    port map (
            O => \N__6173\,
            I => \N__6159\
        );

    \I__1401\ : InMux
    port map (
            O => \N__6172\,
            I => \N__6156\
        );

    \I__1400\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6153\
        );

    \I__1399\ : InMux
    port map (
            O => \N__6170\,
            I => \N__6150\
        );

    \I__1398\ : Span4Mux_v
    port map (
            O => \N__6167\,
            I => \N__6147\
        );

    \I__1397\ : Span4Mux_s3_h
    port map (
            O => \N__6162\,
            I => \N__6140\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__6159\,
            I => \N__6140\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__6156\,
            I => \N__6140\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__6153\,
            I => \N__6137\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__6150\,
            I => \N__6134\
        );

    \I__1392\ : Span4Mux_h
    port map (
            O => \N__6147\,
            I => \N__6129\
        );

    \I__1391\ : Span4Mux_v
    port map (
            O => \N__6140\,
            I => \N__6129\
        );

    \I__1390\ : Span4Mux_v
    port map (
            O => \N__6137\,
            I => \N__6126\
        );

    \I__1389\ : Odrv12
    port map (
            O => \N__6134\,
            I => \SIZ_c_1\
        );

    \I__1388\ : Odrv4
    port map (
            O => \N__6129\,
            I => \SIZ_c_1\
        );

    \I__1387\ : Odrv4
    port map (
            O => \N__6126\,
            I => \SIZ_c_1\
        );

    \I__1386\ : CascadeMux
    port map (
            O => \N__6119\,
            I => \N__6115\
        );

    \I__1385\ : InMux
    port map (
            O => \N__6118\,
            I => \N__6109\
        );

    \I__1384\ : InMux
    port map (
            O => \N__6115\,
            I => \N__6106\
        );

    \I__1383\ : InMux
    port map (
            O => \N__6114\,
            I => \N__6103\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__6113\,
            I => \N__6100\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__6112\,
            I => \N__6097\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__6109\,
            I => \N__6094\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__6106\,
            I => \N__6089\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__6103\,
            I => \N__6089\
        );

    \I__1377\ : InMux
    port map (
            O => \N__6100\,
            I => \N__6084\
        );

    \I__1376\ : InMux
    port map (
            O => \N__6097\,
            I => \N__6084\
        );

    \I__1375\ : Span4Mux_s3_v
    port map (
            O => \N__6094\,
            I => \N__6077\
        );

    \I__1374\ : Span4Mux_v
    port map (
            O => \N__6089\,
            I => \N__6077\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__6084\,
            I => \N__6074\
        );

    \I__1372\ : InMux
    port map (
            O => \N__6083\,
            I => \N__6071\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__6082\,
            I => \N__6068\
        );

    \I__1370\ : Span4Mux_h
    port map (
            O => \N__6077\,
            I => \N__6061\
        );

    \I__1369\ : Span4Mux_s3_v
    port map (
            O => \N__6074\,
            I => \N__6061\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__6071\,
            I => \N__6061\
        );

    \I__1367\ : InMux
    port map (
            O => \N__6068\,
            I => \N__6058\
        );

    \I__1366\ : Span4Mux_s3_h
    port map (
            O => \N__6061\,
            I => \N__6052\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__6058\,
            I => \N__6052\
        );

    \I__1364\ : InMux
    port map (
            O => \N__6057\,
            I => \N__6049\
        );

    \I__1363\ : Span4Mux_v
    port map (
            O => \N__6052\,
            I => \N__6044\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__6049\,
            I => \N__6044\
        );

    \I__1361\ : Odrv4
    port map (
            O => \N__6044\,
            I => \SIZ_c_0\
        );

    \I__1360\ : CascadeMux
    port map (
            O => \N__6041\,
            I => \N__6038\
        );

    \I__1359\ : InMux
    port map (
            O => \N__6038\,
            I => \N__6035\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__6035\,
            I => \N__6032\
        );

    \I__1357\ : Span4Mux_v
    port map (
            O => \N__6032\,
            I => \N__6029\
        );

    \I__1356\ : Odrv4
    port map (
            O => \N__6029\,
            I => \U400_BYTE_ENABLE.N_54_i\
        );

    \I__1355\ : InMux
    port map (
            O => \N__6026\,
            I => \N__6022\
        );

    \I__1354\ : InMux
    port map (
            O => \N__6025\,
            I => \N__6018\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__6022\,
            I => \N__6015\
        );

    \I__1352\ : InMux
    port map (
            O => \N__6021\,
            I => \N__6012\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__6018\,
            I => \N__6009\
        );

    \I__1350\ : Span4Mux_v
    port map (
            O => \N__6015\,
            I => \N__6004\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__6012\,
            I => \N__6004\
        );

    \I__1348\ : Span4Mux_v
    port map (
            O => \N__6009\,
            I => \N__6001\
        );

    \I__1347\ : Sp12to4
    port map (
            O => \N__6004\,
            I => \N__5998\
        );

    \I__1346\ : Span4Mux_v
    port map (
            O => \N__6001\,
            I => \N__5995\
        );

    \I__1345\ : Span12Mux_v
    port map (
            O => \N__5998\,
            I => \N__5992\
        );

    \I__1344\ : Span4Mux_h
    port map (
            O => \N__5995\,
            I => \N__5989\
        );

    \I__1343\ : Odrv12
    port map (
            O => \N__5992\,
            I => \A_c_0\
        );

    \I__1342\ : Odrv4
    port map (
            O => \N__5989\,
            I => \A_c_0\
        );

    \I__1341\ : IoInMux
    port map (
            O => \N__5984\,
            I => \N__5981\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__5981\,
            I => \N__5975\
        );

    \I__1339\ : InMux
    port map (
            O => \N__5980\,
            I => \N__5972\
        );

    \I__1338\ : InMux
    port map (
            O => \N__5979\,
            I => \N__5969\
        );

    \I__1337\ : CascadeMux
    port map (
            O => \N__5978\,
            I => \N__5966\
        );

    \I__1336\ : IoSpan4Mux
    port map (
            O => \N__5975\,
            I => \N__5963\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__5972\,
            I => \N__5960\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__5969\,
            I => \N__5957\
        );

    \I__1333\ : InMux
    port map (
            O => \N__5966\,
            I => \N__5954\
        );

    \I__1332\ : Span4Mux_s2_h
    port map (
            O => \N__5963\,
            I => \N__5945\
        );

    \I__1331\ : Span4Mux_v
    port map (
            O => \N__5960\,
            I => \N__5945\
        );

    \I__1330\ : Span4Mux_h
    port map (
            O => \N__5957\,
            I => \N__5945\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__5954\,
            I => \N__5945\
        );

    \I__1328\ : Span4Mux_v
    port map (
            O => \N__5945\,
            I => \N__5942\
        );

    \I__1327\ : Span4Mux_h
    port map (
            O => \N__5942\,
            I => \N__5939\
        );

    \I__1326\ : Odrv4
    port map (
            O => \N__5939\,
            I => \RAM_SPACE_i_o3dup\
        );

    \I__1325\ : CascadeMux
    port map (
            O => \N__5936\,
            I => \U400_BYTE_ENABLE.N_54_i_cascade_\
        );

    \I__1324\ : InMux
    port map (
            O => \N__5933\,
            I => \N__5927\
        );

    \I__1323\ : InMux
    port map (
            O => \N__5932\,
            I => \N__5927\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__5927\,
            I => \N__5923\
        );

    \I__1321\ : InMux
    port map (
            O => \N__5926\,
            I => \N__5920\
        );

    \I__1320\ : Span4Mux_v
    port map (
            O => \N__5923\,
            I => \N__5914\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__5920\,
            I => \N__5914\
        );

    \I__1318\ : InMux
    port map (
            O => \N__5919\,
            I => \N__5911\
        );

    \I__1317\ : Span4Mux_v
    port map (
            O => \N__5914\,
            I => \N__5908\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__5911\,
            I => \N__5905\
        );

    \I__1315\ : Span4Mux_v
    port map (
            O => \N__5908\,
            I => \N__5902\
        );

    \I__1314\ : Sp12to4
    port map (
            O => \N__5905\,
            I => \N__5899\
        );

    \I__1313\ : Sp12to4
    port map (
            O => \N__5902\,
            I => \N__5894\
        );

    \I__1312\ : Span12Mux_v
    port map (
            O => \N__5899\,
            I => \N__5894\
        );

    \I__1311\ : Odrv12
    port map (
            O => \N__5894\,
            I => \A_c_1\
        );

    \I__1310\ : IoInMux
    port map (
            O => \N__5891\,
            I => \N__5888\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__5888\,
            I => \N__5885\
        );

    \I__1308\ : Span12Mux_s7_v
    port map (
            O => \N__5885\,
            I => \N__5882\
        );

    \I__1307\ : Odrv12
    port map (
            O => \N__5882\,
            I => \N_49\
        );

    \I__1306\ : InMux
    port map (
            O => \N__5879\,
            I => \N__5875\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__5878\,
            I => \N__5869\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__5875\,
            I => \N__5863\
        );

    \I__1303\ : InMux
    port map (
            O => \N__5874\,
            I => \N__5858\
        );

    \I__1302\ : InMux
    port map (
            O => \N__5873\,
            I => \N__5853\
        );

    \I__1301\ : InMux
    port map (
            O => \N__5872\,
            I => \N__5853\
        );

    \I__1300\ : InMux
    port map (
            O => \N__5869\,
            I => \N__5850\
        );

    \I__1299\ : InMux
    port map (
            O => \N__5868\,
            I => \N__5847\
        );

    \I__1298\ : InMux
    port map (
            O => \N__5867\,
            I => \N__5844\
        );

    \I__1297\ : InMux
    port map (
            O => \N__5866\,
            I => \N__5840\
        );

    \I__1296\ : Span4Mux_s1_v
    port map (
            O => \N__5863\,
            I => \N__5837\
        );

    \I__1295\ : InMux
    port map (
            O => \N__5862\,
            I => \N__5832\
        );

    \I__1294\ : InMux
    port map (
            O => \N__5861\,
            I => \N__5832\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__5858\,
            I => \N__5828\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__5853\,
            I => \N__5825\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__5850\,
            I => \N__5818\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__5847\,
            I => \N__5818\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5844\,
            I => \N__5818\
        );

    \I__1288\ : InMux
    port map (
            O => \N__5843\,
            I => \N__5815\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__5840\,
            I => \N__5808\
        );

    \I__1286\ : Span4Mux_h
    port map (
            O => \N__5837\,
            I => \N__5808\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__5832\,
            I => \N__5808\
        );

    \I__1284\ : InMux
    port map (
            O => \N__5831\,
            I => \N__5805\
        );

    \I__1283\ : Span4Mux_s3_h
    port map (
            O => \N__5828\,
            I => \N__5802\
        );

    \I__1282\ : Span4Mux_s3_h
    port map (
            O => \N__5825\,
            I => \N__5799\
        );

    \I__1281\ : Span12Mux_s8_h
    port map (
            O => \N__5818\,
            I => \N__5796\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__5815\,
            I => \N__5791\
        );

    \I__1279\ : Span4Mux_v
    port map (
            O => \N__5808\,
            I => \N__5791\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__5805\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_1\
        );

    \I__1277\ : Odrv4
    port map (
            O => \N__5802\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_1\
        );

    \I__1276\ : Odrv4
    port map (
            O => \N__5799\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_1\
        );

    \I__1275\ : Odrv12
    port map (
            O => \N__5796\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_1\
        );

    \I__1274\ : Odrv4
    port map (
            O => \N__5791\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_1\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__5780\,
            I => \N__5777\
        );

    \I__1272\ : InMux
    port map (
            O => \N__5777\,
            I => \N__5774\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__5774\,
            I => \N__5771\
        );

    \I__1270\ : IoSpan4Mux
    port map (
            O => \N__5771\,
            I => \N__5768\
        );

    \I__1269\ : Odrv4
    port map (
            O => \N__5768\,
            I => \A_c_14\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5765\,
            I => \N__5760\
        );

    \I__1267\ : InMux
    port map (
            O => \N__5764\,
            I => \N__5755\
        );

    \I__1266\ : InMux
    port map (
            O => \N__5763\,
            I => \N__5755\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__5760\,
            I => \N__5748\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__5755\,
            I => \N__5745\
        );

    \I__1263\ : InMux
    port map (
            O => \N__5754\,
            I => \N__5742\
        );

    \I__1262\ : InMux
    port map (
            O => \N__5753\,
            I => \N__5739\
        );

    \I__1261\ : InMux
    port map (
            O => \N__5752\,
            I => \N__5736\
        );

    \I__1260\ : InMux
    port map (
            O => \N__5751\,
            I => \N__5733\
        );

    \I__1259\ : Span4Mux_s1_v
    port map (
            O => \N__5748\,
            I => \N__5726\
        );

    \I__1258\ : Span4Mux_h
    port map (
            O => \N__5745\,
            I => \N__5726\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__5742\,
            I => \N__5726\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__5739\,
            I => \N__5717\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__5736\,
            I => \N__5717\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__5733\,
            I => \N__5714\
        );

    \I__1253\ : Span4Mux_v
    port map (
            O => \N__5726\,
            I => \N__5710\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5725\,
            I => \N__5707\
        );

    \I__1251\ : InMux
    port map (
            O => \N__5724\,
            I => \N__5702\
        );

    \I__1250\ : InMux
    port map (
            O => \N__5723\,
            I => \N__5702\
        );

    \I__1249\ : InMux
    port map (
            O => \N__5722\,
            I => \N__5699\
        );

    \I__1248\ : Span4Mux_v
    port map (
            O => \N__5717\,
            I => \N__5696\
        );

    \I__1247\ : Span4Mux_h
    port map (
            O => \N__5714\,
            I => \N__5693\
        );

    \I__1246\ : InMux
    port map (
            O => \N__5713\,
            I => \N__5690\
        );

    \I__1245\ : Span4Mux_h
    port map (
            O => \N__5710\,
            I => \N__5687\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__5707\,
            I => \N__5682\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__5702\,
            I => \N__5682\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__5699\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_0\
        );

    \I__1241\ : Odrv4
    port map (
            O => \N__5696\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_0\
        );

    \I__1240\ : Odrv4
    port map (
            O => \N__5693\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_0\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__5690\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_0\
        );

    \I__1238\ : Odrv4
    port map (
            O => \N__5687\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_0\
        );

    \I__1237\ : Odrv12
    port map (
            O => \N__5682\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_0\
        );

    \I__1236\ : InMux
    port map (
            O => \N__5669\,
            I => \N__5664\
        );

    \I__1235\ : InMux
    port map (
            O => \N__5668\,
            I => \N__5661\
        );

    \I__1234\ : InMux
    port map (
            O => \N__5667\,
            I => \N__5658\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__5664\,
            I => \N__5655\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__5661\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_1\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__5658\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_1\
        );

    \I__1230\ : Odrv4
    port map (
            O => \N__5655\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_1\
        );

    \I__1229\ : InMux
    port map (
            O => \N__5648\,
            I => \N__5645\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__5645\,
            I => \U400_SDRAM.TA_OUT_5_0\
        );

    \I__1227\ : CascadeMux
    port map (
            O => \N__5642\,
            I => \N__5639\
        );

    \I__1226\ : InMux
    port map (
            O => \N__5639\,
            I => \N__5636\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__5636\,
            I => \N__5633\
        );

    \I__1224\ : Span4Mux_s2_v
    port map (
            O => \N__5633\,
            I => \N__5630\
        );

    \I__1223\ : Sp12to4
    port map (
            O => \N__5630\,
            I => \N__5627\
        );

    \I__1222\ : Span12Mux_s10_h
    port map (
            O => \N__5627\,
            I => \N__5624\
        );

    \I__1221\ : Span12Mux_v
    port map (
            O => \N__5624\,
            I => \N__5621\
        );

    \I__1220\ : Odrv12
    port map (
            O => \N__5621\,
            I => \A_c_24\
        );

    \I__1219\ : IoInMux
    port map (
            O => \N__5618\,
            I => \N__5615\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__5615\,
            I => \N__5612\
        );

    \I__1217\ : Odrv4
    port map (
            O => \N__5612\,
            I => \MA_c_11\
        );

    \I__1216\ : InMux
    port map (
            O => \N__5609\,
            I => \N__5606\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__5606\,
            I => \N__5603\
        );

    \I__1214\ : Odrv12
    port map (
            O => \N__5603\,
            I => \A_c_11\
        );

    \I__1213\ : IoInMux
    port map (
            O => \N__5600\,
            I => \N__5597\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__5597\,
            I => \N__5594\
        );

    \I__1211\ : Span4Mux_s1_v
    port map (
            O => \N__5594\,
            I => \N__5591\
        );

    \I__1210\ : Odrv4
    port map (
            O => \N__5591\,
            I => \MA_c_9\
        );

    \I__1209\ : InMux
    port map (
            O => \N__5588\,
            I => \N__5585\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__5585\,
            I => \N__5582\
        );

    \I__1207\ : Span12Mux_s11_v
    port map (
            O => \N__5582\,
            I => \N__5579\
        );

    \I__1206\ : Odrv12
    port map (
            O => \N__5579\,
            I => \A_c_25\
        );

    \I__1205\ : CascadeMux
    port map (
            O => \N__5576\,
            I => \N__5573\
        );

    \I__1204\ : InMux
    port map (
            O => \N__5573\,
            I => \N__5570\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__5570\,
            I => \N__5567\
        );

    \I__1202\ : Odrv12
    port map (
            O => \N__5567\,
            I => \A_c_10\
        );

    \I__1201\ : IoInMux
    port map (
            O => \N__5564\,
            I => \N__5561\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__5561\,
            I => \N__5558\
        );

    \I__1199\ : IoSpan4Mux
    port map (
            O => \N__5558\,
            I => \N__5555\
        );

    \I__1198\ : Odrv4
    port map (
            O => \N__5555\,
            I => \MA_c_8\
        );

    \I__1197\ : InMux
    port map (
            O => \N__5552\,
            I => \N__5547\
        );

    \I__1196\ : InMux
    port map (
            O => \N__5551\,
            I => \N__5544\
        );

    \I__1195\ : InMux
    port map (
            O => \N__5550\,
            I => \N__5541\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__5547\,
            I => \N__5538\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__5544\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_4\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__5541\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_4\
        );

    \I__1191\ : Odrv4
    port map (
            O => \N__5538\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_4\
        );

    \I__1190\ : InMux
    port map (
            O => \N__5531\,
            I => \N__5528\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5528\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_5\
        );

    \I__1188\ : InMux
    port map (
            O => \N__5525\,
            I => \N__5520\
        );

    \I__1187\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5515\
        );

    \I__1186\ : InMux
    port map (
            O => \N__5523\,
            I => \N__5515\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__5520\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_2\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__5515\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_2\
        );

    \I__1183\ : InMux
    port map (
            O => \N__5510\,
            I => \N__5506\
        );

    \I__1182\ : InMux
    port map (
            O => \N__5509\,
            I => \N__5503\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__5506\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_3\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__5503\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_3\
        );

    \I__1179\ : ClkMux
    port map (
            O => \N__5498\,
            I => \N__5423\
        );

    \I__1178\ : ClkMux
    port map (
            O => \N__5497\,
            I => \N__5423\
        );

    \I__1177\ : ClkMux
    port map (
            O => \N__5496\,
            I => \N__5423\
        );

    \I__1176\ : ClkMux
    port map (
            O => \N__5495\,
            I => \N__5423\
        );

    \I__1175\ : ClkMux
    port map (
            O => \N__5494\,
            I => \N__5423\
        );

    \I__1174\ : ClkMux
    port map (
            O => \N__5493\,
            I => \N__5423\
        );

    \I__1173\ : ClkMux
    port map (
            O => \N__5492\,
            I => \N__5423\
        );

    \I__1172\ : ClkMux
    port map (
            O => \N__5491\,
            I => \N__5423\
        );

    \I__1171\ : ClkMux
    port map (
            O => \N__5490\,
            I => \N__5423\
        );

    \I__1170\ : ClkMux
    port map (
            O => \N__5489\,
            I => \N__5423\
        );

    \I__1169\ : ClkMux
    port map (
            O => \N__5488\,
            I => \N__5423\
        );

    \I__1168\ : ClkMux
    port map (
            O => \N__5487\,
            I => \N__5423\
        );

    \I__1167\ : ClkMux
    port map (
            O => \N__5486\,
            I => \N__5423\
        );

    \I__1166\ : ClkMux
    port map (
            O => \N__5485\,
            I => \N__5423\
        );

    \I__1165\ : ClkMux
    port map (
            O => \N__5484\,
            I => \N__5423\
        );

    \I__1164\ : ClkMux
    port map (
            O => \N__5483\,
            I => \N__5423\
        );

    \I__1163\ : ClkMux
    port map (
            O => \N__5482\,
            I => \N__5423\
        );

    \I__1162\ : ClkMux
    port map (
            O => \N__5481\,
            I => \N__5423\
        );

    \I__1161\ : ClkMux
    port map (
            O => \N__5480\,
            I => \N__5423\
        );

    \I__1160\ : ClkMux
    port map (
            O => \N__5479\,
            I => \N__5423\
        );

    \I__1159\ : ClkMux
    port map (
            O => \N__5478\,
            I => \N__5423\
        );

    \I__1158\ : ClkMux
    port map (
            O => \N__5477\,
            I => \N__5423\
        );

    \I__1157\ : ClkMux
    port map (
            O => \N__5476\,
            I => \N__5423\
        );

    \I__1156\ : ClkMux
    port map (
            O => \N__5475\,
            I => \N__5423\
        );

    \I__1155\ : ClkMux
    port map (
            O => \N__5474\,
            I => \N__5423\
        );

    \I__1154\ : GlobalMux
    port map (
            O => \N__5423\,
            I => \N__5420\
        );

    \I__1153\ : gio2CtrlBuf
    port map (
            O => \N__5420\,
            I => \CLK40_c_g\
        );

    \I__1152\ : InMux
    port map (
            O => \N__5417\,
            I => \N__5413\
        );

    \I__1151\ : InMux
    port map (
            O => \N__5416\,
            I => \N__5410\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__5413\,
            I => \N__5407\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__5410\,
            I => \N__5402\
        );

    \I__1148\ : Span4Mux_h
    port map (
            O => \N__5407\,
            I => \N__5399\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5406\,
            I => \N__5396\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5405\,
            I => \N__5393\
        );

    \I__1145\ : Odrv12
    port map (
            O => \N__5402\,
            I => \U400_SDRAM.SDRAM_CMD_1_sqmuxa_1\
        );

    \I__1144\ : Odrv4
    port map (
            O => \N__5399\,
            I => \U400_SDRAM.SDRAM_CMD_1_sqmuxa_1\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__5396\,
            I => \U400_SDRAM.SDRAM_CMD_1_sqmuxa_1\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__5393\,
            I => \U400_SDRAM.SDRAM_CMD_1_sqmuxa_1\
        );

    \I__1141\ : InMux
    port map (
            O => \N__5384\,
            I => \N__5378\
        );

    \I__1140\ : InMux
    port map (
            O => \N__5383\,
            I => \N__5375\
        );

    \I__1139\ : InMux
    port map (
            O => \N__5382\,
            I => \N__5372\
        );

    \I__1138\ : InMux
    port map (
            O => \N__5381\,
            I => \N__5369\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__5378\,
            I => \U400_SDRAM.BURSTZ0\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__5375\,
            I => \U400_SDRAM.BURSTZ0\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__5372\,
            I => \U400_SDRAM.BURSTZ0\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__5369\,
            I => \U400_SDRAM.BURSTZ0\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5360\,
            I => \N__5357\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__5357\,
            I => \U400_SDRAM.TA_COUNTER_srsts_0_a4_0_0\
        );

    \I__1131\ : InMux
    port map (
            O => \N__5354\,
            I => \N__5351\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__5351\,
            I => \U400_SDRAM.N_243_0\
        );

    \I__1129\ : InMux
    port map (
            O => \N__5348\,
            I => \N__5343\
        );

    \I__1128\ : InMux
    port map (
            O => \N__5347\,
            I => \N__5340\
        );

    \I__1127\ : InMux
    port map (
            O => \N__5346\,
            I => \N__5332\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__5343\,
            I => \N__5327\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__5340\,
            I => \N__5327\
        );

    \I__1124\ : InMux
    port map (
            O => \N__5339\,
            I => \N__5324\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__5338\,
            I => \N__5319\
        );

    \I__1122\ : InMux
    port map (
            O => \N__5337\,
            I => \N__5316\
        );

    \I__1121\ : InMux
    port map (
            O => \N__5336\,
            I => \N__5313\
        );

    \I__1120\ : CascadeMux
    port map (
            O => \N__5335\,
            I => \N__5310\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__5332\,
            I => \N__5305\
        );

    \I__1118\ : Span4Mux_v
    port map (
            O => \N__5327\,
            I => \N__5300\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__5324\,
            I => \N__5300\
        );

    \I__1116\ : InMux
    port map (
            O => \N__5323\,
            I => \N__5297\
        );

    \I__1115\ : CascadeMux
    port map (
            O => \N__5322\,
            I => \N__5293\
        );

    \I__1114\ : InMux
    port map (
            O => \N__5319\,
            I => \N__5289\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__5316\,
            I => \N__5286\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__5313\,
            I => \N__5283\
        );

    \I__1111\ : InMux
    port map (
            O => \N__5310\,
            I => \N__5280\
        );

    \I__1110\ : InMux
    port map (
            O => \N__5309\,
            I => \N__5277\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__5308\,
            I => \N__5274\
        );

    \I__1108\ : Span4Mux_h
    port map (
            O => \N__5305\,
            I => \N__5266\
        );

    \I__1107\ : Span4Mux_h
    port map (
            O => \N__5300\,
            I => \N__5266\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__5297\,
            I => \N__5266\
        );

    \I__1105\ : InMux
    port map (
            O => \N__5296\,
            I => \N__5263\
        );

    \I__1104\ : InMux
    port map (
            O => \N__5293\,
            I => \N__5258\
        );

    \I__1103\ : InMux
    port map (
            O => \N__5292\,
            I => \N__5258\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__5289\,
            I => \N__5255\
        );

    \I__1101\ : Span4Mux_h
    port map (
            O => \N__5286\,
            I => \N__5246\
        );

    \I__1100\ : Span4Mux_v
    port map (
            O => \N__5283\,
            I => \N__5246\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__5280\,
            I => \N__5246\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__5277\,
            I => \N__5246\
        );

    \I__1097\ : InMux
    port map (
            O => \N__5274\,
            I => \N__5241\
        );

    \I__1096\ : InMux
    port map (
            O => \N__5273\,
            I => \N__5241\
        );

    \I__1095\ : Span4Mux_h
    port map (
            O => \N__5266\,
            I => \N__5234\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__5263\,
            I => \N__5234\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__5258\,
            I => \N__5234\
        );

    \I__1092\ : Sp12to4
    port map (
            O => \N__5255\,
            I => \N__5231\
        );

    \I__1091\ : Span4Mux_v
    port map (
            O => \N__5246\,
            I => \N__5228\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__5241\,
            I => \N__5225\
        );

    \I__1089\ : Span4Mux_v
    port map (
            O => \N__5234\,
            I => \N__5222\
        );

    \I__1088\ : Span12Mux_s8_v
    port map (
            O => \N__5231\,
            I => \N__5219\
        );

    \I__1087\ : Sp12to4
    port map (
            O => \N__5228\,
            I => \N__5214\
        );

    \I__1086\ : Span12Mux_s8_v
    port map (
            O => \N__5225\,
            I => \N__5214\
        );

    \I__1085\ : Span4Mux_h
    port map (
            O => \N__5222\,
            I => \N__5211\
        );

    \I__1084\ : Odrv12
    port map (
            O => \N__5219\,
            I => \RESETn_c\
        );

    \I__1083\ : Odrv12
    port map (
            O => \N__5214\,
            I => \RESETn_c\
        );

    \I__1082\ : Odrv4
    port map (
            O => \N__5211\,
            I => \RESETn_c\
        );

    \I__1081\ : InMux
    port map (
            O => \N__5204\,
            I => \N__5199\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5203\,
            I => \N__5196\
        );

    \I__1079\ : InMux
    port map (
            O => \N__5202\,
            I => \N__5193\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__5199\,
            I => \N__5190\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__5196\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_0\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__5193\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_0\
        );

    \I__1075\ : Odrv4
    port map (
            O => \N__5190\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_0\
        );

    \I__1074\ : CascadeMux
    port map (
            O => \N__5183\,
            I => \U400_SDRAM.N_243_0_cascade_\
        );

    \I__1073\ : InMux
    port map (
            O => \N__5180\,
            I => \N__5175\
        );

    \I__1072\ : InMux
    port map (
            O => \N__5179\,
            I => \N__5169\
        );

    \I__1071\ : InMux
    port map (
            O => \N__5178\,
            I => \N__5169\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__5175\,
            I => \N__5166\
        );

    \I__1069\ : InMux
    port map (
            O => \N__5174\,
            I => \N__5162\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__5169\,
            I => \N__5159\
        );

    \I__1067\ : Span4Mux_v
    port map (
            O => \N__5166\,
            I => \N__5156\
        );

    \I__1066\ : InMux
    port map (
            O => \N__5165\,
            I => \N__5153\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__5162\,
            I => \U400_SDRAM.TACKZ0\
        );

    \I__1064\ : Odrv4
    port map (
            O => \N__5159\,
            I => \U400_SDRAM.TACKZ0\
        );

    \I__1063\ : Odrv4
    port map (
            O => \N__5156\,
            I => \U400_SDRAM.TACKZ0\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__5153\,
            I => \U400_SDRAM.TACKZ0\
        );

    \I__1061\ : InMux
    port map (
            O => \N__5144\,
            I => \N__5141\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__5141\,
            I => \U400_SDRAM.N_241_0_en\
        );

    \I__1059\ : CascadeMux
    port map (
            O => \N__5138\,
            I => \N__5134\
        );

    \I__1058\ : InMux
    port map (
            O => \N__5137\,
            I => \N__5131\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5134\,
            I => \N__5128\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__5131\,
            I => \U400_SDRAM.un1_TA_COUNTER_6_0_0\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__5128\,
            I => \U400_SDRAM.un1_TA_COUNTER_6_0_0\
        );

    \I__1054\ : InMux
    port map (
            O => \N__5123\,
            I => \N__5119\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5122\,
            I => \N__5116\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__5119\,
            I => \U400_SDRAM.N_244_0\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__5116\,
            I => \U400_SDRAM.N_244_0\
        );

    \I__1050\ : IoInMux
    port map (
            O => \N__5111\,
            I => \N__5107\
        );

    \I__1049\ : CascadeMux
    port map (
            O => \N__5110\,
            I => \N__5104\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__5107\,
            I => \N__5101\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5104\,
            I => \N__5098\
        );

    \I__1046\ : Odrv12
    port map (
            O => \N__5101\,
            I => \TA_OUT\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__5098\,
            I => \TA_OUT\
        );

    \I__1044\ : IoInMux
    port map (
            O => \N__5093\,
            I => \N__5090\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__5090\,
            I => \N__5087\
        );

    \I__1042\ : Odrv12
    port map (
            O => \N__5087\,
            I => \N_53\
        );

    \I__1041\ : CascadeMux
    port map (
            O => \N__5084\,
            I => \N__5078\
        );

    \I__1040\ : InMux
    port map (
            O => \N__5083\,
            I => \N__5074\
        );

    \I__1039\ : InMux
    port map (
            O => \N__5082\,
            I => \N__5069\
        );

    \I__1038\ : InMux
    port map (
            O => \N__5081\,
            I => \N__5069\
        );

    \I__1037\ : InMux
    port map (
            O => \N__5078\,
            I => \N__5063\
        );

    \I__1036\ : InMux
    port map (
            O => \N__5077\,
            I => \N__5060\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__5074\,
            I => \N__5055\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__5069\,
            I => \N__5055\
        );

    \I__1033\ : InMux
    port map (
            O => \N__5068\,
            I => \N__5044\
        );

    \I__1032\ : InMux
    port map (
            O => \N__5067\,
            I => \N__5039\
        );

    \I__1031\ : InMux
    port map (
            O => \N__5066\,
            I => \N__5039\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__5063\,
            I => \N__5032\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__5060\,
            I => \N__5032\
        );

    \I__1028\ : Span4Mux_h
    port map (
            O => \N__5055\,
            I => \N__5032\
        );

    \I__1027\ : InMux
    port map (
            O => \N__5054\,
            I => \N__5027\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5053\,
            I => \N__5027\
        );

    \I__1025\ : InMux
    port map (
            O => \N__5052\,
            I => \N__5020\
        );

    \I__1024\ : InMux
    port map (
            O => \N__5051\,
            I => \N__5020\
        );

    \I__1023\ : InMux
    port map (
            O => \N__5050\,
            I => \N__5020\
        );

    \I__1022\ : InMux
    port map (
            O => \N__5049\,
            I => \N__5017\
        );

    \I__1021\ : InMux
    port map (
            O => \N__5048\,
            I => \N__5014\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5047\,
            I => \N__5011\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__5044\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__5039\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1017\ : Odrv4
    port map (
            O => \N__5032\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__5027\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__5020\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__5017\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__5014\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__5011\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1011\ : InMux
    port map (
            O => \N__4994\,
            I => \N__4991\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__4991\,
            I => \U400_SDRAM.N_28\
        );

    \I__1009\ : InMux
    port map (
            O => \N__4988\,
            I => \N__4985\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__4985\,
            I => \U400_SDRAM.N_110\
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__4982\,
            I => \N__4979\
        );

    \I__1006\ : InMux
    port map (
            O => \N__4979\,
            I => \N__4973\
        );

    \I__1005\ : InMux
    port map (
            O => \N__4978\,
            I => \N__4973\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__4973\,
            I => \N__4965\
        );

    \I__1003\ : InMux
    port map (
            O => \N__4972\,
            I => \N__4958\
        );

    \I__1002\ : InMux
    port map (
            O => \N__4971\,
            I => \N__4958\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4970\,
            I => \N__4958\
        );

    \I__1000\ : InMux
    port map (
            O => \N__4969\,
            I => \N__4953\
        );

    \I__999\ : InMux
    port map (
            O => \N__4968\,
            I => \N__4950\
        );

    \I__998\ : Span4Mux_h
    port map (
            O => \N__4965\,
            I => \N__4947\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__4958\,
            I => \N__4944\
        );

    \I__996\ : InMux
    port map (
            O => \N__4957\,
            I => \N__4939\
        );

    \I__995\ : InMux
    port map (
            O => \N__4956\,
            I => \N__4939\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__4953\,
            I => \N__4934\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__4950\,
            I => \N__4934\
        );

    \I__992\ : Odrv4
    port map (
            O => \N__4947\,
            I => \U400_SDRAM.WRITE_CYCLEZ0\
        );

    \I__991\ : Odrv4
    port map (
            O => \N__4944\,
            I => \U400_SDRAM.WRITE_CYCLEZ0\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__4939\,
            I => \U400_SDRAM.WRITE_CYCLEZ0\
        );

    \I__989\ : Odrv4
    port map (
            O => \N__4934\,
            I => \U400_SDRAM.WRITE_CYCLEZ0\
        );

    \I__988\ : InMux
    port map (
            O => \N__4925\,
            I => \N__4922\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__4922\,
            I => \U400_SDRAM.N_13\
        );

    \I__986\ : InMux
    port map (
            O => \N__4919\,
            I => \N__4909\
        );

    \I__985\ : InMux
    port map (
            O => \N__4918\,
            I => \N__4904\
        );

    \I__984\ : InMux
    port map (
            O => \N__4917\,
            I => \N__4904\
        );

    \I__983\ : InMux
    port map (
            O => \N__4916\,
            I => \N__4901\
        );

    \I__982\ : InMux
    port map (
            O => \N__4915\,
            I => \N__4897\
        );

    \I__981\ : InMux
    port map (
            O => \N__4914\,
            I => \N__4890\
        );

    \I__980\ : InMux
    port map (
            O => \N__4913\,
            I => \N__4890\
        );

    \I__979\ : InMux
    port map (
            O => \N__4912\,
            I => \N__4890\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__4909\,
            I => \N__4881\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__4904\,
            I => \N__4881\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__4901\,
            I => \N__4881\
        );

    \I__975\ : InMux
    port map (
            O => \N__4900\,
            I => \N__4878\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__4897\,
            I => \N__4873\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__4890\,
            I => \N__4873\
        );

    \I__972\ : InMux
    port map (
            O => \N__4889\,
            I => \N__4870\
        );

    \I__971\ : InMux
    port map (
            O => \N__4888\,
            I => \N__4867\
        );

    \I__970\ : Odrv4
    port map (
            O => \N__4881\,
            I => \U400_SDRAM.N_44\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__4878\,
            I => \U400_SDRAM.N_44\
        );

    \I__968\ : Odrv4
    port map (
            O => \N__4873\,
            I => \U400_SDRAM.N_44\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__4870\,
            I => \U400_SDRAM.N_44\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4867\,
            I => \U400_SDRAM.N_44\
        );

    \I__965\ : CascadeMux
    port map (
            O => \N__4856\,
            I => \N__4852\
        );

    \I__964\ : InMux
    port map (
            O => \N__4855\,
            I => \N__4847\
        );

    \I__963\ : InMux
    port map (
            O => \N__4852\,
            I => \N__4847\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__4847\,
            I => \N__4844\
        );

    \I__961\ : Odrv12
    port map (
            O => \N__4844\,
            I => \U400_SDRAM.N_8\
        );

    \I__960\ : CascadeMux
    port map (
            O => \N__4841\,
            I => \U400_SDRAM.N_13_cascade_\
        );

    \I__959\ : InMux
    port map (
            O => \N__4838\,
            I => \N__4835\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__4835\,
            I => \N__4832\
        );

    \I__957\ : Span4Mux_h
    port map (
            O => \N__4832\,
            I => \N__4829\
        );

    \I__956\ : Odrv4
    port map (
            O => \N__4829\,
            I => \U400_SDRAM.N_76\
        );

    \I__955\ : InMux
    port map (
            O => \N__4826\,
            I => \N__4823\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4823\,
            I => \N__4820\
        );

    \I__953\ : Odrv12
    port map (
            O => \N__4820\,
            I => \U400_SDRAM.un1_SDRAM_COUNTER59_1_1_0\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__4817\,
            I => \N__4814\
        );

    \I__951\ : InMux
    port map (
            O => \N__4814\,
            I => \N__4809\
        );

    \I__950\ : CascadeMux
    port map (
            O => \N__4813\,
            I => \N__4806\
        );

    \I__949\ : InMux
    port map (
            O => \N__4812\,
            I => \N__4802\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__4809\,
            I => \N__4799\
        );

    \I__947\ : InMux
    port map (
            O => \N__4806\,
            I => \N__4796\
        );

    \I__946\ : InMux
    port map (
            O => \N__4805\,
            I => \N__4793\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4802\,
            I => \U400_SDRAM.N_46\
        );

    \I__944\ : Odrv4
    port map (
            O => \N__4799\,
            I => \U400_SDRAM.N_46\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__4796\,
            I => \U400_SDRAM.N_46\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__4793\,
            I => \U400_SDRAM.N_46\
        );

    \I__941\ : CascadeMux
    port map (
            O => \N__4784\,
            I => \U400_SDRAM.N_33_cascade_\
        );

    \I__940\ : InMux
    port map (
            O => \N__4781\,
            I => \N__4778\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__4778\,
            I => \N__4774\
        );

    \I__938\ : CascadeMux
    port map (
            O => \N__4777\,
            I => \N__4770\
        );

    \I__937\ : Span4Mux_v
    port map (
            O => \N__4774\,
            I => \N__4767\
        );

    \I__936\ : InMux
    port map (
            O => \N__4773\,
            I => \N__4762\
        );

    \I__935\ : InMux
    port map (
            O => \N__4770\,
            I => \N__4762\
        );

    \I__934\ : Odrv4
    port map (
            O => \N__4767\,
            I => \U400_SDRAM.N_67\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4762\,
            I => \U400_SDRAM.N_67\
        );

    \I__932\ : InMux
    port map (
            O => \N__4757\,
            I => \N__4754\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4754\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_1_66_i_0_1\
        );

    \I__930\ : InMux
    port map (
            O => \N__4751\,
            I => \N__4745\
        );

    \I__929\ : InMux
    port map (
            O => \N__4750\,
            I => \N__4732\
        );

    \I__928\ : InMux
    port map (
            O => \N__4749\,
            I => \N__4732\
        );

    \I__927\ : InMux
    port map (
            O => \N__4748\,
            I => \N__4729\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__4745\,
            I => \N__4721\
        );

    \I__925\ : InMux
    port map (
            O => \N__4744\,
            I => \N__4714\
        );

    \I__924\ : InMux
    port map (
            O => \N__4743\,
            I => \N__4714\
        );

    \I__923\ : InMux
    port map (
            O => \N__4742\,
            I => \N__4714\
        );

    \I__922\ : InMux
    port map (
            O => \N__4741\,
            I => \N__4711\
        );

    \I__921\ : InMux
    port map (
            O => \N__4740\,
            I => \N__4708\
        );

    \I__920\ : InMux
    port map (
            O => \N__4739\,
            I => \N__4703\
        );

    \I__919\ : InMux
    port map (
            O => \N__4738\,
            I => \N__4703\
        );

    \I__918\ : InMux
    port map (
            O => \N__4737\,
            I => \N__4700\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__4732\,
            I => \N__4695\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4729\,
            I => \N__4695\
        );

    \I__915\ : InMux
    port map (
            O => \N__4728\,
            I => \N__4688\
        );

    \I__914\ : InMux
    port map (
            O => \N__4727\,
            I => \N__4688\
        );

    \I__913\ : InMux
    port map (
            O => \N__4726\,
            I => \N__4688\
        );

    \I__912\ : InMux
    port map (
            O => \N__4725\,
            I => \N__4685\
        );

    \I__911\ : InMux
    port map (
            O => \N__4724\,
            I => \N__4682\
        );

    \I__910\ : Span4Mux_h
    port map (
            O => \N__4721\,
            I => \N__4677\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__4714\,
            I => \N__4677\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4711\,
            I => \N__4674\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__4708\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__4703\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__4700\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__904\ : Odrv4
    port map (
            O => \N__4695\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4688\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__4685\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4682\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__900\ : Odrv4
    port map (
            O => \N__4677\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__899\ : Odrv4
    port map (
            O => \N__4674\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__898\ : InMux
    port map (
            O => \N__4655\,
            I => \N__4638\
        );

    \I__897\ : InMux
    port map (
            O => \N__4654\,
            I => \N__4635\
        );

    \I__896\ : InMux
    port map (
            O => \N__4653\,
            I => \N__4630\
        );

    \I__895\ : InMux
    port map (
            O => \N__4652\,
            I => \N__4630\
        );

    \I__894\ : InMux
    port map (
            O => \N__4651\,
            I => \N__4627\
        );

    \I__893\ : InMux
    port map (
            O => \N__4650\,
            I => \N__4622\
        );

    \I__892\ : InMux
    port map (
            O => \N__4649\,
            I => \N__4622\
        );

    \I__891\ : InMux
    port map (
            O => \N__4648\,
            I => \N__4619\
        );

    \I__890\ : InMux
    port map (
            O => \N__4647\,
            I => \N__4616\
        );

    \I__889\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4611\
        );

    \I__888\ : InMux
    port map (
            O => \N__4645\,
            I => \N__4611\
        );

    \I__887\ : InMux
    port map (
            O => \N__4644\,
            I => \N__4606\
        );

    \I__886\ : InMux
    port map (
            O => \N__4643\,
            I => \N__4606\
        );

    \I__885\ : InMux
    port map (
            O => \N__4642\,
            I => \N__4594\
        );

    \I__884\ : InMux
    port map (
            O => \N__4641\,
            I => \N__4594\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__4638\,
            I => \N__4589\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__4635\,
            I => \N__4589\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__4630\,
            I => \N__4578\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4627\,
            I => \N__4578\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__4622\,
            I => \N__4578\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__4619\,
            I => \N__4578\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__4616\,
            I => \N__4578\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__4611\,
            I => \N__4574\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4606\,
            I => \N__4571\
        );

    \I__874\ : InMux
    port map (
            O => \N__4605\,
            I => \N__4564\
        );

    \I__873\ : InMux
    port map (
            O => \N__4604\,
            I => \N__4564\
        );

    \I__872\ : InMux
    port map (
            O => \N__4603\,
            I => \N__4564\
        );

    \I__871\ : InMux
    port map (
            O => \N__4602\,
            I => \N__4557\
        );

    \I__870\ : InMux
    port map (
            O => \N__4601\,
            I => \N__4557\
        );

    \I__869\ : InMux
    port map (
            O => \N__4600\,
            I => \N__4557\
        );

    \I__868\ : InMux
    port map (
            O => \N__4599\,
            I => \N__4554\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4594\,
            I => \N__4549\
        );

    \I__866\ : Span4Mux_v
    port map (
            O => \N__4589\,
            I => \N__4544\
        );

    \I__865\ : Span4Mux_v
    port map (
            O => \N__4578\,
            I => \N__4544\
        );

    \I__864\ : InMux
    port map (
            O => \N__4577\,
            I => \N__4541\
        );

    \I__863\ : Span4Mux_s3_h
    port map (
            O => \N__4574\,
            I => \N__4538\
        );

    \I__862\ : Span4Mux_h
    port map (
            O => \N__4571\,
            I => \N__4535\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4564\,
            I => \N__4528\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__4557\,
            I => \N__4528\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__4554\,
            I => \N__4528\
        );

    \I__858\ : InMux
    port map (
            O => \N__4553\,
            I => \N__4523\
        );

    \I__857\ : InMux
    port map (
            O => \N__4552\,
            I => \N__4523\
        );

    \I__856\ : Odrv12
    port map (
            O => \N__4549\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__855\ : Odrv4
    port map (
            O => \N__4544\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__4541\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__853\ : Odrv4
    port map (
            O => \N__4538\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__852\ : Odrv4
    port map (
            O => \N__4535\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__851\ : Odrv4
    port map (
            O => \N__4528\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__4523\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__849\ : InMux
    port map (
            O => \N__4508\,
            I => \N__4504\
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__4507\,
            I => \N__4497\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4504\,
            I => \N__4493\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__4503\,
            I => \N__4490\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__4502\,
            I => \N__4487\
        );

    \I__844\ : InMux
    port map (
            O => \N__4501\,
            I => \N__4484\
        );

    \I__843\ : InMux
    port map (
            O => \N__4500\,
            I => \N__4479\
        );

    \I__842\ : InMux
    port map (
            O => \N__4497\,
            I => \N__4479\
        );

    \I__841\ : CascadeMux
    port map (
            O => \N__4496\,
            I => \N__4472\
        );

    \I__840\ : Span4Mux_h
    port map (
            O => \N__4493\,
            I => \N__4464\
        );

    \I__839\ : InMux
    port map (
            O => \N__4490\,
            I => \N__4459\
        );

    \I__838\ : InMux
    port map (
            O => \N__4487\,
            I => \N__4459\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4484\,
            I => \N__4454\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__4479\,
            I => \N__4454\
        );

    \I__835\ : InMux
    port map (
            O => \N__4478\,
            I => \N__4451\
        );

    \I__834\ : InMux
    port map (
            O => \N__4477\,
            I => \N__4446\
        );

    \I__833\ : InMux
    port map (
            O => \N__4476\,
            I => \N__4446\
        );

    \I__832\ : InMux
    port map (
            O => \N__4475\,
            I => \N__4443\
        );

    \I__831\ : InMux
    port map (
            O => \N__4472\,
            I => \N__4440\
        );

    \I__830\ : InMux
    port map (
            O => \N__4471\,
            I => \N__4437\
        );

    \I__829\ : InMux
    port map (
            O => \N__4470\,
            I => \N__4434\
        );

    \I__828\ : InMux
    port map (
            O => \N__4469\,
            I => \N__4427\
        );

    \I__827\ : InMux
    port map (
            O => \N__4468\,
            I => \N__4427\
        );

    \I__826\ : InMux
    port map (
            O => \N__4467\,
            I => \N__4427\
        );

    \I__825\ : Odrv4
    port map (
            O => \N__4464\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__4459\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__823\ : Odrv4
    port map (
            O => \N__4454\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__4451\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4446\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__4443\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__4440\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__4437\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__4434\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__4427\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__815\ : InMux
    port map (
            O => \N__4406\,
            I => \N__4397\
        );

    \I__814\ : InMux
    port map (
            O => \N__4405\,
            I => \N__4392\
        );

    \I__813\ : InMux
    port map (
            O => \N__4404\,
            I => \N__4392\
        );

    \I__812\ : InMux
    port map (
            O => \N__4403\,
            I => \N__4389\
        );

    \I__811\ : InMux
    port map (
            O => \N__4402\,
            I => \N__4379\
        );

    \I__810\ : InMux
    port map (
            O => \N__4401\,
            I => \N__4379\
        );

    \I__809\ : InMux
    port map (
            O => \N__4400\,
            I => \N__4374\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4397\,
            I => \N__4369\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__4392\,
            I => \N__4369\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__4389\,
            I => \N__4366\
        );

    \I__805\ : InMux
    port map (
            O => \N__4388\,
            I => \N__4363\
        );

    \I__804\ : InMux
    port map (
            O => \N__4387\,
            I => \N__4360\
        );

    \I__803\ : InMux
    port map (
            O => \N__4386\,
            I => \N__4355\
        );

    \I__802\ : InMux
    port map (
            O => \N__4385\,
            I => \N__4355\
        );

    \I__801\ : InMux
    port map (
            O => \N__4384\,
            I => \N__4352\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4379\,
            I => \N__4349\
        );

    \I__799\ : InMux
    port map (
            O => \N__4378\,
            I => \N__4341\
        );

    \I__798\ : InMux
    port map (
            O => \N__4377\,
            I => \N__4338\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__4374\,
            I => \N__4335\
        );

    \I__796\ : Span4Mux_v
    port map (
            O => \N__4369\,
            I => \N__4328\
        );

    \I__795\ : Span4Mux_v
    port map (
            O => \N__4366\,
            I => \N__4328\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__4363\,
            I => \N__4328\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__4360\,
            I => \N__4323\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__4355\,
            I => \N__4323\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__4352\,
            I => \N__4318\
        );

    \I__790\ : Span4Mux_h
    port map (
            O => \N__4349\,
            I => \N__4318\
        );

    \I__789\ : InMux
    port map (
            O => \N__4348\,
            I => \N__4311\
        );

    \I__788\ : InMux
    port map (
            O => \N__4347\,
            I => \N__4311\
        );

    \I__787\ : InMux
    port map (
            O => \N__4346\,
            I => \N__4311\
        );

    \I__786\ : InMux
    port map (
            O => \N__4345\,
            I => \N__4306\
        );

    \I__785\ : InMux
    port map (
            O => \N__4344\,
            I => \N__4306\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__4341\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__4338\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__782\ : Odrv4
    port map (
            O => \N__4335\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__781\ : Odrv4
    port map (
            O => \N__4328\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__780\ : Odrv4
    port map (
            O => \N__4323\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__779\ : Odrv4
    port map (
            O => \N__4318\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__4311\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__4306\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__776\ : InMux
    port map (
            O => \N__4289\,
            I => \N__4286\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__4286\,
            I => \U400_SDRAM.N_30\
        );

    \I__774\ : InMux
    port map (
            O => \N__4283\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_0\
        );

    \I__773\ : InMux
    port map (
            O => \N__4280\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_1\
        );

    \I__772\ : CascadeMux
    port map (
            O => \N__4277\,
            I => \N__4274\
        );

    \I__771\ : InMux
    port map (
            O => \N__4274\,
            I => \N__4271\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__4271\,
            I => \U400_SDRAM.SDRAM_COUNTER_s_3\
        );

    \I__769\ : InMux
    port map (
            O => \N__4268\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_2\
        );

    \I__768\ : InMux
    port map (
            O => \N__4265\,
            I => \N__4261\
        );

    \I__767\ : InMux
    port map (
            O => \N__4264\,
            I => \N__4258\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__4261\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__4258\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__764\ : InMux
    port map (
            O => \N__4253\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_3\
        );

    \I__763\ : InMux
    port map (
            O => \N__4250\,
            I => \N__4245\
        );

    \I__762\ : InMux
    port map (
            O => \N__4249\,
            I => \N__4242\
        );

    \I__761\ : InMux
    port map (
            O => \N__4248\,
            I => \N__4239\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__4245\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__4242\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__4239\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__757\ : InMux
    port map (
            O => \N__4232\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_4\
        );

    \I__756\ : InMux
    port map (
            O => \N__4229\,
            I => \N__4224\
        );

    \I__755\ : InMux
    port map (
            O => \N__4228\,
            I => \N__4221\
        );

    \I__754\ : InMux
    port map (
            O => \N__4227\,
            I => \N__4218\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__4224\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__4221\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4218\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__750\ : InMux
    port map (
            O => \N__4211\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_5\
        );

    \I__749\ : InMux
    port map (
            O => \N__4208\,
            I => \N__4205\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__4205\,
            I => \N__4195\
        );

    \I__747\ : InMux
    port map (
            O => \N__4204\,
            I => \N__4192\
        );

    \I__746\ : InMux
    port map (
            O => \N__4203\,
            I => \N__4183\
        );

    \I__745\ : InMux
    port map (
            O => \N__4202\,
            I => \N__4183\
        );

    \I__744\ : InMux
    port map (
            O => \N__4201\,
            I => \N__4183\
        );

    \I__743\ : InMux
    port map (
            O => \N__4200\,
            I => \N__4183\
        );

    \I__742\ : InMux
    port map (
            O => \N__4199\,
            I => \N__4178\
        );

    \I__741\ : InMux
    port map (
            O => \N__4198\,
            I => \N__4178\
        );

    \I__740\ : Odrv4
    port map (
            O => \N__4195\,
            I => \U400_SDRAM.N_29\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__4192\,
            I => \U400_SDRAM.N_29\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__4183\,
            I => \U400_SDRAM.N_29\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__4178\,
            I => \U400_SDRAM.N_29\
        );

    \I__736\ : InMux
    port map (
            O => \N__4169\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_6\
        );

    \I__735\ : CascadeMux
    port map (
            O => \N__4166\,
            I => \N__4162\
        );

    \I__734\ : InMux
    port map (
            O => \N__4165\,
            I => \N__4159\
        );

    \I__733\ : InMux
    port map (
            O => \N__4162\,
            I => \N__4156\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__4159\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__4156\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__730\ : CEMux
    port map (
            O => \N__4151\,
            I => \N__4146\
        );

    \I__729\ : CEMux
    port map (
            O => \N__4150\,
            I => \N__4143\
        );

    \I__728\ : CEMux
    port map (
            O => \N__4149\,
            I => \N__4140\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__4146\,
            I => \N__4137\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__4143\,
            I => \N__4134\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__4140\,
            I => \N__4131\
        );

    \I__724\ : Span4Mux_v
    port map (
            O => \N__4137\,
            I => \N__4124\
        );

    \I__723\ : Span4Mux_h
    port map (
            O => \N__4134\,
            I => \N__4124\
        );

    \I__722\ : Span4Mux_h
    port map (
            O => \N__4131\,
            I => \N__4124\
        );

    \I__721\ : Odrv4
    port map (
            O => \N__4124\,
            I => \U400_SDRAM.SDRAM_COUNTERe_0_i\
        );

    \I__720\ : InMux
    port map (
            O => \N__4121\,
            I => \N__4117\
        );

    \I__719\ : InMux
    port map (
            O => \N__4120\,
            I => \N__4114\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__4117\,
            I => \U400_SDRAM.N_336_1\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__4114\,
            I => \U400_SDRAM.N_336_1\
        );

    \I__716\ : CascadeMux
    port map (
            O => \N__4109\,
            I => \U400_SDRAM.N_56_cascade_\
        );

    \I__715\ : CascadeMux
    port map (
            O => \N__4106\,
            I => \N__4103\
        );

    \I__714\ : InMux
    port map (
            O => \N__4103\,
            I => \N__4100\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__4100\,
            I => \N__4097\
        );

    \I__712\ : Span4Mux_h
    port map (
            O => \N__4097\,
            I => \N__4094\
        );

    \I__711\ : Odrv4
    port map (
            O => \N__4094\,
            I => \U400_SDRAM.TACK_7_iv_i_0\
        );

    \I__710\ : CascadeMux
    port map (
            O => \N__4091\,
            I => \U400_SDRAM.N_8_cascade_\
        );

    \I__709\ : InMux
    port map (
            O => \N__4088\,
            I => \N__4085\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__4085\,
            I => \U400_SDRAM.un1_SDRAM_COUNTER59_4_i_1\
        );

    \I__707\ : CascadeMux
    port map (
            O => \N__4082\,
            I => \U400_SDRAM.N_15_cascade_\
        );

    \I__706\ : InMux
    port map (
            O => \N__4079\,
            I => \N__4076\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__4076\,
            I => \N__4073\
        );

    \I__704\ : Odrv4
    port map (
            O => \N__4073\,
            I => \U400_SDRAM.N_87\
        );

    \I__703\ : InMux
    port map (
            O => \N__4070\,
            I => \N__4067\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__4067\,
            I => \U400_SDRAM.N_25\
        );

    \I__701\ : InMux
    port map (
            O => \N__4064\,
            I => \N__4061\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__4061\,
            I => \U400_SDRAM.N_84\
        );

    \I__699\ : InMux
    port map (
            O => \N__4058\,
            I => \N__4055\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__4055\,
            I => \U400_SDRAM.N_88\
        );

    \I__697\ : InMux
    port map (
            O => \N__4052\,
            I => \N__4047\
        );

    \I__696\ : InMux
    port map (
            O => \N__4051\,
            I => \N__4044\
        );

    \I__695\ : InMux
    port map (
            O => \N__4050\,
            I => \N__4041\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__4047\,
            I => \U400_SDRAM.N_48\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__4044\,
            I => \U400_SDRAM.N_48\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__4041\,
            I => \U400_SDRAM.N_48\
        );

    \I__691\ : CascadeMux
    port map (
            O => \N__4034\,
            I => \N__4031\
        );

    \I__690\ : InMux
    port map (
            O => \N__4031\,
            I => \N__4028\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__4028\,
            I => \N__4025\
        );

    \I__688\ : Span4Mux_h
    port map (
            O => \N__4025\,
            I => \N__4022\
        );

    \I__687\ : Odrv4
    port map (
            O => \N__4022\,
            I => \U400_SDRAM.SDRAM_COUNTER_s_1\
        );

    \I__686\ : CascadeMux
    port map (
            O => \N__4019\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_3_cascade_\
        );

    \I__685\ : InMux
    port map (
            O => \N__4016\,
            I => \N__4009\
        );

    \I__684\ : InMux
    port map (
            O => \N__4015\,
            I => \N__4009\
        );

    \I__683\ : InMux
    port map (
            O => \N__4014\,
            I => \N__4006\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__4009\,
            I => \U400_SDRAM.N_38\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__4006\,
            I => \U400_SDRAM.N_38\
        );

    \I__680\ : CascadeMux
    port map (
            O => \N__4001\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_a2_2_0_cascade_\
        );

    \I__679\ : InMux
    port map (
            O => \N__3998\,
            I => \N__3995\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__3995\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_2\
        );

    \I__677\ : InMux
    port map (
            O => \N__3992\,
            I => \N__3989\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__3989\,
            I => \N__3986\
        );

    \I__675\ : Odrv12
    port map (
            O => \N__3986\,
            I => \A_c_5\
        );

    \I__674\ : InMux
    port map (
            O => \N__3983\,
            I => \N__3980\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__3980\,
            I => \N__3977\
        );

    \I__672\ : Span4Mux_v
    port map (
            O => \N__3977\,
            I => \N__3974\
        );

    \I__671\ : Span4Mux_v
    port map (
            O => \N__3974\,
            I => \N__3971\
        );

    \I__670\ : Sp12to4
    port map (
            O => \N__3971\,
            I => \N__3968\
        );

    \I__669\ : Odrv12
    port map (
            O => \N__3968\,
            I => \A_c_16\
        );

    \I__668\ : IoInMux
    port map (
            O => \N__3965\,
            I => \N__3962\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__3962\,
            I => \N__3959\
        );

    \I__666\ : Span12Mux_s3_v
    port map (
            O => \N__3959\,
            I => \N__3956\
        );

    \I__665\ : Odrv12
    port map (
            O => \N__3956\,
            I => \MA_c_3\
        );

    \I__664\ : CascadeMux
    port map (
            O => \N__3953\,
            I => \N__3950\
        );

    \I__663\ : InMux
    port map (
            O => \N__3950\,
            I => \N__3947\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__3947\,
            I => \N__3944\
        );

    \I__661\ : Span4Mux_h
    port map (
            O => \N__3944\,
            I => \N__3941\
        );

    \I__660\ : Sp12to4
    port map (
            O => \N__3941\,
            I => \N__3938\
        );

    \I__659\ : Span12Mux_v
    port map (
            O => \N__3938\,
            I => \N__3935\
        );

    \I__658\ : Odrv12
    port map (
            O => \N__3935\,
            I => \A_c_26\
        );

    \I__657\ : IoInMux
    port map (
            O => \N__3932\,
            I => \N__3929\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__3929\,
            I => \N__3926\
        );

    \I__655\ : Span4Mux_s0_v
    port map (
            O => \N__3926\,
            I => \N__3923\
        );

    \I__654\ : Odrv4
    port map (
            O => \N__3923\,
            I => \MA_c_12\
        );

    \I__653\ : InMux
    port map (
            O => \N__3920\,
            I => \N__3917\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__3917\,
            I => \N__3914\
        );

    \I__651\ : Span4Mux_v
    port map (
            O => \N__3914\,
            I => \N__3911\
        );

    \I__650\ : Span4Mux_h
    port map (
            O => \N__3911\,
            I => \N__3908\
        );

    \I__649\ : Odrv4
    port map (
            O => \N__3908\,
            I => \A_c_7\
        );

    \I__648\ : InMux
    port map (
            O => \N__3905\,
            I => \N__3902\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__3902\,
            I => \N__3899\
        );

    \I__646\ : Odrv12
    port map (
            O => \N__3899\,
            I => \U400_SDRAM.MA_5_iv_0_5\
        );

    \I__645\ : IoInMux
    port map (
            O => \N__3896\,
            I => \N__3893\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3893\,
            I => \N__3890\
        );

    \I__643\ : Span4Mux_s3_v
    port map (
            O => \N__3890\,
            I => \N__3887\
        );

    \I__642\ : Odrv4
    port map (
            O => \N__3887\,
            I => \MA_c_5\
        );

    \I__641\ : CascadeMux
    port map (
            O => \N__3884\,
            I => \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_a2_0_0_cascade_\
        );

    \I__640\ : CascadeMux
    port map (
            O => \N__3881\,
            I => \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_1_cascade_\
        );

    \I__639\ : InMux
    port map (
            O => \N__3878\,
            I => \N__3875\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__3875\,
            I => \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_3\
        );

    \I__637\ : CascadeMux
    port map (
            O => \N__3872\,
            I => \N__3869\
        );

    \I__636\ : InMux
    port map (
            O => \N__3869\,
            I => \N__3866\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__3866\,
            I => \U400_SDRAM.N_60\
        );

    \I__634\ : CascadeMux
    port map (
            O => \N__3863\,
            I => \U400_SDRAM.N_97_cascade_\
        );

    \I__633\ : InMux
    port map (
            O => \N__3860\,
            I => \N__3857\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__3857\,
            I => \N__3853\
        );

    \I__631\ : InMux
    port map (
            O => \N__3856\,
            I => \N__3850\
        );

    \I__630\ : Odrv4
    port map (
            O => \N__3853\,
            I => \U400_SDRAM.N_20\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__3850\,
            I => \U400_SDRAM.N_20\
        );

    \I__628\ : CascadeMux
    port map (
            O => \N__3845\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_1_66_i_0_2_cascade_\
        );

    \I__627\ : CascadeMux
    port map (
            O => \N__3842\,
            I => \N__3839\
        );

    \I__626\ : InMux
    port map (
            O => \N__3839\,
            I => \N__3836\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3836\,
            I => \N__3833\
        );

    \I__624\ : Span4Mux_v
    port map (
            O => \N__3833\,
            I => \N__3830\
        );

    \I__623\ : Span4Mux_h
    port map (
            O => \N__3830\,
            I => \N__3827\
        );

    \I__622\ : Odrv4
    port map (
            O => \N__3827\,
            I => \A_c_18\
        );

    \I__621\ : InMux
    port map (
            O => \N__3824\,
            I => \N__3820\
        );

    \I__620\ : InMux
    port map (
            O => \N__3823\,
            I => \N__3817\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__3820\,
            I => \N__3813\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__3817\,
            I => \N__3810\
        );

    \I__617\ : InMux
    port map (
            O => \N__3816\,
            I => \N__3807\
        );

    \I__616\ : Odrv4
    port map (
            O => \N__3813\,
            I => \U400_SDRAM.N_11\
        );

    \I__615\ : Odrv4
    port map (
            O => \N__3810\,
            I => \U400_SDRAM.N_11\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__3807\,
            I => \U400_SDRAM.N_11\
        );

    \I__613\ : InMux
    port map (
            O => \N__3800\,
            I => \N__3797\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__3797\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_1\
        );

    \I__611\ : CascadeMux
    port map (
            O => \N__3794\,
            I => \U400_SDRAM.N_44_cascade_\
        );

    \I__610\ : InMux
    port map (
            O => \N__3791\,
            I => \N__3784\
        );

    \I__609\ : InMux
    port map (
            O => \N__3790\,
            I => \N__3784\
        );

    \I__608\ : InMux
    port map (
            O => \N__3789\,
            I => \N__3781\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__3784\,
            I => \N__3777\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3781\,
            I => \N__3773\
        );

    \I__605\ : InMux
    port map (
            O => \N__3780\,
            I => \N__3770\
        );

    \I__604\ : Span4Mux_h
    port map (
            O => \N__3777\,
            I => \N__3767\
        );

    \I__603\ : InMux
    port map (
            O => \N__3776\,
            I => \N__3764\
        );

    \I__602\ : Odrv4
    port map (
            O => \N__3773\,
            I => \U400_SDRAM.N_108\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3770\,
            I => \U400_SDRAM.N_108\
        );

    \I__600\ : Odrv4
    port map (
            O => \N__3767\,
            I => \U400_SDRAM.N_108\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3764\,
            I => \U400_SDRAM.N_108\
        );

    \I__598\ : CascadeMux
    port map (
            O => \N__3755\,
            I => \U400_SDRAM.N_108_cascade_\
        );

    \I__597\ : InMux
    port map (
            O => \N__3752\,
            I => \N__3749\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3749\,
            I => \N__3746\
        );

    \I__595\ : Span4Mux_h
    port map (
            O => \N__3746\,
            I => \N__3742\
        );

    \I__594\ : InMux
    port map (
            O => \N__3745\,
            I => \N__3739\
        );

    \I__593\ : Odrv4
    port map (
            O => \N__3742\,
            I => \U400_SDRAM.N_109\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__3739\,
            I => \U400_SDRAM.N_109\
        );

    \I__591\ : InMux
    port map (
            O => \N__3734\,
            I => \N__3727\
        );

    \I__590\ : InMux
    port map (
            O => \N__3733\,
            I => \N__3727\
        );

    \I__589\ : InMux
    port map (
            O => \N__3732\,
            I => \N__3724\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3727\,
            I => \N__3721\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__3724\,
            I => \U400_SDRAM.N_52\
        );

    \I__586\ : Odrv4
    port map (
            O => \N__3721\,
            I => \U400_SDRAM.N_52\
        );

    \I__585\ : InMux
    port map (
            O => \N__3716\,
            I => \N__3713\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__3713\,
            I => \N__3710\
        );

    \I__583\ : Span4Mux_h
    port map (
            O => \N__3710\,
            I => \N__3707\
        );

    \I__582\ : Span4Mux_s1_h
    port map (
            O => \N__3707\,
            I => \N__3704\
        );

    \I__581\ : Odrv4
    port map (
            O => \N__3704\,
            I => \U400_SDRAM.SDRAM_COUNTER_s_0\
        );

    \I__580\ : InMux
    port map (
            O => \N__3701\,
            I => \N__3698\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__3698\,
            I => \N__3695\
        );

    \I__578\ : Odrv4
    port map (
            O => \N__3695\,
            I => \U400_SDRAM.N_86\
        );

    \I__577\ : CascadeMux
    port map (
            O => \N__3692\,
            I => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_1_0_cascade_\
        );

    \I__576\ : InMux
    port map (
            O => \N__3689\,
            I => \N__3684\
        );

    \I__575\ : InMux
    port map (
            O => \N__3688\,
            I => \N__3681\
        );

    \I__574\ : InMux
    port map (
            O => \N__3687\,
            I => \N__3678\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__3684\,
            I => \U400_SDRAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3681\,
            I => \U400_SDRAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3678\,
            I => \U400_SDRAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__570\ : InMux
    port map (
            O => \N__3671\,
            I => \N__3668\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__3668\,
            I => \N__3664\
        );

    \I__568\ : InMux
    port map (
            O => \N__3667\,
            I => \N__3661\
        );

    \I__567\ : Span4Mux_v
    port map (
            O => \N__3664\,
            I => \N__3656\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__3661\,
            I => \N__3656\
        );

    \I__565\ : Span4Mux_h
    port map (
            O => \N__3656\,
            I => \N__3652\
        );

    \I__564\ : InMux
    port map (
            O => \N__3655\,
            I => \N__3649\
        );

    \I__563\ : Odrv4
    port map (
            O => \N__3652\,
            I => \U400_SDRAM.N_118\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3649\,
            I => \U400_SDRAM.N_118\
        );

    \I__561\ : InMux
    port map (
            O => \N__3644\,
            I => \N__3641\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3641\,
            I => \U400_SDRAM.SDRAM_COUNTER_3_sqmuxa_0_a3_0_a2_0\
        );

    \I__559\ : CascadeMux
    port map (
            O => \N__3638\,
            I => \U400_SDRAM.N_46_cascade_\
        );

    \I__558\ : InMux
    port map (
            O => \N__3635\,
            I => \N__3632\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3632\,
            I => \N__3628\
        );

    \I__556\ : InMux
    port map (
            O => \N__3631\,
            I => \N__3622\
        );

    \I__555\ : Span4Mux_s2_v
    port map (
            O => \N__3628\,
            I => \N__3619\
        );

    \I__554\ : InMux
    port map (
            O => \N__3627\,
            I => \N__3614\
        );

    \I__553\ : InMux
    port map (
            O => \N__3626\,
            I => \N__3614\
        );

    \I__552\ : InMux
    port map (
            O => \N__3625\,
            I => \N__3607\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3622\,
            I => \N__3600\
        );

    \I__550\ : Span4Mux_v
    port map (
            O => \N__3619\,
            I => \N__3600\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3614\,
            I => \N__3600\
        );

    \I__548\ : InMux
    port map (
            O => \N__3613\,
            I => \N__3591\
        );

    \I__547\ : InMux
    port map (
            O => \N__3612\,
            I => \N__3591\
        );

    \I__546\ : InMux
    port map (
            O => \N__3611\,
            I => \N__3591\
        );

    \I__545\ : InMux
    port map (
            O => \N__3610\,
            I => \N__3591\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__3607\,
            I => \U400_SDRAM.RAM_CYCLE_STARTZ0\
        );

    \I__543\ : Odrv4
    port map (
            O => \N__3600\,
            I => \U400_SDRAM.RAM_CYCLE_STARTZ0\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__3591\,
            I => \U400_SDRAM.RAM_CYCLE_STARTZ0\
        );

    \I__541\ : InMux
    port map (
            O => \N__3584\,
            I => \N__3581\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__3581\,
            I => \U400_SDRAM.SDRAM_COUNTER_4_sqmuxa_0_a3_0\
        );

    \I__539\ : InMux
    port map (
            O => \N__3578\,
            I => \N__3575\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3575\,
            I => \N__3572\
        );

    \I__537\ : Span4Mux_v
    port map (
            O => \N__3572\,
            I => \N__3569\
        );

    \I__536\ : Span4Mux_h
    port map (
            O => \N__3569\,
            I => \N__3566\
        );

    \I__535\ : Odrv4
    port map (
            O => \N__3566\,
            I => \RnW_c\
        );

    \I__534\ : InMux
    port map (
            O => \N__3563\,
            I => \N__3560\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3560\,
            I => \N__3554\
        );

    \I__532\ : InMux
    port map (
            O => \N__3559\,
            I => \N__3549\
        );

    \I__531\ : InMux
    port map (
            O => \N__3558\,
            I => \N__3549\
        );

    \I__530\ : InMux
    port map (
            O => \N__3557\,
            I => \N__3546\
        );

    \I__529\ : Odrv4
    port map (
            O => \N__3554\,
            I => \U400_SDRAM.N_113\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__3549\,
            I => \U400_SDRAM.N_113\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3546\,
            I => \U400_SDRAM.N_113\
        );

    \I__526\ : InMux
    port map (
            O => \N__3539\,
            I => \N__3536\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3536\,
            I => \U400_SDRAM.N_63\
        );

    \I__524\ : CascadeMux
    port map (
            O => \N__3533\,
            I => \U400_SDRAM.N_20_cascade_\
        );

    \I__523\ : InMux
    port map (
            O => \N__3530\,
            I => \N__3527\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__3527\,
            I => \N__3524\
        );

    \I__521\ : Odrv12
    port map (
            O => \N__3524\,
            I => \U400_SDRAM.N_35\
        );

    \I__520\ : InMux
    port map (
            O => \N__3521\,
            I => \N__3518\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3518\,
            I => \N__3514\
        );

    \I__518\ : InMux
    port map (
            O => \N__3517\,
            I => \N__3511\
        );

    \I__517\ : Odrv12
    port map (
            O => \N__3514\,
            I => \U400_SDRAM.N_39\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__3511\,
            I => \U400_SDRAM.N_39\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__3506\,
            I => \U400_SDRAM.N_35_cascade_\
        );

    \I__514\ : CascadeMux
    port map (
            O => \N__3503\,
            I => \U400_SDRAM.N_12_cascade_\
        );

    \I__513\ : CascadeMux
    port map (
            O => \N__3500\,
            I => \U400_SDRAM.N_91_cascade_\
        );

    \I__512\ : InMux
    port map (
            O => \N__3497\,
            I => \N__3494\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3494\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_0_103_i_i_a3_0_0\
        );

    \I__510\ : InMux
    port map (
            O => \N__3491\,
            I => \N__3488\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3488\,
            I => \U400_SDRAM.N_89\
        );

    \I__508\ : CascadeMux
    port map (
            O => \N__3485\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_0_103_i_i_0_cascade_\
        );

    \I__507\ : InMux
    port map (
            O => \N__3482\,
            I => \N__3479\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__3479\,
            I => \N__3476\
        );

    \I__505\ : Span4Mux_v
    port map (
            O => \N__3476\,
            I => \N__3473\
        );

    \I__504\ : Span4Mux_h
    port map (
            O => \N__3473\,
            I => \N__3470\
        );

    \I__503\ : Odrv4
    port map (
            O => \N__3470\,
            I => \A_c_8\
        );

    \I__502\ : CascadeMux
    port map (
            O => \N__3467\,
            I => \N__3464\
        );

    \I__501\ : InMux
    port map (
            O => \N__3464\,
            I => \N__3461\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__3461\,
            I => \N__3458\
        );

    \I__499\ : Span4Mux_v
    port map (
            O => \N__3458\,
            I => \N__3455\
        );

    \I__498\ : Span4Mux_v
    port map (
            O => \N__3455\,
            I => \N__3452\
        );

    \I__497\ : Odrv4
    port map (
            O => \N__3452\,
            I => \A_c_19\
        );

    \I__496\ : IoInMux
    port map (
            O => \N__3449\,
            I => \N__3446\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__3446\,
            I => \N__3443\
        );

    \I__494\ : Odrv12
    port map (
            O => \N__3443\,
            I => \MA_c_6\
        );

    \I__493\ : InMux
    port map (
            O => \N__3440\,
            I => \N__3437\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3437\,
            I => \N__3434\
        );

    \I__491\ : Odrv12
    port map (
            O => \N__3434\,
            I => \A_c_6\
        );

    \I__490\ : CascadeMux
    port map (
            O => \N__3431\,
            I => \N__3428\
        );

    \I__489\ : InMux
    port map (
            O => \N__3428\,
            I => \N__3425\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__3425\,
            I => \N__3422\
        );

    \I__487\ : Span12Mux_s8_v
    port map (
            O => \N__3422\,
            I => \N__3419\
        );

    \I__486\ : Odrv12
    port map (
            O => \N__3419\,
            I => \A_c_17\
        );

    \I__485\ : IoInMux
    port map (
            O => \N__3416\,
            I => \N__3413\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3413\,
            I => \N__3410\
        );

    \I__483\ : Span4Mux_s3_v
    port map (
            O => \N__3410\,
            I => \N__3407\
        );

    \I__482\ : Odrv4
    port map (
            O => \N__3407\,
            I => \MA_c_4\
        );

    \I__481\ : InMux
    port map (
            O => \N__3404\,
            I => \N__3401\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3401\,
            I => \N__3398\
        );

    \I__479\ : Span4Mux_v
    port map (
            O => \N__3398\,
            I => \N__3395\
        );

    \I__478\ : Span4Mux_v
    port map (
            O => \N__3395\,
            I => \N__3392\
        );

    \I__477\ : Span4Mux_v
    port map (
            O => \N__3392\,
            I => \N__3389\
        );

    \I__476\ : Odrv4
    port map (
            O => \N__3389\,
            I => \A_c_20\
        );

    \I__475\ : CascadeMux
    port map (
            O => \N__3386\,
            I => \N__3383\
        );

    \I__474\ : InMux
    port map (
            O => \N__3383\,
            I => \N__3380\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__3380\,
            I => \N__3377\
        );

    \I__472\ : Span12Mux_s4_v
    port map (
            O => \N__3377\,
            I => \N__3374\
        );

    \I__471\ : Odrv12
    port map (
            O => \N__3374\,
            I => \A_c_9\
        );

    \I__470\ : IoInMux
    port map (
            O => \N__3371\,
            I => \N__3368\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3368\,
            I => \N__3365\
        );

    \I__468\ : Odrv12
    port map (
            O => \N__3365\,
            I => \MA_c_7\
        );

    \I__467\ : CascadeMux
    port map (
            O => \N__3362\,
            I => \U400_SDRAM.N_113_cascade_\
        );

    \I__466\ : CascadeMux
    port map (
            O => \N__3359\,
            I => \U400_SDRAM.N_39_cascade_\
        );

    \I__465\ : InMux
    port map (
            O => \N__3356\,
            I => \N__3353\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__3353\,
            I => \N__3350\
        );

    \I__463\ : Odrv4
    port map (
            O => \N__3350\,
            I => \U400_SDRAM.SDRAM_COUNTER_1_sqmuxa_i_0_1\
        );

    \I__462\ : InMux
    port map (
            O => \N__3347\,
            I => \N__3344\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__3344\,
            I => \N__3341\
        );

    \I__460\ : Span4Mux_s2_h
    port map (
            O => \N__3341\,
            I => \N__3338\
        );

    \I__459\ : Odrv4
    port map (
            O => \N__3338\,
            I => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_a2_1_0_0\
        );

    \I__458\ : CascadeMux
    port map (
            O => \N__3335\,
            I => \U400_SDRAM.N_78_cascade_\
        );

    \I__457\ : InMux
    port map (
            O => \N__3332\,
            I => \N__3326\
        );

    \I__456\ : InMux
    port map (
            O => \N__3331\,
            I => \N__3326\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__3326\,
            I => \N__3321\
        );

    \I__454\ : CascadeMux
    port map (
            O => \N__3325\,
            I => \N__3318\
        );

    \I__453\ : InMux
    port map (
            O => \N__3324\,
            I => \N__3314\
        );

    \I__452\ : Span4Mux_v
    port map (
            O => \N__3321\,
            I => \N__3311\
        );

    \I__451\ : InMux
    port map (
            O => \N__3318\,
            I => \N__3306\
        );

    \I__450\ : InMux
    port map (
            O => \N__3317\,
            I => \N__3306\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__3314\,
            I => \U400_SDRAM.N_337_1\
        );

    \I__448\ : Odrv4
    port map (
            O => \N__3311\,
            I => \U400_SDRAM.N_337_1\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__3306\,
            I => \U400_SDRAM.N_337_1\
        );

    \I__446\ : IoInMux
    port map (
            O => \N__3299\,
            I => \N__3296\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__3296\,
            I => \N__3293\
        );

    \I__444\ : Odrv4
    port map (
            O => \N__3293\,
            I => \RASn_c\
        );

    \I__443\ : CascadeMux
    port map (
            O => \N__3290\,
            I => \N__3287\
        );

    \I__442\ : InMux
    port map (
            O => \N__3287\,
            I => \N__3284\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__3284\,
            I => \N__3280\
        );

    \I__440\ : InMux
    port map (
            O => \N__3283\,
            I => \N__3277\
        );

    \I__439\ : Odrv12
    port map (
            O => \N__3280\,
            I => \U400_SDRAM.CS0_ENZ0\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__3277\,
            I => \U400_SDRAM.CS0_ENZ0\
        );

    \I__437\ : IoInMux
    port map (
            O => \N__3272\,
            I => \N__3269\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__3269\,
            I => \N__3266\
        );

    \I__435\ : Odrv4
    port map (
            O => \N__3266\,
            I => \CS0n_c\
        );

    \I__434\ : InMux
    port map (
            O => \N__3263\,
            I => \N__3260\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__3260\,
            I => \N__3257\
        );

    \I__432\ : Span4Mux_h
    port map (
            O => \N__3257\,
            I => \N__3254\
        );

    \I__431\ : Odrv4
    port map (
            O => \N__3254\,
            I => \A_c_31\
        );

    \I__430\ : InMux
    port map (
            O => \N__3251\,
            I => \N__3248\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__3248\,
            I => \N__3245\
        );

    \I__428\ : Span4Mux_h
    port map (
            O => \N__3245\,
            I => \N__3242\
        );

    \I__427\ : Odrv4
    port map (
            O => \N__3242\,
            I => \A_c_30\
        );

    \I__426\ : InMux
    port map (
            O => \N__3239\,
            I => \N__3236\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__3236\,
            I => \N__3233\
        );

    \I__424\ : Span4Mux_h
    port map (
            O => \N__3233\,
            I => \N__3230\
        );

    \I__423\ : Odrv4
    port map (
            O => \N__3230\,
            I => \A_c_29\
        );

    \I__422\ : InMux
    port map (
            O => \N__3227\,
            I => \N__3224\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3224\,
            I => \A_c_28\
        );

    \I__420\ : InMux
    port map (
            O => \N__3221\,
            I => \N__3218\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__3218\,
            I => \N__3215\
        );

    \I__418\ : Span12Mux_s6_v
    port map (
            O => \N__3215\,
            I => \N__3212\
        );

    \I__417\ : Odrv12
    port map (
            O => \N__3212\,
            I => \TSn_c\
        );

    \I__416\ : InMux
    port map (
            O => \N__3209\,
            I => \N__3206\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__3206\,
            I => \N__3203\
        );

    \I__414\ : Span4Mux_v
    port map (
            O => \N__3203\,
            I => \N__3200\
        );

    \I__413\ : Odrv4
    port map (
            O => \N__3200\,
            I => \U400_SDRAM.N_101\
        );

    \I__412\ : InMux
    port map (
            O => \N__3197\,
            I => \N__3193\
        );

    \I__411\ : InMux
    port map (
            O => \N__3196\,
            I => \N__3190\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__3193\,
            I => \N__3185\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__3190\,
            I => \N__3185\
        );

    \I__408\ : Odrv4
    port map (
            O => \N__3185\,
            I => \U400_ADDRESS_DECODE_RAM_SPACE_i_o3_2\
        );

    \I__407\ : CascadeMux
    port map (
            O => \N__3182\,
            I => \N__3178\
        );

    \I__406\ : InMux
    port map (
            O => \N__3181\,
            I => \N__3173\
        );

    \I__405\ : InMux
    port map (
            O => \N__3178\,
            I => \N__3173\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__3173\,
            I => \N__3170\
        );

    \I__403\ : Span12Mux_v
    port map (
            O => \N__3170\,
            I => \N__3167\
        );

    \I__402\ : Odrv12
    port map (
            O => \N__3167\,
            I => \A_c_27\
        );

    \I__401\ : CascadeMux
    port map (
            O => \N__3164\,
            I => \N__3161\
        );

    \I__400\ : InMux
    port map (
            O => \N__3161\,
            I => \N__3155\
        );

    \I__399\ : InMux
    port map (
            O => \N__3160\,
            I => \N__3155\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__3155\,
            I => \N__3152\
        );

    \I__397\ : Odrv4
    port map (
            O => \N__3152\,
            I => \U400_ADDRESS_DECODE_RAM_SPACE_i_o3_1\
        );

    \I__396\ : CascadeMux
    port map (
            O => \N__3149\,
            I => \U400_SDRAM.N_72_cascade_\
        );

    \I__395\ : InMux
    port map (
            O => \N__3146\,
            I => \N__3143\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__3143\,
            I => \U400_SDRAM.N_40\
        );

    \I__393\ : CascadeMux
    port map (
            O => \N__3140\,
            I => \N__3137\
        );

    \I__392\ : InMux
    port map (
            O => \N__3137\,
            I => \N__3131\
        );

    \I__391\ : InMux
    port map (
            O => \N__3136\,
            I => \N__3131\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3131\,
            I => \N__3128\
        );

    \I__389\ : Span4Mux_h
    port map (
            O => \N__3128\,
            I => \N__3125\
        );

    \I__388\ : Span4Mux_v
    port map (
            O => \N__3125\,
            I => \N__3122\
        );

    \I__387\ : Odrv4
    port map (
            O => \N__3122\,
            I => \A_c_23\
        );

    \I__386\ : CascadeMux
    port map (
            O => \N__3119\,
            I => \U400_SDRAM.N_40_cascade_\
        );

    \I__385\ : InMux
    port map (
            O => \N__3116\,
            I => \N__3113\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__3113\,
            I => \U400_SDRAM.CS0_EN_0\
        );

    \I__383\ : CascadeMux
    port map (
            O => \N__3110\,
            I => \N__3105\
        );

    \I__382\ : InMux
    port map (
            O => \N__3109\,
            I => \N__3102\
        );

    \I__381\ : InMux
    port map (
            O => \N__3108\,
            I => \N__3097\
        );

    \I__380\ : InMux
    port map (
            O => \N__3105\,
            I => \N__3097\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__3102\,
            I => \U400_SDRAM.N_115\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__3097\,
            I => \U400_SDRAM.N_115\
        );

    \I__377\ : CascadeMux
    port map (
            O => \N__3092\,
            I => \N__3089\
        );

    \I__376\ : InMux
    port map (
            O => \N__3089\,
            I => \N__3085\
        );

    \I__375\ : InMux
    port map (
            O => \N__3088\,
            I => \N__3082\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__3085\,
            I => \U400_SDRAM.RAM_CYCLEZ0\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__3082\,
            I => \U400_SDRAM.RAM_CYCLEZ0\
        );

    \I__372\ : CascadeMux
    port map (
            O => \N__3077\,
            I => \N__3074\
        );

    \I__371\ : InMux
    port map (
            O => \N__3074\,
            I => \N__3071\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__3071\,
            I => \N__3067\
        );

    \I__369\ : InMux
    port map (
            O => \N__3070\,
            I => \N__3064\
        );

    \I__368\ : Span4Mux_v
    port map (
            O => \N__3067\,
            I => \N__3061\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__3064\,
            I => \N__3058\
        );

    \I__366\ : Odrv4
    port map (
            O => \N__3061\,
            I => \U400_SDRAM.CS1_ENZ0\
        );

    \I__365\ : Odrv4
    port map (
            O => \N__3058\,
            I => \U400_SDRAM.CS1_ENZ0\
        );

    \I__364\ : IoInMux
    port map (
            O => \N__3053\,
            I => \N__3050\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__3050\,
            I => \N__3047\
        );

    \I__362\ : Span4Mux_s3_v
    port map (
            O => \N__3047\,
            I => \N__3044\
        );

    \I__361\ : Span4Mux_v
    port map (
            O => \N__3044\,
            I => \N__3041\
        );

    \I__360\ : Odrv4
    port map (
            O => \N__3041\,
            I => \CS1n_c\
        );

    \I__359\ : IoInMux
    port map (
            O => \N__3038\,
            I => \N__3035\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__3035\,
            I => \N__3032\
        );

    \I__357\ : Odrv4
    port map (
            O => \N__3032\,
            I => \CASn_c\
        );

    \I__356\ : IoInMux
    port map (
            O => \N__3029\,
            I => \N__3026\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__3026\,
            I => \N__3023\
        );

    \I__354\ : Odrv12
    port map (
            O => \N__3023\,
            I => \WEn_c\
        );

    \I__353\ : InMux
    port map (
            O => \N__3020\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_7\
        );

    \I__352\ : SRMux
    port map (
            O => \N__3017\,
            I => \N__3014\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__3014\,
            I => \N__3010\
        );

    \I__350\ : SRMux
    port map (
            O => \N__3013\,
            I => \N__3007\
        );

    \I__349\ : Span4Mux_h
    port map (
            O => \N__3010\,
            I => \N__3004\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__3007\,
            I => \N__3001\
        );

    \I__347\ : Span4Mux_s0_h
    port map (
            O => \N__3004\,
            I => \N__2996\
        );

    \I__346\ : Span4Mux_h
    port map (
            O => \N__3001\,
            I => \N__2996\
        );

    \I__345\ : Odrv4
    port map (
            O => \N__2996\,
            I => \U400_SDRAM.SDRAM_COUNTER_RNIV59H2Z0Z_1\
        );

    \I__344\ : InMux
    port map (
            O => \N__2993\,
            I => \N__2989\
        );

    \I__343\ : InMux
    port map (
            O => \N__2992\,
            I => \N__2986\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2989\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__2986\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__340\ : InMux
    port map (
            O => \N__2981\,
            I => \N__2977\
        );

    \I__339\ : InMux
    port map (
            O => \N__2980\,
            I => \N__2974\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__2977\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2974\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__336\ : InMux
    port map (
            O => \N__2969\,
            I => \N__2965\
        );

    \I__335\ : InMux
    port map (
            O => \N__2968\,
            I => \N__2962\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__2965\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2962\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__332\ : InMux
    port map (
            O => \N__2957\,
            I => \N__2953\
        );

    \I__331\ : InMux
    port map (
            O => \N__2956\,
            I => \N__2950\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__2953\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2950\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__328\ : InMux
    port map (
            O => \N__2945\,
            I => \N__2941\
        );

    \I__327\ : InMux
    port map (
            O => \N__2944\,
            I => \N__2938\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__2941\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_8\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__2938\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_8\
        );

    \I__324\ : CascadeMux
    port map (
            O => \N__2933\,
            I => \U400_SDRAM.un1_REFRESH_COUNTERlt7_0_cascade_\
        );

    \I__323\ : InMux
    port map (
            O => \N__2930\,
            I => \N__2926\
        );

    \I__322\ : InMux
    port map (
            O => \N__2929\,
            I => \N__2923\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__2926\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2923\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__319\ : CascadeMux
    port map (
            O => \N__2918\,
            I => \U400_SDRAM.N_337_1_cascade_\
        );

    \I__318\ : CascadeMux
    port map (
            O => \N__2915\,
            I => \U400_SDRAM.N_64_cascade_\
        );

    \I__317\ : InMux
    port map (
            O => \N__2912\,
            I => \N__2909\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__2909\,
            I => \U400_SDRAM.CS1_EN_0\
        );

    \I__315\ : InMux
    port map (
            O => \N__2906\,
            I => \N__2901\
        );

    \I__314\ : InMux
    port map (
            O => \N__2905\,
            I => \N__2898\
        );

    \I__313\ : InMux
    port map (
            O => \N__2904\,
            I => \N__2895\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__2901\,
            I => \N__2892\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2898\,
            I => \U400_SDRAM.N_64\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__2895\,
            I => \U400_SDRAM.N_64\
        );

    \I__309\ : Odrv4
    port map (
            O => \N__2892\,
            I => \U400_SDRAM.N_64\
        );

    \I__308\ : IoInMux
    port map (
            O => \N__2885\,
            I => \N__2882\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2882\,
            I => \RESETn_c_i\
        );

    \I__306\ : InMux
    port map (
            O => \N__2879\,
            I => \N__2875\
        );

    \I__305\ : InMux
    port map (
            O => \N__2878\,
            I => \N__2872\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__2875\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__2872\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__302\ : CascadeMux
    port map (
            O => \N__2867\,
            I => \N__2862\
        );

    \I__301\ : InMux
    port map (
            O => \N__2866\,
            I => \N__2857\
        );

    \I__300\ : InMux
    port map (
            O => \N__2865\,
            I => \N__2857\
        );

    \I__299\ : InMux
    port map (
            O => \N__2862\,
            I => \N__2854\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__2857\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__2854\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__296\ : InMux
    port map (
            O => \N__2849\,
            I => \N__2846\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2846\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__294\ : InMux
    port map (
            O => \N__2843\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_1\
        );

    \I__293\ : InMux
    port map (
            O => \N__2840\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_2\
        );

    \I__292\ : InMux
    port map (
            O => \N__2837\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_3\
        );

    \I__291\ : InMux
    port map (
            O => \N__2834\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_4\
        );

    \I__290\ : InMux
    port map (
            O => \N__2831\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_5\
        );

    \I__289\ : InMux
    port map (
            O => \N__2828\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_6\
        );

    \I__288\ : CascadeMux
    port map (
            O => \N__2825\,
            I => \N__2822\
        );

    \I__287\ : InMux
    port map (
            O => \N__2822\,
            I => \N__2819\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__2819\,
            I => \A_c_21\
        );

    \I__285\ : IoInMux
    port map (
            O => \N__2816\,
            I => \N__2813\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__2813\,
            I => \N__2810\
        );

    \I__283\ : IoSpan4Mux
    port map (
            O => \N__2810\,
            I => \N__2807\
        );

    \I__282\ : Span4Mux_s0_h
    port map (
            O => \N__2807\,
            I => \N__2804\
        );

    \I__281\ : Span4Mux_v
    port map (
            O => \N__2804\,
            I => \N__2800\
        );

    \I__280\ : InMux
    port map (
            O => \N__2803\,
            I => \N__2797\
        );

    \I__279\ : Odrv4
    port map (
            O => \N__2800\,
            I => \BANK0_c\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2797\,
            I => \BANK0_c\
        );

    \I__277\ : IoInMux
    port map (
            O => \N__2792\,
            I => \N__2789\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__2789\,
            I => \N__2786\
        );

    \I__275\ : Span4Mux_s0_h
    port map (
            O => \N__2786\,
            I => \N__2783\
        );

    \I__274\ : Span4Mux_v
    port map (
            O => \N__2783\,
            I => \N__2779\
        );

    \I__273\ : InMux
    port map (
            O => \N__2782\,
            I => \N__2776\
        );

    \I__272\ : Span4Mux_v
    port map (
            O => \N__2779\,
            I => \N__2771\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__2776\,
            I => \N__2771\
        );

    \I__270\ : Odrv4
    port map (
            O => \N__2771\,
            I => \CONSTANT_ONE_NET\
        );

    \I__269\ : CascadeMux
    port map (
            O => \N__2768\,
            I => \N__2765\
        );

    \I__268\ : InMux
    port map (
            O => \N__2765\,
            I => \N__2762\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__2762\,
            I => \N__2759\
        );

    \I__266\ : Span12Mux_s2_h
    port map (
            O => \N__2759\,
            I => \N__2756\
        );

    \I__265\ : Odrv12
    port map (
            O => \N__2756\,
            I => \A_c_22\
        );

    \I__264\ : IoInMux
    port map (
            O => \N__2753\,
            I => \N__2750\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__2750\,
            I => \N__2747\
        );

    \I__262\ : IoSpan4Mux
    port map (
            O => \N__2747\,
            I => \N__2744\
        );

    \I__261\ : IoSpan4Mux
    port map (
            O => \N__2744\,
            I => \N__2740\
        );

    \I__260\ : InMux
    port map (
            O => \N__2743\,
            I => \N__2737\
        );

    \I__259\ : Odrv4
    port map (
            O => \N__2740\,
            I => \BANK1_c\
        );

    \I__258\ : LocalMux
    port map (
            O => \N__2737\,
            I => \BANK1_c\
        );

    \I__257\ : InMux
    port map (
            O => \N__2732\,
            I => \N__2726\
        );

    \I__256\ : InMux
    port map (
            O => \N__2731\,
            I => \N__2726\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__2726\,
            I => \U400_SDRAM.un1_SDRAM_COUNTER59_0\
        );

    \I__254\ : InMux
    port map (
            O => \N__2723\,
            I => \N__2720\
        );

    \I__253\ : LocalMux
    port map (
            O => \N__2720\,
            I => \U400_SDRAM.SDRAM_CMD_5_sqmuxa\
        );

    \I__252\ : IoInMux
    port map (
            O => \N__2717\,
            I => \N__2714\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__2714\,
            I => \N__2711\
        );

    \I__250\ : IoSpan4Mux
    port map (
            O => \N__2711\,
            I => \N__2708\
        );

    \I__249\ : IoSpan4Mux
    port map (
            O => \N__2708\,
            I => \N__2705\
        );

    \I__248\ : Span4Mux_s2_h
    port map (
            O => \N__2705\,
            I => \N__2702\
        );

    \I__247\ : Sp12to4
    port map (
            O => \N__2702\,
            I => \N__2699\
        );

    \I__246\ : Odrv12
    port map (
            O => \N__2699\,
            I => \CLK40_ibuf_gb_io_gb_input\
        );

    \INVU400_SDRAM.MA_nesr_1C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_1C_net\,
            I => \N__5498\
        );

    \INVU400_SDRAM.MA_nesr_10C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_10C_net\,
            I => \N__5497\
        );

    \INVU400_SDRAM.BURSTC\ : INV
    port map (
            O => \INVU400_SDRAM.BURSTC_net\,
            I => \N__5493\
        );

    \INVU400_SDRAM.MA_nesr_11C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_11C_net\,
            I => \N__5496\
        );

    \INVU400_SDRAM.SDRAM_COUNTER_2C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            I => \N__5490\
        );

    \INVU400_SDRAM.MA_nesr_3C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_3C_net\,
            I => \N__5489\
        );

    \INVU400_SDRAM.SDRAM_CMD_0C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_CMD_0C_net\,
            I => \N__5483\
        );

    \INVU400_SDRAM.SDRAM_COUNTER_0C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_COUNTER_0C_net\,
            I => \N__5487\
        );

    \INVU400_SDRAM.TACKC\ : INV
    port map (
            O => \INVU400_SDRAM.TACKC_net\,
            I => \N__5491\
        );

    \INVU400_SDRAM.MA_nesr_6C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_6C_net\,
            I => \N__5485\
        );

    \INVU400_SDRAM.SDRAM_CMD_1C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_CMD_1C_net\,
            I => \N__5480\
        );

    \INVU400_SDRAM.SDRAM_CONFIGUREDC\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_CONFIGUREDC_net\,
            I => \N__5486\
        );

    \INVU400_SDRAM.SDRAM_COUNTER_1C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_COUNTER_1C_net\,
            I => \N__5488\
        );

    \INVU400_SDRAM.RASnC\ : INV
    port map (
            O => \INVU400_SDRAM.RASnC_net\,
            I => \N__5476\
        );

    \INVU400_SDRAM.CS1nC\ : INV
    port map (
            O => \INVU400_SDRAM.CS1nC_net\,
            I => \N__5474\
        );

    \INVU400_SDRAM.CS0_ENC\ : INV
    port map (
            O => \INVU400_SDRAM.CS0_ENC_net\,
            I => \N__5482\
        );

    \INVU400_SDRAM.REFRESH_COUNTER_2C\ : INV
    port map (
            O => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            I => \N__5484\
        );

    \INVU400_SDRAM.RAM_CYCLEC\ : INV
    port map (
            O => \INVU400_SDRAM.RAM_CYCLEC_net\,
            I => \N__5475\
        );

    \INVU400_SDRAM.CS1_ENC\ : INV
    port map (
            O => \INVU400_SDRAM.CS1_ENC_net\,
            I => \N__5477\
        );

    \INVU400_SDRAM.BANK0C\ : INV
    port map (
            O => \INVU400_SDRAM.BANK0C_net\,
            I => \N__5479\
        );

    \INVU400_SDRAM.REFRESH_COUNTER_1C\ : INV
    port map (
            O => \INVU400_SDRAM.REFRESH_COUNTER_1C_net\,
            I => \N__5481\
        );

    \IN_MUX_bfv_2_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_4_0_\
        );

    \IN_MUX_bfv_6_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_6_0_\
        );

    \CLK40_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2717\,
            GLOBALBUFFEROUTPUT => \CLK40_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2885\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_1_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__2866\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2879\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__3013\
        );

    \U400_SDRAM.REFRESH_COUNTER_0_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2865\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__3013\
        );

    \U400_SDRAM.BANK0_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__2803\,
            in1 => \N__5082\,
            in2 => \N__2825\,
            in3 => \N__2731\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.BANK0C_net\,
            ce => 'H',
            sr => \N__6348\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__2782\,
            in1 => \N__5081\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.BANK1_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__2732\,
            in1 => \N__2743\,
            in2 => \N__2768\,
            in3 => \N__5083\,
            lcout => \BANK1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.BANK0C_net\,
            ce => 'H',
            sr => \N__6348\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIV59H2_1_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__5337\,
            in1 => \N__3530\,
            in2 => \_gnd_net_\,
            in3 => \N__4655\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_RNIV59H2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.CS1_EN_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__3108\,
            in1 => \N__2905\,
            in2 => \_gnd_net_\,
            in3 => \N__2912\,
            lcout => \U400_SDRAM.CS1_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS1_ENC_net\,
            ce => 'H',
            sr => \N__6345\
        );

    \U400_SDRAM.RAM_CYCLE_RNO_0_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__4406\,
            in1 => \N__3324\,
            in2 => \N__3110\,
            in3 => \N__3625\,
            lcout => \U400_SDRAM.SDRAM_CMD_5_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.WRITE_CYCLE_RNIF1VQ5_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3521\,
            in2 => \_gnd_net_\,
            in3 => \N__5405\,
            lcout => \U400_SDRAM.un1_SDRAM_COUNTER59_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__4826\,
            in1 => \N__5406\,
            in2 => \N__3092\,
            in3 => \N__2723\,
            lcout => \U400_SDRAM.RAM_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.RAM_CYCLEC_net\,
            ce => 'H',
            sr => \N__6344\
        );

    \RESETn_ibuf_RNIM9SF_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5347\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.un3_REFRESH_COUNTER_cry_1_c_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2878\,
            in2 => \N__2867\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_4_0_\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_2_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2849\,
            in2 => \_gnd_net_\,
            in3 => \N__2843\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un3_REFRESH_COUNTER_cry_1\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_2\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3017\
        );

    \U400_SDRAM.REFRESH_COUNTER_3_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2993\,
            in2 => \_gnd_net_\,
            in3 => \N__2840\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un3_REFRESH_COUNTER_cry_2\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_3\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3017\
        );

    \U400_SDRAM.REFRESH_COUNTER_4_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2969\,
            in2 => \_gnd_net_\,
            in3 => \N__2837\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un3_REFRESH_COUNTER_cry_3\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_4\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3017\
        );

    \U400_SDRAM.REFRESH_COUNTER_5_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2981\,
            in2 => \_gnd_net_\,
            in3 => \N__2834\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un3_REFRESH_COUNTER_cry_4\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_5\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3017\
        );

    \U400_SDRAM.REFRESH_COUNTER_6_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2957\,
            in2 => \_gnd_net_\,
            in3 => \N__2831\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un3_REFRESH_COUNTER_cry_5\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_6\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3017\
        );

    \U400_SDRAM.REFRESH_COUNTER_7_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2930\,
            in2 => \_gnd_net_\,
            in3 => \N__2828\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un3_REFRESH_COUNTER_cry_6\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_7\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3017\
        );

    \U400_SDRAM.REFRESH_COUNTER_8_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2945\,
            in2 => \_gnd_net_\,
            in3 => \N__3020\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3017\
        );

    \U400_SDRAM.CS0_EN_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__3109\,
            in1 => \N__2904\,
            in2 => \_gnd_net_\,
            in3 => \N__3116\,
            lcout => \U400_SDRAM.CS0_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS0_ENC_net\,
            ce => 'H',
            sr => \N__6350\
        );

    \U400_SDRAM.REFRESH_COUNTER_RNILA301_3_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__2992\,
            in1 => \N__2980\,
            in2 => \_gnd_net_\,
            in3 => \N__2968\,
            lcout => OPEN,
            ltout => \U400_SDRAM.un1_REFRESH_COUNTERlt7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_RNIJU602_8_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__2956\,
            in1 => \N__2944\,
            in2 => \N__2933\,
            in3 => \N__2929\,
            lcout => \U400_SDRAM.N_337_1\,
            ltout => \U400_SDRAM.N_337_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNIS9I32_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2918\,
            in3 => \N__4388\,
            lcout => \U400_SDRAM.N_64\,
            ltout => \U400_SDRAM.N_64_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI6JJA4_1_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__5346\,
            in1 => \N__3789\,
            in2 => \N__2915\,
            in3 => \N__4654\,
            lcout => \U400_SDRAM.N_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.CS1_EN_RNO_0_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__3070\,
            in1 => \N__3734\,
            in2 => \N__3140\,
            in3 => \N__3146\,
            lcout => \U400_SDRAM.CS1_EN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_RNIP6F34_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4405\,
            in1 => \N__3752\,
            in2 => \N__3325\,
            in3 => \N__3611\,
            lcout => \U400_SDRAM.SDRAM_CMD_1_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__3612\,
            in1 => \N__3347\,
            in2 => \_gnd_net_\,
            in3 => \N__2906\,
            lcout => \U400_SDRAM.N_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_RNI8DRF2_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__3317\,
            in1 => \N__4645\,
            in2 => \_gnd_net_\,
            in3 => \N__3610\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_72_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNI9NVF9_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__3356\,
            in1 => \N__3791\,
            in2 => \N__3149\,
            in3 => \N__4404\,
            lcout => \U400_SDRAM.N_40\,
            ltout => \U400_SDRAM.N_40_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.CS0_EN_RNO_0_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__3733\,
            in1 => \N__3136\,
            in2 => \N__3119\,
            in3 => \N__3283\,
            lcout => \U400_SDRAM.CS0_EN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIA9172_1_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__4646\,
            in1 => \N__5348\,
            in2 => \_gnd_net_\,
            in3 => \N__3790\,
            lcout => \U400_SDRAM.N_115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_RNIFGBJ4_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__3655\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3613\,
            lcout => \U400_SDRAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__3209\,
            in1 => \N__3088\,
            in2 => \_gnd_net_\,
            in3 => \N__3631\,
            lcout => \U400_SDRAM.RAM_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5478\,
            ce => 'H',
            sr => \N__6346\
        );

    \U400_SDRAM.CS1n_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__6593\,
            in1 => \N__5872\,
            in2 => \N__3077\,
            in3 => \N__5753\,
            lcout => \CS1n_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS1nC_net\,
            ce => 'H',
            sr => \N__6347\
        );

    \U400_SDRAM.CASn_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5873\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS1nC_net\,
            ce => 'H',
            sr => \N__6347\
        );

    \U400_SDRAM.WEn_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5751\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS1nC_net\,
            ce => 'H',
            sr => \N__6347\
        );

    \U400_SDRAM.RASn_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6595\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.RASnC_net\,
            ce => 'H',
            sr => \N__6349\
        );

    \U400_SDRAM.CS0n_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__6594\,
            in1 => \N__5874\,
            in2 => \N__3290\,
            in3 => \N__5752\,
            lcout => \CS0n_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.RASnC_net\,
            ce => 'H',
            sr => \N__6349\
        );

    \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_2_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3263\,
            in2 => \_gnd_net_\,
            in3 => \N__3251\,
            lcout => \U400_ADDRESS_DECODE_RAM_SPACE_i_o3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_1_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__3239\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3227\,
            lcout => \U400_ADDRESS_DECODE_RAM_SPACE_i_o3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__3197\,
            in1 => \N__3181\,
            in2 => \N__3164\,
            in3 => \N__3221\,
            lcout => \U400_SDRAM.N_101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.RAM_SPACE_i_o3dup_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__3196\,
            in1 => \N__5336\,
            in2 => \N__3182\,
            in3 => \N__3160\,
            lcout => \RAM_SPACE_i_o3dup\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_1_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__3584\,
            in1 => \N__4204\,
            in2 => \N__4034\,
            in3 => \N__3667\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_1C_net\,
            ce => \N__4151\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4378\,
            in2 => \_gnd_net_\,
            in3 => \N__3689\,
            lcout => \U400_SDRAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_CONFIGUREDC_net\,
            ce => 'H',
            sr => \N__6351\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIQQB91_0_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__4741\,
            in1 => \N__5049\,
            in2 => \_gnd_net_\,
            in3 => \N__4889\,
            lcout => \U400_SDRAM.N_113\,
            ltout => \U400_SDRAM.N_113_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.WRITE_CYCLE_RNIMQFN1_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__4968\,
            in1 => \N__4600\,
            in2 => \N__3362\,
            in3 => \N__4347\,
            lcout => \U400_SDRAM.N_39\,
            ltout => \U400_SDRAM.N_39_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNIGGGC5_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__4348\,
            in1 => \N__3745\,
            in2 => \N__3359\,
            in3 => \N__3687\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_1_sqmuxa_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6190\,
            in1 => \N__3780\,
            in2 => \N__6119\,
            in3 => \N__4601\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_a2_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNINU7A_3_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__4346\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4471\,
            lcout => \U400_SDRAM.N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI6C8G1_1_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3557\,
            in2 => \_gnd_net_\,
            in3 => \N__4602\,
            lcout => \U400_SDRAM.N_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_5_2_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4475\,
            in2 => \_gnd_net_\,
            in3 => \N__4603\,
            lcout => \U400_SDRAM.N_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__3332\,
            in1 => \N__4604\,
            in2 => \_gnd_net_\,
            in3 => \N__5066\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_78_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5309\,
            in1 => \N__4751\,
            in2 => \N__3335\,
            in3 => \N__4384\,
            lcout => \U400_SDRAM.N_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_RNI2IKT2_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3331\,
            in1 => \N__5067\,
            in2 => \N__4813\,
            in3 => \N__3626\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI4LJ09_1_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__4605\,
            in1 => \N__3878\,
            in2 => \N__3503\,
            in3 => \N__4916\,
            lcout => \U400_SDRAM.N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6114\,
            in1 => \N__6170\,
            in2 => \_gnd_net_\,
            in3 => \N__3627\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_3_sqmuxa_0_a3_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_4_1_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__4120\,
            in1 => \N__4508\,
            in2 => \_gnd_net_\,
            in3 => \N__4641\,
            lcout => \U400_SDRAM.SDRAM_CMD_cnst_0_0_103_i_i_a3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_3_1_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__4642\,
            in1 => \N__3563\,
            in2 => \N__5308\,
            in3 => \N__3823\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_91_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__4919\,
            in1 => \N__5273\,
            in2 => \N__3500\,
            in3 => \N__3497\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_0_0_103_i_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_1_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__3491\,
            in1 => \N__5831\,
            in2 => \N__3485\,
            in3 => \N__4014\,
            lcout => \U400_SDRAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_CMD_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_6_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__3482\,
            in1 => \N__6591\,
            in2 => \N__3467\,
            in3 => \N__6461\,
            lcout => \MA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_6C_net\,
            ce => \N__6421\,
            sr => \N__6352\
        );

    \U400_SDRAM.MA_nesr_4_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__3440\,
            in1 => \N__6590\,
            in2 => \N__3431\,
            in3 => \N__6460\,
            lcout => \MA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_6C_net\,
            ce => \N__6421\,
            sr => \N__6352\
        );

    \U400_SDRAM.MA_nesr_7_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__6462\,
            in1 => \N__3404\,
            in2 => \N__3386\,
            in3 => \N__6592\,
            lcout => \MA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_6C_net\,
            ce => \N__6421\,
            sr => \N__6352\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__6118\,
            in1 => \N__6191\,
            in2 => \_gnd_net_\,
            in3 => \N__3635\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_4_sqmuxa_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111010"
        )
    port map (
            in0 => \N__3539\,
            in1 => \N__5174\,
            in2 => \N__4106\,
            in3 => \N__4070\,
            lcout => \U400_SDRAM.TACKZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.TACKC_net\,
            ce => 'H',
            sr => \N__6353\
        );

    \U400_SDRAM.WRITE_CYCLE_RNIJKOA_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4956\,
            in2 => \_gnd_net_\,
            in3 => \N__4577\,
            lcout => \U400_SDRAM.N_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.WRITE_CYCLE_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__4957\,
            in1 => \N__3578\,
            in2 => \_gnd_net_\,
            in3 => \N__5417\,
            lcout => \U400_SDRAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.TACKC_net\,
            ce => 'H',
            sr => \N__6353\
        );

    \U400_SDRAM.RAM_CYCLE_RNO_2_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__4468\,
            in1 => \N__3558\,
            in2 => \N__4777\,
            in3 => \N__4345\,
            lcout => \U400_SDRAM.N_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_1_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__3559\,
            in1 => \N__4773\,
            in2 => \_gnd_net_\,
            in3 => \N__4469\,
            lcout => \U400_SDRAM.N_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNILS7A_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4552\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4344\,
            lcout => \U400_SDRAM.N_20\,
            ltout => \U400_SDRAM.N_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNITAGQ1_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3533\,
            in3 => \N__3776\,
            lcout => \U400_SDRAM.N_35\,
            ltout => \U400_SDRAM.N_35_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.WRITE_CYCLE_RNI6QCS5_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__5339\,
            in1 => \N__3517\,
            in2 => \N__3506\,
            in3 => \N__3688\,
            lcout => \U400_SDRAM.N_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4227\,
            in1 => \N__4248\,
            in2 => \N__4166\,
            in3 => \N__4264\,
            lcout => \U400_SDRAM.N_44\,
            ltout => \U400_SDRAM.N_44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_0_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4467\,
            in1 => \N__4724\,
            in2 => \N__3794\,
            in3 => \N__5048\,
            lcout => \U400_SDRAM.N_108\,
            ltout => \U400_SDRAM.N_108_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_1_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3755\,
            in3 => \N__4553\,
            lcout => \U400_SDRAM.N_109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111001111"
        )
    port map (
            in0 => \N__3732\,
            in1 => \N__4064\,
            in2 => \N__5335\,
            in3 => \N__4377\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_0_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__3716\,
            in1 => \N__3701\,
            in2 => \N__3692\,
            in3 => \N__4199\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_0C_net\,
            ce => \N__4149\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNITAGQ1_3_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__4725\,
            in1 => \N__3856\,
            in2 => \N__4496\,
            in3 => \N__4050\,
            lcout => \U400_SDRAM.SDRAM_CMD_3_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_3_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__4198\,
            in1 => \N__3671\,
            in2 => \N__4277\,
            in3 => \N__3644\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_0C_net\,
            ce => \N__4149\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIR5PD_3_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4470\,
            in2 => \_gnd_net_\,
            in3 => \N__4742\,
            lcout => \U400_SDRAM.N_46\,
            ltout => \U400_SDRAM.N_46_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNII7IR_0_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__4599\,
            in1 => \_gnd_net_\,
            in2 => \N__3638\,
            in3 => \N__5053\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI189H2_0_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001111111111"
        )
    port map (
            in0 => \N__4915\,
            in1 => \N__5296\,
            in2 => \N__3884\,
            in3 => \N__3816\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNIKPF05_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__4386\,
            in1 => \N__4051\,
            in2 => \N__3881\,
            in3 => \N__4988\,
            lcout => \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIO2PD_0_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4743\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5054\,
            lcout => \U400_SDRAM.N_336_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_4_2_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__4969\,
            in1 => \N__4744\,
            in2 => \N__3872\,
            in3 => \N__4385\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_97_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_3_2_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4812\,
            in2 => \N__3863\,
            in3 => \N__3860\,
            lcout => \U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_1_0_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101111"
        )
    port map (
            in0 => \N__4757\,
            in1 => \_gnd_net_\,
            in2 => \N__5322\,
            in3 => \N__4918\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_0_1_66_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_0_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011100100"
        )
    port map (
            in0 => \N__4016\,
            in1 => \N__5722\,
            in2 => \N__3845\,
            in3 => \N__4994\,
            lcout => \U400_SDRAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_CMD_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_RNO_0_5_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100101110"
        )
    port map (
            in0 => \N__5843\,
            in1 => \N__6529\,
            in2 => \N__3842\,
            in3 => \N__5713\,
            lcout => \U400_SDRAM.MA_5_iv_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111010000"
        )
    port map (
            in0 => \N__4750\,
            in1 => \N__3824\,
            in2 => \N__5084\,
            in3 => \N__3800\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_2_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010101010"
        )
    port map (
            in0 => \N__6538\,
            in1 => \N__3998\,
            in2 => \N__4019\,
            in3 => \N__4015\,
            lcout => \U400_SDRAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_CMD_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__4749\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5077\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_a2_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110101"
        )
    port map (
            in0 => \N__5292\,
            in1 => \N__4387\,
            in2 => \N__4001\,
            in3 => \N__4917\,
            lcout => \U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_3_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__6456\,
            in1 => \N__3992\,
            in2 => \N__6578\,
            in3 => \N__3983\,
            lcout => \MA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_3C_net\,
            ce => \N__6418\,
            sr => \N__6355\
        );

    \U400_SDRAM.MA_nesr_12_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6549\,
            in1 => \N__5866\,
            in2 => \N__3953\,
            in3 => \N__5725\,
            lcout => \MA_c_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_3C_net\,
            ce => \N__6418\,
            sr => \N__6355\
        );

    \U400_SDRAM.MA_nesr_5_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__3920\,
            in1 => \N__3905\,
            in2 => \_gnd_net_\,
            in3 => \N__6455\,
            lcout => \MA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_3C_net\,
            ce => \N__6418\,
            sr => \N__6355\
        );

    \U400_SDRAM.SDRAM_CMD_RNIMFKP_0_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011011110111"
        )
    port map (
            in0 => \N__6577\,
            in1 => \N__5861\,
            in2 => \N__6371\,
            in3 => \N__5723\,
            lcout => \U400_SDRAM.un1_MA21_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6576\,
            in1 => \N__5862\,
            in2 => \_gnd_net_\,
            in3 => \N__5724\,
            lcout => \U400_SDRAM.MA20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_6_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110110011"
        )
    port map (
            in0 => \N__4738\,
            in1 => \N__4400\,
            in2 => \N__4502\,
            in3 => \N__4900\,
            lcout => \U400_SDRAM.un1_SDRAM_COUNTER59_4_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI5LLK_0_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000100010"
        )
    port map (
            in0 => \N__4476\,
            in1 => \N__4643\,
            in2 => \_gnd_net_\,
            in3 => \N__5050\,
            lcout => \U400_SDRAM.N_8\,
            ltout => \U400_SDRAM.N_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_4_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__4249\,
            in1 => \N__4978\,
            in2 => \N__4091\,
            in3 => \N__4228\,
            lcout => \U400_SDRAM.N_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_RNIPSFM_0_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5204\,
            in2 => \_gnd_net_\,
            in3 => \N__5165\,
            lcout => \U400_SDRAM.N_244_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_3_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001011110000"
        )
    port map (
            in0 => \N__5052\,
            in1 => \N__4737\,
            in2 => \N__4817\,
            in3 => \N__4649\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_0_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__4058\,
            in1 => \N__4088\,
            in2 => \N__4082\,
            in3 => \N__4079\,
            lcout => \U400_SDRAM.N_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__4739\,
            in1 => \N__4650\,
            in2 => \N__4503\,
            in3 => \N__4052\,
            lcout => \U400_SDRAM.N_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_5_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4477\,
            in1 => \N__4644\,
            in2 => \N__4982\,
            in3 => \N__5051\,
            lcout => \U400_SDRAM.N_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNID8F21_0_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5047\,
            in2 => \_gnd_net_\,
            in3 => \N__4888\,
            lcout => \U400_SDRAM.N_48\,
            ltout => OPEN,
            carryin => \bfn_6_6_0_\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_1_1_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4651\,
            in2 => \_gnd_net_\,
            in3 => \N__4283\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_s_1\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_0\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_2_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4200\,
            in1 => \N__4740\,
            in2 => \_gnd_net_\,
            in3 => \N__4280\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_1\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_2\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__4150\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_1_3_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4501\,
            in2 => \_gnd_net_\,
            in3 => \N__4268\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_s_3\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_2\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_4_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4201\,
            in1 => \N__4265\,
            in2 => \_gnd_net_\,
            in3 => \N__4253\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_3\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_4\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__4150\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_5_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4208\,
            in1 => \N__4250\,
            in2 => \_gnd_net_\,
            in3 => \N__4232\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_4\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_5\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__4150\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_6_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4202\,
            in1 => \N__4229\,
            in2 => \_gnd_net_\,
            in3 => \N__4211\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_5\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_6\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__4150\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_7_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__4165\,
            in1 => \N__4203\,
            in2 => \_gnd_net_\,
            in3 => \N__4169\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__4150\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_7_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4971\,
            in1 => \N__4728\,
            in2 => \N__4856\,
            in3 => \N__4913\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_56_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_2_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__4121\,
            in1 => \N__4972\,
            in2 => \N__4109\,
            in3 => \N__4653\,
            lcout => \U400_SDRAM.TACK_7_iv_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_0_0_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__4925\,
            in1 => \N__4652\,
            in2 => \_gnd_net_\,
            in3 => \N__5068\,
            lcout => \U400_SDRAM.N_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNITTB91_3_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__4478\,
            in1 => \N__4726\,
            in2 => \_gnd_net_\,
            in3 => \N__4912\,
            lcout => \U400_SDRAM.N_110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.WRITE_CYCLE_RNIT04E_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__4970\,
            in1 => \N__4727\,
            in2 => \_gnd_net_\,
            in3 => \N__4403\,
            lcout => \U400_SDRAM.N_13\,
            ltout => \U400_SDRAM.N_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_RNO_1_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__4914\,
            in1 => \N__4855\,
            in2 => \N__4841\,
            in3 => \N__4838\,
            lcout => \U400_SDRAM.un1_SDRAM_COUNTER59_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_4_0_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__4402\,
            in1 => \N__4805\,
            in2 => \_gnd_net_\,
            in3 => \N__4648\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_33_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_2_0_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__4500\,
            in1 => \N__4289\,
            in2 => \N__4784\,
            in3 => \N__4781\,
            lcout => \U400_SDRAM.SDRAM_CMD_cnst_0_1_66_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_3_0_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011010"
        )
    port map (
            in0 => \N__4748\,
            in1 => \N__4647\,
            in2 => \N__4507\,
            in3 => \N__4401\,
            lcout => \U400_SDRAM.N_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_0_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010000011111111"
        )
    port map (
            in0 => \N__5360\,
            in1 => \N__5179\,
            in2 => \N__5138\,
            in3 => \N__5354\,
            lcout => \U400_SDRAM.TA_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5494\,
            ce => 'H',
            sr => \N__6357\
        );

    \U400_SDRAM.TA_EN_i_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011111110101010"
        )
    port map (
            in0 => \N__6223\,
            in1 => \N__5122\,
            in2 => \N__5338\,
            in3 => \N__5144\,
            lcout => \TA_EN_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5494\,
            ce => 'H',
            sr => \N__6357\
        );

    \U400_SDRAM.TA_COUNTER_2_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5668\,
            lcout => \U400_SDRAM.TA_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5494\,
            ce => 'H',
            sr => \N__6357\
        );

    \U400_SDRAM.TA_COUNTER_1_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5203\,
            in2 => \_gnd_net_\,
            in3 => \N__5178\,
            lcout => \U400_SDRAM.TA_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5494\,
            ce => 'H',
            sr => \N__6357\
        );

    \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5524\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5509\,
            lcout => \U400_SDRAM.TA_COUNTER_srsts_0_a4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_RNINB8O_1_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5550\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5667\,
            lcout => \U400_SDRAM.un1_TA_COUNTER_6_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_RNIMKDP_5_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__5531\,
            in1 => \N__5523\,
            in2 => \_gnd_net_\,
            in3 => \N__5381\,
            lcout => \U400_SDRAM.N_243_0\,
            ltout => \U400_SDRAM.N_243_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_EN_i_RNO_0_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__5323\,
            in1 => \N__5202\,
            in2 => \N__5183\,
            in3 => \N__5180\,
            lcout => \U400_SDRAM.N_241_0_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_OUT_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001110110001"
        )
    port map (
            in0 => \N__5137\,
            in1 => \N__5648\,
            in2 => \N__5110\,
            in3 => \N__5123\,
            lcout => \TA_OUT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5492\,
            ce => 'H',
            sr => \N__6354\
        );

    \U400_BYTE_ENABLE.un1_UUBEn_i_0_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__5979\,
            in1 => \N__5919\,
            in2 => \N__6041\,
            in3 => \N__6025\,
            lcout => \N_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_OUT_RNO_0_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__5552\,
            in1 => \N__5669\,
            in2 => \_gnd_net_\,
            in3 => \N__5382\,
            lcout => \U400_SDRAM.TA_OUT_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_11_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6612\,
            in1 => \N__5868\,
            in2 => \N__5642\,
            in3 => \N__5763\,
            lcout => \MA_c_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_11C_net\,
            ce => \N__6422\,
            sr => \N__6362\
        );

    \U400_SDRAM.MA_nesr_9_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6613\,
            in1 => \N__5764\,
            in2 => \N__5878\,
            in3 => \N__5609\,
            lcout => \MA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_11C_net\,
            ce => \N__6422\,
            sr => \N__6362\
        );

    \U400_SDRAM.MA_nesr_8_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__5588\,
            in1 => \N__6614\,
            in2 => \N__5576\,
            in3 => \N__6481\,
            lcout => \MA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_11C_net\,
            ce => \N__6422\,
            sr => \N__6362\
        );

    \U400_SDRAM.TA_COUNTER_4_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5510\,
            lcout => \U400_SDRAM.TA_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5495\,
            ce => 'H',
            sr => \N__6358\
        );

    \U400_SDRAM.TA_COUNTER_5_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5551\,
            lcout => \U400_SDRAM.TA_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5495\,
            ce => 'H',
            sr => \N__6358\
        );

    \U400_SDRAM.TA_COUNTER_3_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5525\,
            in2 => \_gnd_net_\,
            in3 => \N__5383\,
            lcout => \U400_SDRAM.TA_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5495\,
            ce => 'H',
            sr => \N__6358\
        );

    \U400_SDRAM.BURST_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__6172\,
            in1 => \N__5384\,
            in2 => \N__6082\,
            in3 => \N__5416\,
            lcout => \U400_SDRAM.BURSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.BURSTC_net\,
            ce => 'H',
            sr => \N__6356\
        );

    \U400_SDRAM.MA_nesr_10_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001000100"
        )
    port map (
            in0 => \N__6616\,
            in1 => \N__5879\,
            in2 => \N__6299\,
            in3 => \N__5765\,
            lcout => \MA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_10C_net\,
            ce => \N__6419\,
            sr => \N__6363\
        );

    \U400_SDRAM.MA_nesr_0_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__6278\,
            in1 => \N__6615\,
            in2 => \N__6266\,
            in3 => \N__6482\,
            lcout => \MA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_10C_net\,
            ce => \N__6419\,
            sr => \N__6363\
        );

    \U400_BYTE_ENABLE.un1_UMBEn_i_0_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100101000"
        )
    port map (
            in0 => \N__5933\,
            in1 => \N__6186\,
            in2 => \N__6113\,
            in3 => \N__6200\,
            lcout => \N_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_BYTE_ENABLE.un1_LLBEn_i_0_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010100"
        )
    port map (
            in0 => \N__5932\,
            in1 => \N__6185\,
            in2 => \N__6112\,
            in3 => \N__6199\,
            lcout => \N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TAn_obuft_RNO_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6227\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_542_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_BYTE_ENABLE.un1_LLBEn_i_o3_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__6173\,
            in1 => \N__6083\,
            in2 => \N__5978\,
            in3 => \N__6026\,
            lcout => \U400_BYTE_ENABLE.N_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_BYTE_ENABLE.un1_LLBEn_i_x2_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__6171\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6057\,
            lcout => \U400_BYTE_ENABLE.N_54_i\,
            ltout => \U400_BYTE_ENABLE.N_54_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_BYTE_ENABLE.un1_LMBEn_i_0_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011111100"
        )
    port map (
            in0 => \N__6021\,
            in1 => \N__5980\,
            in2 => \N__5936\,
            in3 => \N__5926\,
            lcout => \N_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_RNO_0_1_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101001110"
        )
    port map (
            in0 => \N__6596\,
            in1 => \N__5867\,
            in2 => \N__5780\,
            in3 => \N__5754\,
            lcout => \U400_SDRAM.MA_5_iv_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_1_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__6656\,
            in1 => \N__6644\,
            in2 => \_gnd_net_\,
            in3 => \N__6479\,
            lcout => \MA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_1C_net\,
            ce => \N__6420\,
            sr => \N__6364\
        );

    \U400_SDRAM.MA_nesr_2_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__6632\,
            in1 => \N__6617\,
            in2 => \N__6491\,
            in3 => \N__6480\,
            lcout => \MA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_1C_net\,
            ce => \N__6420\,
            sr => \N__6364\
        );
end \INTERFACE\;

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 22 2025 01:34:21

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U400_TOP" view "INTERFACE"

module U400_TOP (
    SIZ,
    MA,
    A,
    LBENn,
    CS0n,
    UUBEn,
    TAn,
    CLK40,
    RnW,
    BANK1,
    UMBEn,
    WEn,
    LLBEn,
    TSn,
    LMBEn,
    RASn,
    CS1n,
    RESETn,
    CLK_EN,
    CASn,
    BANK0);

    input [1:0] SIZ;
    output [12:0] MA;
    input [31:0] A;
    output LBENn;
    output CS0n;
    output UUBEn;
    output TAn;
    input CLK40;
    input RnW;
    output BANK1;
    output UMBEn;
    output WEn;
    output LLBEn;
    input TSn;
    output LMBEn;
    output RASn;
    output CS1n;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;

    wire N__7004;
    wire N__7003;
    wire N__7002;
    wire N__6995;
    wire N__6994;
    wire N__6993;
    wire N__6986;
    wire N__6985;
    wire N__6984;
    wire N__6977;
    wire N__6976;
    wire N__6975;
    wire N__6968;
    wire N__6967;
    wire N__6966;
    wire N__6959;
    wire N__6958;
    wire N__6957;
    wire N__6950;
    wire N__6949;
    wire N__6948;
    wire N__6941;
    wire N__6940;
    wire N__6939;
    wire N__6932;
    wire N__6931;
    wire N__6930;
    wire N__6923;
    wire N__6922;
    wire N__6921;
    wire N__6914;
    wire N__6913;
    wire N__6912;
    wire N__6905;
    wire N__6904;
    wire N__6903;
    wire N__6896;
    wire N__6895;
    wire N__6894;
    wire N__6887;
    wire N__6886;
    wire N__6885;
    wire N__6878;
    wire N__6877;
    wire N__6876;
    wire N__6869;
    wire N__6868;
    wire N__6867;
    wire N__6860;
    wire N__6859;
    wire N__6858;
    wire N__6851;
    wire N__6850;
    wire N__6849;
    wire N__6842;
    wire N__6841;
    wire N__6840;
    wire N__6833;
    wire N__6832;
    wire N__6831;
    wire N__6824;
    wire N__6823;
    wire N__6822;
    wire N__6815;
    wire N__6814;
    wire N__6813;
    wire N__6806;
    wire N__6805;
    wire N__6804;
    wire N__6797;
    wire N__6796;
    wire N__6795;
    wire N__6788;
    wire N__6787;
    wire N__6786;
    wire N__6779;
    wire N__6778;
    wire N__6777;
    wire N__6770;
    wire N__6769;
    wire N__6768;
    wire N__6761;
    wire N__6760;
    wire N__6759;
    wire N__6752;
    wire N__6751;
    wire N__6750;
    wire N__6743;
    wire N__6742;
    wire N__6741;
    wire N__6734;
    wire N__6733;
    wire N__6732;
    wire N__6725;
    wire N__6724;
    wire N__6723;
    wire N__6716;
    wire N__6715;
    wire N__6714;
    wire N__6707;
    wire N__6706;
    wire N__6705;
    wire N__6698;
    wire N__6697;
    wire N__6696;
    wire N__6689;
    wire N__6688;
    wire N__6687;
    wire N__6680;
    wire N__6679;
    wire N__6678;
    wire N__6671;
    wire N__6670;
    wire N__6669;
    wire N__6662;
    wire N__6661;
    wire N__6660;
    wire N__6653;
    wire N__6652;
    wire N__6651;
    wire N__6644;
    wire N__6643;
    wire N__6642;
    wire N__6635;
    wire N__6634;
    wire N__6633;
    wire N__6626;
    wire N__6625;
    wire N__6624;
    wire N__6617;
    wire N__6616;
    wire N__6615;
    wire N__6608;
    wire N__6607;
    wire N__6606;
    wire N__6599;
    wire N__6598;
    wire N__6597;
    wire N__6590;
    wire N__6589;
    wire N__6588;
    wire N__6581;
    wire N__6580;
    wire N__6579;
    wire N__6572;
    wire N__6571;
    wire N__6570;
    wire N__6563;
    wire N__6562;
    wire N__6561;
    wire N__6554;
    wire N__6553;
    wire N__6552;
    wire N__6545;
    wire N__6544;
    wire N__6543;
    wire N__6536;
    wire N__6535;
    wire N__6534;
    wire N__6527;
    wire N__6526;
    wire N__6525;
    wire N__6518;
    wire N__6517;
    wire N__6516;
    wire N__6509;
    wire N__6508;
    wire N__6507;
    wire N__6500;
    wire N__6499;
    wire N__6498;
    wire N__6491;
    wire N__6490;
    wire N__6489;
    wire N__6482;
    wire N__6481;
    wire N__6480;
    wire N__6473;
    wire N__6472;
    wire N__6471;
    wire N__6464;
    wire N__6463;
    wire N__6462;
    wire N__6455;
    wire N__6454;
    wire N__6453;
    wire N__6446;
    wire N__6445;
    wire N__6444;
    wire N__6437;
    wire N__6436;
    wire N__6435;
    wire N__6428;
    wire N__6427;
    wire N__6426;
    wire N__6409;
    wire N__6406;
    wire N__6403;
    wire N__6400;
    wire N__6397;
    wire N__6394;
    wire N__6391;
    wire N__6388;
    wire N__6385;
    wire N__6384;
    wire N__6383;
    wire N__6380;
    wire N__6377;
    wire N__6376;
    wire N__6375;
    wire N__6372;
    wire N__6367;
    wire N__6364;
    wire N__6361;
    wire N__6360;
    wire N__6359;
    wire N__6356;
    wire N__6351;
    wire N__6348;
    wire N__6343;
    wire N__6338;
    wire N__6335;
    wire N__6332;
    wire N__6325;
    wire N__6322;
    wire N__6319;
    wire N__6318;
    wire N__6315;
    wire N__6314;
    wire N__6311;
    wire N__6308;
    wire N__6305;
    wire N__6304;
    wire N__6303;
    wire N__6302;
    wire N__6301;
    wire N__6300;
    wire N__6299;
    wire N__6298;
    wire N__6297;
    wire N__6292;
    wire N__6289;
    wire N__6286;
    wire N__6283;
    wire N__6278;
    wire N__6275;
    wire N__6272;
    wire N__6267;
    wire N__6264;
    wire N__6257;
    wire N__6256;
    wire N__6255;
    wire N__6250;
    wire N__6247;
    wire N__6244;
    wire N__6241;
    wire N__6238;
    wire N__6235;
    wire N__6232;
    wire N__6229;
    wire N__6226;
    wire N__6217;
    wire N__6208;
    wire N__6205;
    wire N__6204;
    wire N__6203;
    wire N__6200;
    wire N__6199;
    wire N__6198;
    wire N__6195;
    wire N__6192;
    wire N__6191;
    wire N__6190;
    wire N__6189;
    wire N__6188;
    wire N__6185;
    wire N__6182;
    wire N__6179;
    wire N__6176;
    wire N__6173;
    wire N__6168;
    wire N__6163;
    wire N__6162;
    wire N__6161;
    wire N__6156;
    wire N__6153;
    wire N__6150;
    wire N__6143;
    wire N__6140;
    wire N__6137;
    wire N__6134;
    wire N__6129;
    wire N__6124;
    wire N__6115;
    wire N__6114;
    wire N__6113;
    wire N__6110;
    wire N__6109;
    wire N__6108;
    wire N__6105;
    wire N__6104;
    wire N__6103;
    wire N__6100;
    wire N__6097;
    wire N__6094;
    wire N__6091;
    wire N__6090;
    wire N__6089;
    wire N__6088;
    wire N__6087;
    wire N__6082;
    wire N__6079;
    wire N__6078;
    wire N__6073;
    wire N__6070;
    wire N__6065;
    wire N__6060;
    wire N__6057;
    wire N__6056;
    wire N__6055;
    wire N__6050;
    wire N__6049;
    wire N__6048;
    wire N__6047;
    wire N__6046;
    wire N__6043;
    wire N__6042;
    wire N__6037;
    wire N__6030;
    wire N__6029;
    wire N__6026;
    wire N__6023;
    wire N__6020;
    wire N__6017;
    wire N__6012;
    wire N__6009;
    wire N__6006;
    wire N__6003;
    wire N__5998;
    wire N__5995;
    wire N__5990;
    wire N__5987;
    wire N__5984;
    wire N__5975;
    wire N__5972;
    wire N__5965;
    wire N__5960;
    wire N__5953;
    wire N__5950;
    wire N__5947;
    wire N__5944;
    wire N__5941;
    wire N__5938;
    wire N__5937;
    wire N__5936;
    wire N__5935;
    wire N__5934;
    wire N__5933;
    wire N__5932;
    wire N__5929;
    wire N__5928;
    wire N__5927;
    wire N__5926;
    wire N__5925;
    wire N__5924;
    wire N__5923;
    wire N__5922;
    wire N__5921;
    wire N__5920;
    wire N__5887;
    wire N__5884;
    wire N__5881;
    wire N__5878;
    wire N__5875;
    wire N__5872;
    wire N__5869;
    wire N__5866;
    wire N__5863;
    wire N__5860;
    wire N__5857;
    wire N__5856;
    wire N__5853;
    wire N__5850;
    wire N__5849;
    wire N__5842;
    wire N__5841;
    wire N__5838;
    wire N__5835;
    wire N__5832;
    wire N__5829;
    wire N__5824;
    wire N__5821;
    wire N__5818;
    wire N__5817;
    wire N__5816;
    wire N__5813;
    wire N__5812;
    wire N__5805;
    wire N__5802;
    wire N__5797;
    wire N__5794;
    wire N__5791;
    wire N__5788;
    wire N__5785;
    wire N__5782;
    wire N__5779;
    wire N__5776;
    wire N__5773;
    wire N__5770;
    wire N__5767;
    wire N__5764;
    wire N__5761;
    wire N__5758;
    wire N__5755;
    wire N__5752;
    wire N__5751;
    wire N__5748;
    wire N__5745;
    wire N__5744;
    wire N__5743;
    wire N__5742;
    wire N__5741;
    wire N__5738;
    wire N__5735;
    wire N__5728;
    wire N__5725;
    wire N__5724;
    wire N__5721;
    wire N__5718;
    wire N__5715;
    wire N__5712;
    wire N__5709;
    wire N__5706;
    wire N__5697;
    wire N__5694;
    wire N__5691;
    wire N__5686;
    wire N__5685;
    wire N__5682;
    wire N__5681;
    wire N__5680;
    wire N__5679;
    wire N__5676;
    wire N__5675;
    wire N__5672;
    wire N__5665;
    wire N__5664;
    wire N__5661;
    wire N__5658;
    wire N__5655;
    wire N__5652;
    wire N__5649;
    wire N__5646;
    wire N__5643;
    wire N__5640;
    wire N__5635;
    wire N__5632;
    wire N__5629;
    wire N__5624;
    wire N__5617;
    wire N__5614;
    wire N__5613;
    wire N__5610;
    wire N__5607;
    wire N__5604;
    wire N__5601;
    wire N__5596;
    wire N__5595;
    wire N__5590;
    wire N__5587;
    wire N__5584;
    wire N__5581;
    wire N__5578;
    wire N__5575;
    wire N__5572;
    wire N__5571;
    wire N__5566;
    wire N__5563;
    wire N__5560;
    wire N__5557;
    wire N__5556;
    wire N__5555;
    wire N__5554;
    wire N__5553;
    wire N__5552;
    wire N__5551;
    wire N__5548;
    wire N__5545;
    wire N__5542;
    wire N__5541;
    wire N__5538;
    wire N__5535;
    wire N__5528;
    wire N__5527;
    wire N__5526;
    wire N__5525;
    wire N__5524;
    wire N__5523;
    wire N__5522;
    wire N__5519;
    wire N__5516;
    wire N__5513;
    wire N__5510;
    wire N__5507;
    wire N__5504;
    wire N__5499;
    wire N__5494;
    wire N__5491;
    wire N__5490;
    wire N__5489;
    wire N__5488;
    wire N__5485;
    wire N__5482;
    wire N__5479;
    wire N__5474;
    wire N__5471;
    wire N__5464;
    wire N__5461;
    wire N__5456;
    wire N__5453;
    wire N__5450;
    wire N__5443;
    wire N__5440;
    wire N__5437;
    wire N__5432;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5418;
    wire N__5413;
    wire N__5404;
    wire N__5401;
    wire N__5398;
    wire N__5395;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5334;
    wire N__5331;
    wire N__5328;
    wire N__5325;
    wire N__5320;
    wire N__5319;
    wire N__5316;
    wire N__5315;
    wire N__5314;
    wire N__5311;
    wire N__5308;
    wire N__5305;
    wire N__5302;
    wire N__5299;
    wire N__5294;
    wire N__5291;
    wire N__5286;
    wire N__5281;
    wire N__5280;
    wire N__5277;
    wire N__5276;
    wire N__5275;
    wire N__5274;
    wire N__5273;
    wire N__5272;
    wire N__5271;
    wire N__5270;
    wire N__5269;
    wire N__5268;
    wire N__5267;
    wire N__5266;
    wire N__5263;
    wire N__5260;
    wire N__5257;
    wire N__5252;
    wire N__5243;
    wire N__5242;
    wire N__5241;
    wire N__5240;
    wire N__5237;
    wire N__5236;
    wire N__5233;
    wire N__5232;
    wire N__5229;
    wire N__5226;
    wire N__5225;
    wire N__5220;
    wire N__5213;
    wire N__5210;
    wire N__5205;
    wire N__5202;
    wire N__5199;
    wire N__5196;
    wire N__5193;
    wire N__5188;
    wire N__5185;
    wire N__5178;
    wire N__5161;
    wire N__5160;
    wire N__5159;
    wire N__5156;
    wire N__5153;
    wire N__5152;
    wire N__5151;
    wire N__5150;
    wire N__5149;
    wire N__5146;
    wire N__5143;
    wire N__5142;
    wire N__5139;
    wire N__5136;
    wire N__5135;
    wire N__5132;
    wire N__5131;
    wire N__5128;
    wire N__5127;
    wire N__5122;
    wire N__5119;
    wire N__5116;
    wire N__5113;
    wire N__5110;
    wire N__5103;
    wire N__5098;
    wire N__5093;
    wire N__5080;
    wire N__5079;
    wire N__5078;
    wire N__5077;
    wire N__5076;
    wire N__5075;
    wire N__5074;
    wire N__5073;
    wire N__5072;
    wire N__5065;
    wire N__5062;
    wire N__5059;
    wire N__5056;
    wire N__5053;
    wire N__5050;
    wire N__5047;
    wire N__5044;
    wire N__5043;
    wire N__5042;
    wire N__5041;
    wire N__5040;
    wire N__5039;
    wire N__5038;
    wire N__5033;
    wire N__5028;
    wire N__5023;
    wire N__5022;
    wire N__5021;
    wire N__5018;
    wire N__5013;
    wire N__5010;
    wire N__5007;
    wire N__5004;
    wire N__5001;
    wire N__4994;
    wire N__4989;
    wire N__4972;
    wire N__4969;
    wire N__4966;
    wire N__4963;
    wire N__4962;
    wire N__4961;
    wire N__4960;
    wire N__4959;
    wire N__4952;
    wire N__4951;
    wire N__4950;
    wire N__4949;
    wire N__4948;
    wire N__4947;
    wire N__4946;
    wire N__4941;
    wire N__4940;
    wire N__4939;
    wire N__4938;
    wire N__4935;
    wire N__4930;
    wire N__4929;
    wire N__4928;
    wire N__4927;
    wire N__4926;
    wire N__4923;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4903;
    wire N__4898;
    wire N__4895;
    wire N__4888;
    wire N__4867;
    wire N__4866;
    wire N__4863;
    wire N__4862;
    wire N__4859;
    wire N__4856;
    wire N__4855;
    wire N__4854;
    wire N__4851;
    wire N__4848;
    wire N__4845;
    wire N__4842;
    wire N__4839;
    wire N__4828;
    wire N__4827;
    wire N__4826;
    wire N__4825;
    wire N__4824;
    wire N__4821;
    wire N__4818;
    wire N__4815;
    wire N__4812;
    wire N__4809;
    wire N__4806;
    wire N__4805;
    wire N__4804;
    wire N__4803;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4789;
    wire N__4786;
    wire N__4781;
    wire N__4780;
    wire N__4779;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4767;
    wire N__4762;
    wire N__4757;
    wire N__4754;
    wire N__4741;
    wire N__4738;
    wire N__4735;
    wire N__4734;
    wire N__4731;
    wire N__4728;
    wire N__4723;
    wire N__4720;
    wire N__4717;
    wire N__4714;
    wire N__4713;
    wire N__4712;
    wire N__4711;
    wire N__4710;
    wire N__4709;
    wire N__4708;
    wire N__4707;
    wire N__4706;
    wire N__4703;
    wire N__4700;
    wire N__4697;
    wire N__4694;
    wire N__4691;
    wire N__4688;
    wire N__4685;
    wire N__4684;
    wire N__4681;
    wire N__4680;
    wire N__4677;
    wire N__4674;
    wire N__4671;
    wire N__4668;
    wire N__4661;
    wire N__4660;
    wire N__4659;
    wire N__4654;
    wire N__4647;
    wire N__4642;
    wire N__4641;
    wire N__4640;
    wire N__4635;
    wire N__4630;
    wire N__4629;
    wire N__4628;
    wire N__4627;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4613;
    wire N__4608;
    wire N__4603;
    wire N__4600;
    wire N__4597;
    wire N__4582;
    wire N__4581;
    wire N__4578;
    wire N__4577;
    wire N__4576;
    wire N__4573;
    wire N__4570;
    wire N__4567;
    wire N__4566;
    wire N__4565;
    wire N__4562;
    wire N__4559;
    wire N__4556;
    wire N__4553;
    wire N__4548;
    wire N__4545;
    wire N__4542;
    wire N__4533;
    wire N__4528;
    wire N__4525;
    wire N__4522;
    wire N__4519;
    wire N__4516;
    wire N__4513;
    wire N__4510;
    wire N__4507;
    wire N__4504;
    wire N__4501;
    wire N__4498;
    wire N__4495;
    wire N__4492;
    wire N__4489;
    wire N__4486;
    wire N__4483;
    wire N__4480;
    wire N__4477;
    wire N__4474;
    wire N__4471;
    wire N__4468;
    wire N__4465;
    wire N__4462;
    wire N__4459;
    wire N__4456;
    wire N__4453;
    wire N__4450;
    wire N__4447;
    wire N__4444;
    wire N__4441;
    wire N__4438;
    wire N__4435;
    wire N__4434;
    wire N__4433;
    wire N__4432;
    wire N__4431;
    wire N__4428;
    wire N__4425;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4405;
    wire N__4404;
    wire N__4401;
    wire N__4400;
    wire N__4397;
    wire N__4394;
    wire N__4391;
    wire N__4384;
    wire N__4381;
    wire N__4378;
    wire N__4375;
    wire N__4372;
    wire N__4369;
    wire N__4366;
    wire N__4363;
    wire N__4362;
    wire N__4359;
    wire N__4356;
    wire N__4351;
    wire N__4348;
    wire N__4347;
    wire N__4344;
    wire N__4341;
    wire N__4336;
    wire N__4333;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4321;
    wire N__4318;
    wire N__4317;
    wire N__4316;
    wire N__4315;
    wire N__4314;
    wire N__4307;
    wire N__4306;
    wire N__4305;
    wire N__4304;
    wire N__4301;
    wire N__4298;
    wire N__4295;
    wire N__4292;
    wire N__4287;
    wire N__4276;
    wire N__4273;
    wire N__4270;
    wire N__4267;
    wire N__4264;
    wire N__4261;
    wire N__4258;
    wire N__4255;
    wire N__4252;
    wire N__4249;
    wire N__4246;
    wire N__4243;
    wire N__4242;
    wire N__4241;
    wire N__4240;
    wire N__4239;
    wire N__4236;
    wire N__4233;
    wire N__4230;
    wire N__4225;
    wire N__4216;
    wire N__4213;
    wire N__4210;
    wire N__4207;
    wire N__4204;
    wire N__4201;
    wire N__4198;
    wire N__4195;
    wire N__4192;
    wire N__4189;
    wire N__4186;
    wire N__4183;
    wire N__4180;
    wire N__4177;
    wire N__4174;
    wire N__4171;
    wire N__4168;
    wire N__4165;
    wire N__4162;
    wire N__4159;
    wire N__4156;
    wire N__4153;
    wire N__4150;
    wire N__4147;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4135;
    wire N__4132;
    wire N__4131;
    wire N__4126;
    wire N__4123;
    wire N__4120;
    wire N__4117;
    wire N__4114;
    wire N__4111;
    wire N__4108;
    wire N__4105;
    wire N__4102;
    wire N__4099;
    wire N__4096;
    wire N__4093;
    wire N__4092;
    wire N__4091;
    wire N__4088;
    wire N__4083;
    wire N__4078;
    wire N__4075;
    wire N__4074;
    wire N__4073;
    wire N__4070;
    wire N__4069;
    wire N__4068;
    wire N__4067;
    wire N__4066;
    wire N__4065;
    wire N__4060;
    wire N__4055;
    wire N__4052;
    wire N__4047;
    wire N__4044;
    wire N__4033;
    wire N__4030;
    wire N__4029;
    wire N__4028;
    wire N__4023;
    wire N__4020;
    wire N__4019;
    wire N__4018;
    wire N__4017;
    wire N__4016;
    wire N__4015;
    wire N__4014;
    wire N__4013;
    wire N__4012;
    wire N__4009;
    wire N__4006;
    wire N__4003;
    wire N__3998;
    wire N__3995;
    wire N__3988;
    wire N__3985;
    wire N__3976;
    wire N__3967;
    wire N__3966;
    wire N__3965;
    wire N__3960;
    wire N__3959;
    wire N__3958;
    wire N__3955;
    wire N__3952;
    wire N__3951;
    wire N__3950;
    wire N__3949;
    wire N__3948;
    wire N__3945;
    wire N__3944;
    wire N__3941;
    wire N__3938;
    wire N__3935;
    wire N__3930;
    wire N__3927;
    wire N__3924;
    wire N__3919;
    wire N__3904;
    wire N__3901;
    wire N__3898;
    wire N__3895;
    wire N__3892;
    wire N__3889;
    wire N__3886;
    wire N__3883;
    wire N__3880;
    wire N__3877;
    wire N__3874;
    wire N__3873;
    wire N__3870;
    wire N__3869;
    wire N__3866;
    wire N__3863;
    wire N__3860;
    wire N__3853;
    wire N__3850;
    wire N__3847;
    wire N__3846;
    wire N__3845;
    wire N__3842;
    wire N__3839;
    wire N__3836;
    wire N__3829;
    wire N__3826;
    wire N__3823;
    wire N__3820;
    wire N__3817;
    wire N__3814;
    wire N__3811;
    wire N__3808;
    wire N__3805;
    wire N__3804;
    wire N__3801;
    wire N__3798;
    wire N__3793;
    wire N__3790;
    wire N__3787;
    wire N__3784;
    wire N__3781;
    wire N__3778;
    wire N__3775;
    wire N__3772;
    wire N__3769;
    wire N__3766;
    wire N__3763;
    wire N__3760;
    wire N__3757;
    wire N__3754;
    wire N__3751;
    wire N__3748;
    wire N__3745;
    wire N__3744;
    wire N__3741;
    wire N__3738;
    wire N__3735;
    wire N__3732;
    wire N__3727;
    wire N__3724;
    wire N__3721;
    wire N__3718;
    wire N__3715;
    wire N__3714;
    wire N__3713;
    wire N__3712;
    wire N__3709;
    wire N__3706;
    wire N__3701;
    wire N__3696;
    wire N__3691;
    wire N__3688;
    wire N__3687;
    wire N__3686;
    wire N__3685;
    wire N__3682;
    wire N__3681;
    wire N__3676;
    wire N__3675;
    wire N__3672;
    wire N__3669;
    wire N__3666;
    wire N__3663;
    wire N__3660;
    wire N__3649;
    wire N__3648;
    wire N__3647;
    wire N__3646;
    wire N__3645;
    wire N__3644;
    wire N__3643;
    wire N__3642;
    wire N__3641;
    wire N__3640;
    wire N__3639;
    wire N__3638;
    wire N__3637;
    wire N__3636;
    wire N__3635;
    wire N__3634;
    wire N__3633;
    wire N__3632;
    wire N__3631;
    wire N__3630;
    wire N__3629;
    wire N__3628;
    wire N__3627;
    wire N__3626;
    wire N__3625;
    wire N__3624;
    wire N__3623;
    wire N__3568;
    wire N__3565;
    wire N__3562;
    wire N__3559;
    wire N__3556;
    wire N__3553;
    wire N__3550;
    wire N__3547;
    wire N__3546;
    wire N__3543;
    wire N__3540;
    wire N__3535;
    wire N__3532;
    wire N__3529;
    wire N__3526;
    wire N__3523;
    wire N__3520;
    wire N__3517;
    wire N__3516;
    wire N__3511;
    wire N__3508;
    wire N__3505;
    wire N__3502;
    wire N__3501;
    wire N__3498;
    wire N__3495;
    wire N__3490;
    wire N__3487;
    wire N__3484;
    wire N__3481;
    wire N__3478;
    wire N__3475;
    wire N__3472;
    wire N__3471;
    wire N__3468;
    wire N__3465;
    wire N__3460;
    wire N__3457;
    wire N__3454;
    wire N__3451;
    wire N__3448;
    wire N__3445;
    wire N__3444;
    wire N__3443;
    wire N__3440;
    wire N__3435;
    wire N__3430;
    wire N__3427;
    wire N__3424;
    wire N__3423;
    wire N__3420;
    wire N__3417;
    wire N__3412;
    wire N__3409;
    wire N__3408;
    wire N__3405;
    wire N__3402;
    wire N__3399;
    wire N__3394;
    wire N__3393;
    wire N__3390;
    wire N__3387;
    wire N__3382;
    wire N__3381;
    wire N__3378;
    wire N__3375;
    wire N__3372;
    wire N__3367;
    wire N__3366;
    wire N__3365;
    wire N__3362;
    wire N__3359;
    wire N__3356;
    wire N__3349;
    wire N__3346;
    wire N__3345;
    wire N__3344;
    wire N__3343;
    wire N__3342;
    wire N__3341;
    wire N__3340;
    wire N__3339;
    wire N__3336;
    wire N__3331;
    wire N__3328;
    wire N__3319;
    wire N__3310;
    wire N__3309;
    wire N__3308;
    wire N__3305;
    wire N__3300;
    wire N__3295;
    wire N__3292;
    wire N__3289;
    wire N__3288;
    wire N__3285;
    wire N__3282;
    wire N__3277;
    wire N__3276;
    wire N__3275;
    wire N__3272;
    wire N__3271;
    wire N__3266;
    wire N__3263;
    wire N__3260;
    wire N__3253;
    wire N__3252;
    wire N__3249;
    wire N__3246;
    wire N__3243;
    wire N__3238;
    wire N__3237;
    wire N__3234;
    wire N__3231;
    wire N__3226;
    wire N__3223;
    wire N__3220;
    wire N__3217;
    wire N__3214;
    wire N__3211;
    wire N__3208;
    wire N__3207;
    wire N__3204;
    wire N__3201;
    wire N__3198;
    wire N__3193;
    wire N__3190;
    wire N__3187;
    wire N__3186;
    wire N__3183;
    wire N__3180;
    wire N__3175;
    wire N__3172;
    wire N__3169;
    wire N__3166;
    wire N__3163;
    wire N__3160;
    wire N__3157;
    wire N__3154;
    wire N__3153;
    wire N__3152;
    wire N__3149;
    wire N__3144;
    wire N__3139;
    wire N__3136;
    wire N__3133;
    wire N__3130;
    wire N__3127;
    wire N__3124;
    wire N__3121;
    wire N__3118;
    wire N__3115;
    wire N__3112;
    wire N__3109;
    wire N__3106;
    wire N__3103;
    wire N__3100;
    wire N__3097;
    wire N__3094;
    wire N__3091;
    wire N__3088;
    wire N__3085;
    wire N__3082;
    wire N__3081;
    wire N__3080;
    wire N__3079;
    wire N__3078;
    wire N__3077;
    wire N__3074;
    wire N__3071;
    wire N__3062;
    wire N__3055;
    wire N__3054;
    wire N__3053;
    wire N__3050;
    wire N__3049;
    wire N__3048;
    wire N__3045;
    wire N__3042;
    wire N__3039;
    wire N__3032;
    wire N__3029;
    wire N__3022;
    wire N__3021;
    wire N__3018;
    wire N__3015;
    wire N__3010;
    wire N__3009;
    wire N__3006;
    wire N__3003;
    wire N__2998;
    wire N__2995;
    wire N__2992;
    wire N__2991;
    wire N__2986;
    wire N__2983;
    wire N__2980;
    wire N__2977;
    wire N__2974;
    wire N__2971;
    wire N__2968;
    wire N__2965;
    wire N__2962;
    wire N__2961;
    wire N__2960;
    wire N__2959;
    wire N__2958;
    wire N__2955;
    wire N__2954;
    wire N__2951;
    wire N__2948;
    wire N__2939;
    wire N__2932;
    wire N__2929;
    wire N__2926;
    wire N__2923;
    wire N__2922;
    wire N__2919;
    wire N__2916;
    wire N__2913;
    wire N__2910;
    wire N__2905;
    wire N__2902;
    wire N__2899;
    wire N__2896;
    wire N__2893;
    wire N__2890;
    wire N__2887;
    wire N__2884;
    wire N__2881;
    wire N__2878;
    wire N__2875;
    wire N__2872;
    wire N__2869;
    wire N__2866;
    wire N__2863;
    wire N__2860;
    wire N__2857;
    wire N__2854;
    wire N__2851;
    wire N__2848;
    wire N__2845;
    wire N__2842;
    wire N__2839;
    wire N__2836;
    wire N__2833;
    wire N__2830;
    wire N__2827;
    wire N__2824;
    wire N__2821;
    wire N__2818;
    wire N__2815;
    wire N__2812;
    wire N__2809;
    wire N__2806;
    wire N__2803;
    wire N__2800;
    wire N__2797;
    wire N__2794;
    wire N__2791;
    wire N__2788;
    wire N__2785;
    wire N__2782;
    wire N__2779;
    wire N__2776;
    wire N__2773;
    wire N__2770;
    wire N__2767;
    wire N__2764;
    wire N__2761;
    wire N__2758;
    wire N__2755;
    wire N__2752;
    wire N__2749;
    wire N__2746;
    wire N__2743;
    wire N__2740;
    wire N__2737;
    wire N__2734;
    wire N__2731;
    wire N__2728;
    wire N__2725;
    wire N__2722;
    wire N__2719;
    wire N__2716;
    wire N__2713;
    wire N__2710;
    wire N__2707;
    wire N__2706;
    wire N__2703;
    wire N__2700;
    wire N__2695;
    wire N__2692;
    wire N__2689;
    wire N__2686;
    wire N__2683;
    wire N__2680;
    wire N__2677;
    wire N__2674;
    wire N__2671;
    wire N__2668;
    wire N__2667;
    wire N__2664;
    wire N__2661;
    wire N__2656;
    wire N__2653;
    wire N__2650;
    wire N__2647;
    wire N__2644;
    wire N__2641;
    wire N__2638;
    wire N__2635;
    wire N__2632;
    wire N__2629;
    wire N__2626;
    wire N__2623;
    wire N__2620;
    wire N__2617;
    wire N__2614;
    wire N__2611;
    wire N__2608;
    wire N__2605;
    wire N__2602;
    wire N__2599;
    wire N__2596;
    wire N__2593;
    wire N__2590;
    wire N__2587;
    wire N__2584;
    wire N__2581;
    wire N__2578;
    wire N__2575;
    wire N__2572;
    wire N__2569;
    wire CLK40_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire RESETn_c_i;
    wire A_c_30;
    wire A_c_29;
    wire A_c_28;
    wire A_c_27;
    wire \U400_SDRAM.TA_COUNTER_7_f1_0_0_cascade_ ;
    wire \U400_SDRAM.un1_TA_COUNTER26_0_cascade_ ;
    wire \U400_SDRAM.TA_COUNTER23_cascade_ ;
    wire \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0 ;
    wire \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0_cascade_ ;
    wire \U400_SDRAM.CO1 ;
    wire \U400_SDRAM.CO1_cascade_ ;
    wire A_c_21;
    wire BANK0_c;
    wire A_c_22;
    wire BANK1_c;
    wire \INVU400_SDRAM.BANK0C_net ;
    wire \U400_SDRAM.un1_SDRAM_COUNTER52_4_0_i_a3_0_cascade_ ;
    wire \U400_SDRAM.un1_SDRAM_COUNTER52_4_0_i_1 ;
    wire \U400_SDRAM.N_208_cascade_ ;
    wire \U400_SDRAM.un1_SDRAM_COUNTER52_4_0_i_2 ;
    wire RASn_c;
    wire CASn_c;
    wire WEn_c;
    wire \INVU400_SDRAM.RASnC_net ;
    wire A_c_24;
    wire A_c_18;
    wire MA_c_8;
    wire A_c_17;
    wire A_c_9;
    wire MA_c_7;
    wire \INVU400_SDRAM.MA_8C_net ;
    wire A_c_8;
    wire A_c_16;
    wire MA_c_6;
    wire \INVU400_SDRAM.MA_6C_net ;
    wire bfn_5_3_0_;
    wire \U400_SDRAM.un2_REFRESH_COUNTER_cry_1 ;
    wire \U400_SDRAM.un2_REFRESH_COUNTER_cry_2 ;
    wire \U400_SDRAM.un2_REFRESH_COUNTER_cry_3 ;
    wire \U400_SDRAM.un2_REFRESH_COUNTER_cry_4 ;
    wire \U400_SDRAM.un2_REFRESH_COUNTER_cry_5 ;
    wire \U400_SDRAM.un2_REFRESH_COUNTER_cry_6 ;
    wire \U400_SDRAM.un2_REFRESH_COUNTER_cry_7 ;
    wire \INVU400_SDRAM.REFRESH_COUNTER_2C_net ;
    wire \U400_SDRAM.TA_COUNTERZ0Z_2 ;
    wire \U400_SDRAM.un1_TA_COUNTER26_2_0 ;
    wire TA_OUT;
    wire \U400_SDRAM.TA_COUNTERZ0Z_1 ;
    wire \U400_SDRAM.TA_COUNTERZ0Z_3 ;
    wire \U400_SDRAM.TA_COUNTER_0_sqmuxa ;
    wire \U400_SDRAM.TA_COUNTER27 ;
    wire \U400_SDRAM.TA_COUNTER_0_sqmuxa_cascade_ ;
    wire \INVU400_SDRAM.BURSTC_net ;
    wire \U400_SDRAM.un1_SDRAM_COUNTER52_2_0_i_1_cascade_ ;
    wire \U400_SDRAM.N_23 ;
    wire \U400_SDRAM.N_255 ;
    wire \U400_SDRAM.TACK_7_iv_i_i_0_cascade_ ;
    wire \U400_SDRAM.TACK_7_iv_i_i_1 ;
    wire \U400_SDRAM.N_15 ;
    wire \U400_SDRAM.RAM_CYCLE_e_1 ;
    wire \U400_SDRAM.N_6 ;
    wire RnW_c;
    wire \INVU400_SDRAM.RAM_CYCLEC_net ;
    wire CS0n_c;
    wire A_c_19;
    wire MA_c_9;
    wire \INVU400_SDRAM.CS0_ENC_net ;
    wire \INVU400_SDRAM.REFRESH_COUNTER_0C_net ;
    wire \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2Z0Z_1 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_2 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U400_SDRAM.TA_COUNTERZ0Z_0 ;
    wire \U400_SDRAM.BURSTZ0 ;
    wire \U400_SDRAM.TA_EN11_m ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_0 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U400_SDRAM.N_205_cascade_ ;
    wire \INVU400_SDRAM.SDRAM_CMD_1C_net ;
    wire \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en ;
    wire \U400_SDRAM.un1_REFRESH_COUNTERlto7_4 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_8 ;
    wire \U400_SDRAM.un1_REFRESH_COUNTERlto7_5 ;
    wire \U400_SDRAM.N_189 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_1_32_i_0_i_1_1_cascade_ ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_1_32_i_0_i_1_cascade_ ;
    wire \INVU400_SDRAM.SDRAM_CMD_0C_net ;
    wire \U400_SDRAM.N_128 ;
    wire \U400_SDRAM.N_185 ;
    wire \U400_SDRAM.RAM_CYCLEZ0 ;
    wire \U400_SDRAM.N_75_cascade_ ;
    wire \U400_SDRAM.CS1_EN_0 ;
    wire \U400_SDRAM.CS1_EN_7_i_0_o3_0_cascade_ ;
    wire \U400_SDRAM.N_159 ;
    wire A_c_23;
    wire \U400_SDRAM.CS0_ENZ0 ;
    wire \U400_SDRAM.N_159_cascade_ ;
    wire \U400_SDRAM.N_75 ;
    wire \U400_SDRAM.CS0_EN_0 ;
    wire \U400_SDRAM.N_250 ;
    wire \U400_SDRAM.N_176_cascade_ ;
    wire \U400_SDRAM.CS1_ENZ0 ;
    wire CS1n_c;
    wire A_c_26;
    wire MA_c_12;
    wire \INVU400_SDRAM.CS1nC_net ;
    wire CONSTANT_ONE_NET;
    wire UUBEn_c;
    wire \U400_SDRAM.TA_COUNTER23 ;
    wire \U400_SDRAM.TACKZ0 ;
    wire CLK40_c_g;
    wire \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en_0 ;
    wire \U400_SDRAM.N_252_cascade_ ;
    wire \U400_SDRAM.N_200_cascade_ ;
    wire \U400_SDRAM.N_199 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_61_i_i_1_cascade_ ;
    wire \U400_SDRAM.N_17 ;
    wire \INVU400_SDRAM.SDRAM_CMD_2C_net ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_i_a2_0_1_1 ;
    wire \U400_SDRAM.N_228 ;
    wire \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5Z0Z_0_cascade_ ;
    wire \INVU400_SDRAM.SDRAM_COUNTER_3C_net ;
    wire \U400_SDRAM.N_203 ;
    wire \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_i_0 ;
    wire \U400_SDRAM.N_126_cascade_ ;
    wire \U400_SDRAM.N_129_cascade_ ;
    wire \U400_SDRAM.N_257_cascade_ ;
    wire \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_1_0 ;
    wire \U400_SDRAM.N_133 ;
    wire \U400_SDRAM.N_133_cascade_ ;
    wire \U400_SDRAM.N_139 ;
    wire \U400_SDRAM.N_141_cascade_ ;
    wire \U400_SDRAM.REFRESH_COUNTER_RNIVV903Z0Z_8 ;
    wire \U400_SDRAM.RAM_CYCLE_STARTZ0 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_2_0 ;
    wire \U400_SDRAM.SDRAM_COUNTER_s_0 ;
    wire \U400_SDRAM.N_181_cascade_ ;
    wire \INVU400_SDRAM.SDRAM_COUNTER_0C_net ;
    wire A_c_25;
    wire MA_c_11;
    wire \U400_SDRAM.N_257 ;
    wire \INVU400_SDRAM.MA_11C_net ;
    wire A_c_6;
    wire A_c_14;
    wire MA_c_4;
    wire MA_c_5;
    wire \INVU400_SDRAM.MA_4C_net ;
    wire \U400_SDRAM.N_150 ;
    wire \U400_SDRAM.N_150_cascade_ ;
    wire \U400_SDRAM.N_252 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_61_i_i_a3_1_0_cascade_ ;
    wire \U400_SDRAM.N_201 ;
    wire TA_EN_i_ess;
    wire N_529_i;
    wire \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5Z0Z_0 ;
    wire \INVU400_SDRAM.SDRAM_COUNTER_1C_net ;
    wire \U400_SDRAM.N_129 ;
    wire \U400_SDRAM.N_260 ;
    wire bfn_8_8_0_;
    wire \U400_SDRAM.SDRAM_COUNTER_s_1 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_0 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_1 ;
    wire \U400_SDRAM.SDRAM_COUNTER_s_3 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_2 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_3 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_4 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_5 ;
    wire \U400_SDRAM.N_37 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_6 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_7 ;
    wire \INVU400_SDRAM.SDRAM_COUNTER_2C_net ;
    wire \U400_SDRAM.SDRAM_COUNTERe_0_i ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U400_SDRAM.WRITE_CYCLEZ0 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U400_SDRAM.N_161_cascade_ ;
    wire \U400_SDRAM.N_183 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U400_SDRAM.N_126 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U400_SDRAM.N_138 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_a3_1_0_0 ;
    wire \U400_SDRAM.SDRAM_CONFIGUREDZ0 ;
    wire \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7JZ0 ;
    wire A_c_7;
    wire A_c_15;
    wire \U400_SDRAM.MAc_0_0 ;
    wire A_c_2;
    wire A_c_10;
    wire MA_c_0;
    wire A_c_20;
    wire MA_c_10;
    wire \INVU400_SDRAM.MA_0C_net ;
    wire UMBEn_c;
    wire LLBEn_c;
    wire A_c_1;
    wire A_c_0;
    wire LMBEn_c;
    wire TSn_c;
    wire \U400_SDRAM.N_220 ;
    wire SIZ_c_1;
    wire SIZ_c_0;
    wire \U400_SDRAM.BURST8 ;
    wire A_c_31;
    wire U400_ADDRESS_DECODE_RAM_SPACE_0_a3_3;
    wire RESETn_c;
    wire N_220_3_i;
    wire A_c_5;
    wire A_c_13;
    wire MA_c_3;
    wire \INVU400_SDRAM.MA_3C_net ;
    wire A_c_3;
    wire A_c_11;
    wire A_c_4;
    wire A_c_12;
    wire \U400_SDRAM.MAc_1_0 ;
    wire MA_c_2;
    wire \U400_SDRAM.SDRAM_CMDZ0Z_1 ;
    wire \U400_SDRAM.SDRAM_CMDZ1Z_0 ;
    wire \U400_SDRAM.SDRAM_CMDZ0Z_2 ;
    wire \U400_SDRAM.MAc_9_0 ;
    wire MA_c_1;
    wire _gnd_net_;
    wire \INVU400_SDRAM.MA_2C_net ;
    wire RESETn_c_i_g;

    IO_PAD MA_obuf_7_iopad (
            .OE(N__7004),
            .DIN(N__7003),
            .DOUT(N__7002),
            .PACKAGEPIN(MA[7]));
    defparam MA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_7_preio (
            .PADOEN(N__7004),
            .PADOUT(N__7003),
            .PADIN(N__7002),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2797),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__6995),
            .DIN(N__6994),
            .DOUT(N__6993),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__6995),
            .PADOUT(N__6994),
            .PADIN(N__6993),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__6986),
            .DIN(N__6985),
            .DOUT(N__6984),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__6986),
            .PADOUT(N__6985),
            .PADIN(N__6984),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2881),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__6977),
            .DIN(N__6976),
            .DOUT(N__6975),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__6977),
            .PADOUT(N__6976),
            .PADIN(N__6975),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2677),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_8_iopad (
            .OE(N__6968),
            .DIN(N__6967),
            .DOUT(N__6966),
            .PACKAGEPIN(MA[8]));
    defparam MA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_8_preio (
            .PADOEN(N__6968),
            .PADOUT(N__6967),
            .PADIN(N__6966),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2830),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_10_iopad (
            .OE(N__6959),
            .DIN(N__6958),
            .DOUT(N__6957),
            .PACKAGEPIN(MA[10]));
    defparam MA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_10_preio (
            .PADOEN(N__6959),
            .PADOUT(N__6958),
            .PADIN(N__6957),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5881),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_23_iopad (
            .OE(N__6950),
            .DIN(N__6949),
            .DOUT(N__6948),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__6950),
            .PADOUT(N__6949),
            .PADIN(N__6948),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_2_iopad (
            .OE(N__6941),
            .DIN(N__6940),
            .DOUT(N__6939),
            .PACKAGEPIN(MA[2]));
    defparam MA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_2_preio (
            .PADOEN(N__6941),
            .PADOUT(N__6940),
            .PADIN(N__6939),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6325),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__6932),
            .DIN(N__6931),
            .DOUT(N__6930),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__6932),
            .PADOUT(N__6931),
            .PADIN(N__6930),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__6923),
            .DIN(N__6922),
            .DOUT(N__6921),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__6923),
            .PADOUT(N__6922),
            .PADIN(N__6921),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__6914),
            .DIN(N__6913),
            .DOUT(N__6912),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__6914),
            .PADOUT(N__6913),
            .PADIN(N__6912),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3727),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_24_iopad (
            .OE(N__6905),
            .DIN(N__6904),
            .DOUT(N__6903),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__6905),
            .PADOUT(N__6904),
            .PADIN(N__6903),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_31_iopad (
            .OE(N__6896),
            .DIN(N__6895),
            .DOUT(N__6894),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__6896),
            .PADOUT(N__6895),
            .PADIN(N__6894),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__6887),
            .DIN(N__6886),
            .DOUT(N__6885),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__6887),
            .PADOUT(N__6886),
            .PADIN(N__6885),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_12_iopad (
            .OE(N__6878),
            .DIN(N__6877),
            .DOUT(N__6876),
            .PACKAGEPIN(MA[12]));
    defparam MA_obuf_12_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_12_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_12_preio (
            .PADOEN(N__6878),
            .PADOUT(N__6877),
            .PADIN(N__6876),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3763),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_1_iopad (
            .OE(N__6869),
            .DIN(N__6868),
            .DOUT(N__6867),
            .PACKAGEPIN(MA[1]));
    defparam MA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_1_preio (
            .PADOEN(N__6869),
            .PADOUT(N__6868),
            .PADIN(N__6867),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5947),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__6860),
            .DIN(N__6859),
            .DOUT(N__6858),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__6860),
            .PADOUT(N__6859),
            .PADIN(N__6858),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__6851),
            .DIN(N__6850),
            .DOUT(N__6849),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__6851),
            .PADOUT(N__6850),
            .PADIN(N__6849),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_21_iopad (
            .OE(N__6842),
            .DIN(N__6841),
            .DOUT(N__6840),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__6842),
            .PADOUT(N__6841),
            .PADIN(N__6840),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_4_iopad (
            .OE(N__6833),
            .DIN(N__6832),
            .DOUT(N__6831),
            .PACKAGEPIN(MA[4]));
    defparam MA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_4_preio (
            .PADOEN(N__6833),
            .PADOUT(N__6832),
            .PADIN(N__6831),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4186),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__6824),
            .DIN(N__6823),
            .DOUT(N__6822),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__6824),
            .PADOUT(N__6823),
            .PADIN(N__6822),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__6815),
            .DIN(N__6814),
            .DOUT(N__6813),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__6815),
            .PADOUT(N__6814),
            .PADIN(N__6813),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__6806),
            .DIN(N__6805),
            .DOUT(N__6804),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__6806),
            .PADOUT(N__6805),
            .PADIN(N__6804),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5866),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__6797),
            .DIN(N__6796),
            .DOUT(N__6795),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__6797),
            .PADOUT(N__6796),
            .PADIN(N__6795),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_9_iopad (
            .OE(N__6788),
            .DIN(N__6787),
            .DOUT(N__6786),
            .PACKAGEPIN(MA[9]));
    defparam MA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_9_preio (
            .PADOEN(N__6788),
            .PADOUT(N__6787),
            .PADIN(N__6786),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3091),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__6779),
            .DIN(N__6778),
            .DOUT(N__6777),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__6779),
            .PADOUT(N__6778),
            .PADIN(N__6777),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5875),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__6770),
            .DIN(N__6769),
            .DOUT(N__6768),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__6770),
            .PADOUT(N__6769),
            .PADIN(N__6768),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_29_iopad (
            .OE(N__6761),
            .DIN(N__6760),
            .DOUT(N__6759),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__6761),
            .PADOUT(N__6760),
            .PADIN(N__6759),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__6752),
            .DIN(N__6751),
            .DOUT(N__6750),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__6752),
            .PADOUT(N__6751),
            .PADIN(N__6750),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3751),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__6743),
            .DIN(N__6742),
            .DOUT(N__6741),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__6743),
            .PADOUT(N__6742),
            .PADIN(N__6741),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_22_iopad (
            .OE(N__6734),
            .DIN(N__6733),
            .DOUT(N__6732),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__6734),
            .PADOUT(N__6733),
            .PADIN(N__6732),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_3_iopad (
            .OE(N__6725),
            .DIN(N__6724),
            .DOUT(N__6723),
            .PACKAGEPIN(MA[3]));
    defparam MA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_3_preio (
            .PADOEN(N__6725),
            .PADOUT(N__6724),
            .PADIN(N__6723),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5371),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__6716),
            .DIN(N__6715),
            .DOUT(N__6714),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__6716),
            .PADOUT(N__6715),
            .PADIN(N__6714),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__6707),
            .DIN(N__6706),
            .DOUT(N__6705),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__6707),
            .PADOUT(N__6706),
            .PADIN(N__6705),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_27_iopad (
            .OE(N__6698),
            .DIN(N__6697),
            .DOUT(N__6696),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__6698),
            .PADOUT(N__6697),
            .PADIN(N__6696),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_6_iopad (
            .OE(N__6689),
            .DIN(N__6688),
            .DOUT(N__6687),
            .PACKAGEPIN(MA[6]));
    defparam MA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_6_preio (
            .PADOEN(N__6689),
            .PADOUT(N__6688),
            .PADIN(N__6687),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2761),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__6680),
            .DIN(N__6679),
            .DOUT(N__6678),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__6680),
            .PADOUT(N__6679),
            .PADIN(N__6678),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__6671),
            .DIN(N__6670),
            .DOUT(N__6669),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__6671),
            .PADOUT(N__6670),
            .PADIN(N__6669),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__6662),
            .DIN(N__6661),
            .DOUT(N__6660),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__6662),
            .PADOUT(N__6661),
            .PADIN(N__6660),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__6653),
            .DIN(N__6652),
            .DOUT(N__6651),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__6653),
            .PADOUT(N__6652),
            .PADIN(N__6651),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2893),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__6644),
            .DIN(N__6643),
            .DOUT(N__6642),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__6644),
            .PADOUT(N__6643),
            .PADIN(N__6642),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__6635),
            .DIN(N__6634),
            .DOUT(N__6633),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__6635),
            .PADOUT(N__6634),
            .PADIN(N__6633),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2716),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_11_iopad (
            .OE(N__6626),
            .DIN(N__6625),
            .DOUT(N__6624),
            .PACKAGEPIN(MA[11]));
    defparam MA_obuf_11_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_11_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_11_preio (
            .PADOEN(N__6626),
            .PADOUT(N__6625),
            .PADIN(N__6624),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4258),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TAn_obuft_iopad (
            .OE(N__6617),
            .DIN(N__6616),
            .DOUT(N__6615),
            .PACKAGEPIN(TAn));
    defparam TAn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TAn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TAn_obuft_preio (
            .PADOEN(N__6617),
            .PADOUT(N__6616),
            .PADIN(N__6615),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4117),
            .DIN0(),
            .DOUT0(N__2926),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__6608),
            .DIN(N__6607),
            .DOUT(N__6606),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__6608),
            .PADOUT(N__6607),
            .PADIN(N__6606),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_5_iopad (
            .OE(N__6599),
            .DIN(N__6598),
            .DOUT(N__6597),
            .PACKAGEPIN(MA[5]));
    defparam MA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_5_preio (
            .PADOEN(N__6599),
            .PADOUT(N__6598),
            .PADIN(N__6597),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4171),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__6590),
            .DIN(N__6589),
            .DOUT(N__6588),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__6590),
            .PADOUT(N__6589),
            .PADIN(N__6588),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__6581),
            .DIN(N__6580),
            .DOUT(N__6579),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__6581),
            .PADOUT(N__6580),
            .PADIN(N__6579),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam LBENn_obuf_iopad.PULLUP=1'b1;
    IO_PAD LBENn_obuf_iopad (
            .OE(N__6572),
            .DIN(N__6571),
            .DOUT(N__6570),
            .PACKAGEPIN(LBENn));
    defparam LBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LBENn_obuf_preio (
            .PADOEN(N__6572),
            .PADOUT(N__6571),
            .PADIN(N__6570),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5404),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_25_iopad (
            .OE(N__6563),
            .DIN(N__6562),
            .DOUT(N__6561),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__6563),
            .PADOUT(N__6562),
            .PADIN(N__6561),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CS1n_obuf_iopad (
            .OE(N__6554),
            .DIN(N__6553),
            .DOUT(N__6552),
            .PACKAGEPIN(CS1n));
    defparam CS1n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CS1n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CS1n_obuf_preio (
            .PADOEN(N__6554),
            .PADOUT(N__6553),
            .PADIN(N__6552),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3793),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__6545),
            .DIN(N__6544),
            .DOUT(N__6543),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__6545),
            .PADOUT(N__6544),
            .PADIN(N__6543),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_28_iopad (
            .OE(N__6536),
            .DIN(N__6535),
            .DOUT(N__6534),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__6536),
            .PADOUT(N__6535),
            .PADIN(N__6534),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_30_iopad (
            .OE(N__6527),
            .DIN(N__6526),
            .DOUT(N__6525),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__6527),
            .PADOUT(N__6526),
            .PADIN(N__6525),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__6518),
            .DIN(N__6517),
            .DOUT(N__6516),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__6518),
            .PADOUT(N__6517),
            .PADIN(N__6516),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__6509),
            .DIN(N__6508),
            .DOUT(N__6507),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__6509),
            .PADOUT(N__6508),
            .PADIN(N__6507),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2872),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_0_iopad (
            .OE(N__6500),
            .DIN(N__6499),
            .DOUT(N__6498),
            .PACKAGEPIN(MA[0]));
    defparam MA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_0_preio (
            .PADOEN(N__6500),
            .PADOUT(N__6499),
            .PADIN(N__6498),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4468),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__6491),
            .DIN(N__6490),
            .DOUT(N__6489),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__6491),
            .PADOUT(N__6490),
            .PADIN(N__6489),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__6482),
            .DIN(N__6481),
            .DOUT(N__6480),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__6482),
            .PADOUT(N__6481),
            .PADIN(N__6480),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__6473),
            .DIN(N__6472),
            .DOUT(N__6471),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__6473),
            .PADOUT(N__6472),
            .PADIN(N__6471),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CS0n_obuf_iopad (
            .OE(N__6464),
            .DIN(N__6463),
            .DOUT(N__6462),
            .PACKAGEPIN(CS0n));
    defparam CS0n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CS0n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CS0n_obuf_preio (
            .PADOEN(N__6464),
            .PADOUT(N__6463),
            .PADIN(N__6462),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3124),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_26_iopad (
            .OE(N__6455),
            .DIN(N__6454),
            .DOUT(N__6453),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__6455),
            .PADOUT(N__6454),
            .PADIN(N__6453),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__6446),
            .DIN(N__6445),
            .DOUT(N__6444),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__6446),
            .PADOUT(N__6445),
            .PADIN(N__6444),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5785),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__6437),
            .DIN(N__6436),
            .DOUT(N__6435),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__6437),
            .PADOUT(N__6436),
            .PADIN(N__6435),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_ibuf_gb_io_iopad (
            .OE(N__6428),
            .DIN(N__6427),
            .DOUT(N__6426),
            .PACKAGEPIN(CLK40));
    defparam CLK40_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_ibuf_gb_io_preio (
            .PADOEN(N__6428),
            .PADOUT(N__6427),
            .PADIN(N__6426),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1516 (
            .O(N__6409),
            .I(N__6406));
    LocalMux I__1515 (
            .O(N__6406),
            .I(N__6403));
    Span4Mux_s2_v I__1514 (
            .O(N__6403),
            .I(N__6400));
    IoSpan4Mux I__1513 (
            .O(N__6400),
            .I(N__6397));
    Odrv4 I__1512 (
            .O(N__6397),
            .I(A_c_4));
    CascadeMux I__1511 (
            .O(N__6394),
            .I(N__6391));
    InMux I__1510 (
            .O(N__6391),
            .I(N__6388));
    LocalMux I__1509 (
            .O(N__6388),
            .I(A_c_12));
    InMux I__1508 (
            .O(N__6385),
            .I(N__6380));
    InMux I__1507 (
            .O(N__6384),
            .I(N__6377));
    InMux I__1506 (
            .O(N__6383),
            .I(N__6372));
    LocalMux I__1505 (
            .O(N__6380),
            .I(N__6367));
    LocalMux I__1504 (
            .O(N__6377),
            .I(N__6367));
    InMux I__1503 (
            .O(N__6376),
            .I(N__6364));
    InMux I__1502 (
            .O(N__6375),
            .I(N__6361));
    LocalMux I__1501 (
            .O(N__6372),
            .I(N__6356));
    Span4Mux_h I__1500 (
            .O(N__6367),
            .I(N__6351));
    LocalMux I__1499 (
            .O(N__6364),
            .I(N__6351));
    LocalMux I__1498 (
            .O(N__6361),
            .I(N__6348));
    InMux I__1497 (
            .O(N__6360),
            .I(N__6343));
    InMux I__1496 (
            .O(N__6359),
            .I(N__6343));
    Span4Mux_v I__1495 (
            .O(N__6356),
            .I(N__6338));
    Span4Mux_v I__1494 (
            .O(N__6351),
            .I(N__6338));
    Span4Mux_h I__1493 (
            .O(N__6348),
            .I(N__6335));
    LocalMux I__1492 (
            .O(N__6343),
            .I(N__6332));
    Odrv4 I__1491 (
            .O(N__6338),
            .I(\U400_SDRAM.MAc_1_0 ));
    Odrv4 I__1490 (
            .O(N__6335),
            .I(\U400_SDRAM.MAc_1_0 ));
    Odrv4 I__1489 (
            .O(N__6332),
            .I(\U400_SDRAM.MAc_1_0 ));
    IoInMux I__1488 (
            .O(N__6325),
            .I(N__6322));
    LocalMux I__1487 (
            .O(N__6322),
            .I(MA_c_2));
    CascadeMux I__1486 (
            .O(N__6319),
            .I(N__6315));
    InMux I__1485 (
            .O(N__6318),
            .I(N__6311));
    InMux I__1484 (
            .O(N__6315),
            .I(N__6308));
    InMux I__1483 (
            .O(N__6314),
            .I(N__6305));
    LocalMux I__1482 (
            .O(N__6311),
            .I(N__6292));
    LocalMux I__1481 (
            .O(N__6308),
            .I(N__6292));
    LocalMux I__1480 (
            .O(N__6305),
            .I(N__6289));
    InMux I__1479 (
            .O(N__6304),
            .I(N__6286));
    InMux I__1478 (
            .O(N__6303),
            .I(N__6283));
    InMux I__1477 (
            .O(N__6302),
            .I(N__6278));
    InMux I__1476 (
            .O(N__6301),
            .I(N__6278));
    InMux I__1475 (
            .O(N__6300),
            .I(N__6275));
    InMux I__1474 (
            .O(N__6299),
            .I(N__6272));
    InMux I__1473 (
            .O(N__6298),
            .I(N__6267));
    InMux I__1472 (
            .O(N__6297),
            .I(N__6267));
    Span4Mux_s2_v I__1471 (
            .O(N__6292),
            .I(N__6264));
    Span4Mux_s1_v I__1470 (
            .O(N__6289),
            .I(N__6257));
    LocalMux I__1469 (
            .O(N__6286),
            .I(N__6257));
    LocalMux I__1468 (
            .O(N__6283),
            .I(N__6257));
    LocalMux I__1467 (
            .O(N__6278),
            .I(N__6250));
    LocalMux I__1466 (
            .O(N__6275),
            .I(N__6250));
    LocalMux I__1465 (
            .O(N__6272),
            .I(N__6247));
    LocalMux I__1464 (
            .O(N__6267),
            .I(N__6244));
    Sp12to4 I__1463 (
            .O(N__6264),
            .I(N__6241));
    Span4Mux_h I__1462 (
            .O(N__6257),
            .I(N__6238));
    InMux I__1461 (
            .O(N__6256),
            .I(N__6235));
    InMux I__1460 (
            .O(N__6255),
            .I(N__6232));
    Span4Mux_v I__1459 (
            .O(N__6250),
            .I(N__6229));
    Span4Mux_v I__1458 (
            .O(N__6247),
            .I(N__6226));
    Sp12to4 I__1457 (
            .O(N__6244),
            .I(N__6217));
    Span12Mux_s6_h I__1456 (
            .O(N__6241),
            .I(N__6217));
    Sp12to4 I__1455 (
            .O(N__6238),
            .I(N__6217));
    LocalMux I__1454 (
            .O(N__6235),
            .I(N__6217));
    LocalMux I__1453 (
            .O(N__6232),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1452 (
            .O(N__6229),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1451 (
            .O(N__6226),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_1 ));
    Odrv12 I__1450 (
            .O(N__6217),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_1 ));
    InMux I__1449 (
            .O(N__6208),
            .I(N__6205));
    LocalMux I__1448 (
            .O(N__6205),
            .I(N__6200));
    InMux I__1447 (
            .O(N__6204),
            .I(N__6195));
    InMux I__1446 (
            .O(N__6203),
            .I(N__6192));
    Span4Mux_h I__1445 (
            .O(N__6200),
            .I(N__6185));
    InMux I__1444 (
            .O(N__6199),
            .I(N__6182));
    InMux I__1443 (
            .O(N__6198),
            .I(N__6179));
    LocalMux I__1442 (
            .O(N__6195),
            .I(N__6176));
    LocalMux I__1441 (
            .O(N__6192),
            .I(N__6173));
    InMux I__1440 (
            .O(N__6191),
            .I(N__6168));
    InMux I__1439 (
            .O(N__6190),
            .I(N__6168));
    InMux I__1438 (
            .O(N__6189),
            .I(N__6163));
    InMux I__1437 (
            .O(N__6188),
            .I(N__6163));
    Sp12to4 I__1436 (
            .O(N__6185),
            .I(N__6156));
    LocalMux I__1435 (
            .O(N__6182),
            .I(N__6156));
    LocalMux I__1434 (
            .O(N__6179),
            .I(N__6153));
    Span4Mux_s3_v I__1433 (
            .O(N__6176),
            .I(N__6150));
    Span4Mux_h I__1432 (
            .O(N__6173),
            .I(N__6143));
    LocalMux I__1431 (
            .O(N__6168),
            .I(N__6143));
    LocalMux I__1430 (
            .O(N__6163),
            .I(N__6143));
    InMux I__1429 (
            .O(N__6162),
            .I(N__6140));
    InMux I__1428 (
            .O(N__6161),
            .I(N__6137));
    Span12Mux_s10_v I__1427 (
            .O(N__6156),
            .I(N__6134));
    Span4Mux_h I__1426 (
            .O(N__6153),
            .I(N__6129));
    Span4Mux_v I__1425 (
            .O(N__6150),
            .I(N__6129));
    Sp12to4 I__1424 (
            .O(N__6143),
            .I(N__6124));
    LocalMux I__1423 (
            .O(N__6140),
            .I(N__6124));
    LocalMux I__1422 (
            .O(N__6137),
            .I(\U400_SDRAM.SDRAM_CMDZ1Z_0 ));
    Odrv12 I__1421 (
            .O(N__6134),
            .I(\U400_SDRAM.SDRAM_CMDZ1Z_0 ));
    Odrv4 I__1420 (
            .O(N__6129),
            .I(\U400_SDRAM.SDRAM_CMDZ1Z_0 ));
    Odrv12 I__1419 (
            .O(N__6124),
            .I(\U400_SDRAM.SDRAM_CMDZ1Z_0 ));
    CascadeMux I__1418 (
            .O(N__6115),
            .I(N__6110));
    CascadeMux I__1417 (
            .O(N__6114),
            .I(N__6105));
    InMux I__1416 (
            .O(N__6113),
            .I(N__6100));
    InMux I__1415 (
            .O(N__6110),
            .I(N__6097));
    InMux I__1414 (
            .O(N__6109),
            .I(N__6094));
    CascadeMux I__1413 (
            .O(N__6108),
            .I(N__6091));
    InMux I__1412 (
            .O(N__6105),
            .I(N__6082));
    InMux I__1411 (
            .O(N__6104),
            .I(N__6082));
    InMux I__1410 (
            .O(N__6103),
            .I(N__6079));
    LocalMux I__1409 (
            .O(N__6100),
            .I(N__6073));
    LocalMux I__1408 (
            .O(N__6097),
            .I(N__6073));
    LocalMux I__1407 (
            .O(N__6094),
            .I(N__6070));
    InMux I__1406 (
            .O(N__6091),
            .I(N__6065));
    InMux I__1405 (
            .O(N__6090),
            .I(N__6065));
    InMux I__1404 (
            .O(N__6089),
            .I(N__6060));
    InMux I__1403 (
            .O(N__6088),
            .I(N__6060));
    InMux I__1402 (
            .O(N__6087),
            .I(N__6057));
    LocalMux I__1401 (
            .O(N__6082),
            .I(N__6050));
    LocalMux I__1400 (
            .O(N__6079),
            .I(N__6050));
    InMux I__1399 (
            .O(N__6078),
            .I(N__6043));
    Span4Mux_v I__1398 (
            .O(N__6073),
            .I(N__6037));
    Span4Mux_s3_v I__1397 (
            .O(N__6070),
            .I(N__6037));
    LocalMux I__1396 (
            .O(N__6065),
            .I(N__6030));
    LocalMux I__1395 (
            .O(N__6060),
            .I(N__6030));
    LocalMux I__1394 (
            .O(N__6057),
            .I(N__6030));
    InMux I__1393 (
            .O(N__6056),
            .I(N__6026));
    InMux I__1392 (
            .O(N__6055),
            .I(N__6023));
    Span4Mux_s2_v I__1391 (
            .O(N__6050),
            .I(N__6020));
    InMux I__1390 (
            .O(N__6049),
            .I(N__6017));
    InMux I__1389 (
            .O(N__6048),
            .I(N__6012));
    InMux I__1388 (
            .O(N__6047),
            .I(N__6012));
    InMux I__1387 (
            .O(N__6046),
            .I(N__6009));
    LocalMux I__1386 (
            .O(N__6043),
            .I(N__6006));
    InMux I__1385 (
            .O(N__6042),
            .I(N__6003));
    Span4Mux_h I__1384 (
            .O(N__6037),
            .I(N__5998));
    Span4Mux_s3_v I__1383 (
            .O(N__6030),
            .I(N__5998));
    InMux I__1382 (
            .O(N__6029),
            .I(N__5995));
    LocalMux I__1381 (
            .O(N__6026),
            .I(N__5990));
    LocalMux I__1380 (
            .O(N__6023),
            .I(N__5990));
    Span4Mux_v I__1379 (
            .O(N__6020),
            .I(N__5987));
    LocalMux I__1378 (
            .O(N__6017),
            .I(N__5984));
    LocalMux I__1377 (
            .O(N__6012),
            .I(N__5975));
    LocalMux I__1376 (
            .O(N__6009),
            .I(N__5975));
    Span4Mux_h I__1375 (
            .O(N__6006),
            .I(N__5975));
    LocalMux I__1374 (
            .O(N__6003),
            .I(N__5975));
    Span4Mux_v I__1373 (
            .O(N__5998),
            .I(N__5972));
    LocalMux I__1372 (
            .O(N__5995),
            .I(N__5965));
    Span4Mux_v I__1371 (
            .O(N__5990),
            .I(N__5965));
    Span4Mux_v I__1370 (
            .O(N__5987),
            .I(N__5965));
    Span4Mux_h I__1369 (
            .O(N__5984),
            .I(N__5960));
    Span4Mux_v I__1368 (
            .O(N__5975),
            .I(N__5960));
    Odrv4 I__1367 (
            .O(N__5972),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1366 (
            .O(N__5965),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1365 (
            .O(N__5960),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    InMux I__1364 (
            .O(N__5953),
            .I(N__5950));
    LocalMux I__1363 (
            .O(N__5950),
            .I(\U400_SDRAM.MAc_9_0 ));
    IoInMux I__1362 (
            .O(N__5947),
            .I(N__5944));
    LocalMux I__1361 (
            .O(N__5944),
            .I(MA_c_1));
    InMux I__1360 (
            .O(N__5941),
            .I(N__5938));
    LocalMux I__1359 (
            .O(N__5938),
            .I(N__5929));
    SRMux I__1358 (
            .O(N__5937),
            .I(N__5887));
    SRMux I__1357 (
            .O(N__5936),
            .I(N__5887));
    SRMux I__1356 (
            .O(N__5935),
            .I(N__5887));
    SRMux I__1355 (
            .O(N__5934),
            .I(N__5887));
    SRMux I__1354 (
            .O(N__5933),
            .I(N__5887));
    SRMux I__1353 (
            .O(N__5932),
            .I(N__5887));
    Glb2LocalMux I__1352 (
            .O(N__5929),
            .I(N__5887));
    SRMux I__1351 (
            .O(N__5928),
            .I(N__5887));
    SRMux I__1350 (
            .O(N__5927),
            .I(N__5887));
    SRMux I__1349 (
            .O(N__5926),
            .I(N__5887));
    SRMux I__1348 (
            .O(N__5925),
            .I(N__5887));
    SRMux I__1347 (
            .O(N__5924),
            .I(N__5887));
    SRMux I__1346 (
            .O(N__5923),
            .I(N__5887));
    SRMux I__1345 (
            .O(N__5922),
            .I(N__5887));
    SRMux I__1344 (
            .O(N__5921),
            .I(N__5887));
    SRMux I__1343 (
            .O(N__5920),
            .I(N__5887));
    GlobalMux I__1342 (
            .O(N__5887),
            .I(N__5884));
    gio2CtrlBuf I__1341 (
            .O(N__5884),
            .I(RESETn_c_i_g));
    IoInMux I__1340 (
            .O(N__5881),
            .I(N__5878));
    LocalMux I__1339 (
            .O(N__5878),
            .I(MA_c_10));
    IoInMux I__1338 (
            .O(N__5875),
            .I(N__5872));
    LocalMux I__1337 (
            .O(N__5872),
            .I(N__5869));
    Odrv12 I__1336 (
            .O(N__5869),
            .I(UMBEn_c));
    IoInMux I__1335 (
            .O(N__5866),
            .I(N__5863));
    LocalMux I__1334 (
            .O(N__5863),
            .I(N__5860));
    Odrv4 I__1333 (
            .O(N__5860),
            .I(LLBEn_c));
    CascadeMux I__1332 (
            .O(N__5857),
            .I(N__5853));
    CascadeMux I__1331 (
            .O(N__5856),
            .I(N__5850));
    InMux I__1330 (
            .O(N__5853),
            .I(N__5842));
    InMux I__1329 (
            .O(N__5850),
            .I(N__5842));
    InMux I__1328 (
            .O(N__5849),
            .I(N__5842));
    LocalMux I__1327 (
            .O(N__5842),
            .I(N__5838));
    InMux I__1326 (
            .O(N__5841),
            .I(N__5835));
    Span4Mux_h I__1325 (
            .O(N__5838),
            .I(N__5832));
    LocalMux I__1324 (
            .O(N__5835),
            .I(N__5829));
    Sp12to4 I__1323 (
            .O(N__5832),
            .I(N__5824));
    Sp12to4 I__1322 (
            .O(N__5829),
            .I(N__5824));
    Span12Mux_v I__1321 (
            .O(N__5824),
            .I(N__5821));
    Odrv12 I__1320 (
            .O(N__5821),
            .I(A_c_1));
    CascadeMux I__1319 (
            .O(N__5818),
            .I(N__5813));
    InMux I__1318 (
            .O(N__5817),
            .I(N__5805));
    InMux I__1317 (
            .O(N__5816),
            .I(N__5805));
    InMux I__1316 (
            .O(N__5813),
            .I(N__5805));
    InMux I__1315 (
            .O(N__5812),
            .I(N__5802));
    LocalMux I__1314 (
            .O(N__5805),
            .I(N__5797));
    LocalMux I__1313 (
            .O(N__5802),
            .I(N__5797));
    Span4Mux_h I__1312 (
            .O(N__5797),
            .I(N__5794));
    Sp12to4 I__1311 (
            .O(N__5794),
            .I(N__5791));
    Span12Mux_v I__1310 (
            .O(N__5791),
            .I(N__5788));
    Odrv12 I__1309 (
            .O(N__5788),
            .I(A_c_0));
    IoInMux I__1308 (
            .O(N__5785),
            .I(N__5782));
    LocalMux I__1307 (
            .O(N__5782),
            .I(N__5779));
    Odrv4 I__1306 (
            .O(N__5779),
            .I(LMBEn_c));
    InMux I__1305 (
            .O(N__5776),
            .I(N__5773));
    LocalMux I__1304 (
            .O(N__5773),
            .I(N__5770));
    Span4Mux_v I__1303 (
            .O(N__5770),
            .I(N__5767));
    Odrv4 I__1302 (
            .O(N__5767),
            .I(TSn_c));
    InMux I__1301 (
            .O(N__5764),
            .I(N__5761));
    LocalMux I__1300 (
            .O(N__5761),
            .I(N__5758));
    Span4Mux_h I__1299 (
            .O(N__5758),
            .I(N__5755));
    Odrv4 I__1298 (
            .O(N__5755),
            .I(\U400_SDRAM.N_220 ));
    CascadeMux I__1297 (
            .O(N__5752),
            .I(N__5748));
    InMux I__1296 (
            .O(N__5751),
            .I(N__5745));
    InMux I__1295 (
            .O(N__5748),
            .I(N__5738));
    LocalMux I__1294 (
            .O(N__5745),
            .I(N__5735));
    InMux I__1293 (
            .O(N__5744),
            .I(N__5728));
    InMux I__1292 (
            .O(N__5743),
            .I(N__5728));
    InMux I__1291 (
            .O(N__5742),
            .I(N__5728));
    InMux I__1290 (
            .O(N__5741),
            .I(N__5725));
    LocalMux I__1289 (
            .O(N__5738),
            .I(N__5721));
    Span4Mux_v I__1288 (
            .O(N__5735),
            .I(N__5718));
    LocalMux I__1287 (
            .O(N__5728),
            .I(N__5715));
    LocalMux I__1286 (
            .O(N__5725),
            .I(N__5712));
    InMux I__1285 (
            .O(N__5724),
            .I(N__5709));
    Span4Mux_h I__1284 (
            .O(N__5721),
            .I(N__5706));
    Span4Mux_h I__1283 (
            .O(N__5718),
            .I(N__5697));
    Span4Mux_v I__1282 (
            .O(N__5715),
            .I(N__5697));
    Span4Mux_v I__1281 (
            .O(N__5712),
            .I(N__5697));
    LocalMux I__1280 (
            .O(N__5709),
            .I(N__5697));
    Span4Mux_v I__1279 (
            .O(N__5706),
            .I(N__5694));
    IoSpan4Mux I__1278 (
            .O(N__5697),
            .I(N__5691));
    Odrv4 I__1277 (
            .O(N__5694),
            .I(SIZ_c_1));
    Odrv4 I__1276 (
            .O(N__5691),
            .I(SIZ_c_1));
    CascadeMux I__1275 (
            .O(N__5686),
            .I(N__5682));
    InMux I__1274 (
            .O(N__5685),
            .I(N__5676));
    InMux I__1273 (
            .O(N__5682),
            .I(N__5672));
    InMux I__1272 (
            .O(N__5681),
            .I(N__5665));
    InMux I__1271 (
            .O(N__5680),
            .I(N__5665));
    InMux I__1270 (
            .O(N__5679),
            .I(N__5665));
    LocalMux I__1269 (
            .O(N__5676),
            .I(N__5661));
    InMux I__1268 (
            .O(N__5675),
            .I(N__5658));
    LocalMux I__1267 (
            .O(N__5672),
            .I(N__5655));
    LocalMux I__1266 (
            .O(N__5665),
            .I(N__5652));
    InMux I__1265 (
            .O(N__5664),
            .I(N__5649));
    Sp12to4 I__1264 (
            .O(N__5661),
            .I(N__5646));
    LocalMux I__1263 (
            .O(N__5658),
            .I(N__5643));
    Span4Mux_v I__1262 (
            .O(N__5655),
            .I(N__5640));
    Span4Mux_s3_v I__1261 (
            .O(N__5652),
            .I(N__5635));
    LocalMux I__1260 (
            .O(N__5649),
            .I(N__5635));
    Span12Mux_s7_v I__1259 (
            .O(N__5646),
            .I(N__5632));
    Span4Mux_v I__1258 (
            .O(N__5643),
            .I(N__5629));
    Span4Mux_h I__1257 (
            .O(N__5640),
            .I(N__5624));
    Span4Mux_v I__1256 (
            .O(N__5635),
            .I(N__5624));
    Odrv12 I__1255 (
            .O(N__5632),
            .I(SIZ_c_0));
    Odrv4 I__1254 (
            .O(N__5629),
            .I(SIZ_c_0));
    Odrv4 I__1253 (
            .O(N__5624),
            .I(SIZ_c_0));
    InMux I__1252 (
            .O(N__5617),
            .I(N__5614));
    LocalMux I__1251 (
            .O(N__5614),
            .I(N__5610));
    CascadeMux I__1250 (
            .O(N__5613),
            .I(N__5607));
    Span4Mux_v I__1249 (
            .O(N__5610),
            .I(N__5604));
    InMux I__1248 (
            .O(N__5607),
            .I(N__5601));
    Odrv4 I__1247 (
            .O(N__5604),
            .I(\U400_SDRAM.BURST8 ));
    LocalMux I__1246 (
            .O(N__5601),
            .I(\U400_SDRAM.BURST8 ));
    InMux I__1245 (
            .O(N__5596),
            .I(N__5590));
    InMux I__1244 (
            .O(N__5595),
            .I(N__5590));
    LocalMux I__1243 (
            .O(N__5590),
            .I(N__5587));
    Span4Mux_h I__1242 (
            .O(N__5587),
            .I(N__5584));
    Span4Mux_h I__1241 (
            .O(N__5584),
            .I(N__5581));
    Span4Mux_v I__1240 (
            .O(N__5581),
            .I(N__5578));
    Odrv4 I__1239 (
            .O(N__5578),
            .I(A_c_31));
    CascadeMux I__1238 (
            .O(N__5575),
            .I(N__5572));
    InMux I__1237 (
            .O(N__5572),
            .I(N__5566));
    InMux I__1236 (
            .O(N__5571),
            .I(N__5566));
    LocalMux I__1235 (
            .O(N__5566),
            .I(N__5563));
    Span12Mux_v I__1234 (
            .O(N__5563),
            .I(N__5560));
    Odrv12 I__1233 (
            .O(N__5560),
            .I(U400_ADDRESS_DECODE_RAM_SPACE_0_a3_3));
    CascadeMux I__1232 (
            .O(N__5557),
            .I(N__5548));
    InMux I__1231 (
            .O(N__5556),
            .I(N__5545));
    InMux I__1230 (
            .O(N__5555),
            .I(N__5542));
    CascadeMux I__1229 (
            .O(N__5554),
            .I(N__5538));
    CascadeMux I__1228 (
            .O(N__5553),
            .I(N__5535));
    InMux I__1227 (
            .O(N__5552),
            .I(N__5528));
    InMux I__1226 (
            .O(N__5551),
            .I(N__5528));
    InMux I__1225 (
            .O(N__5548),
            .I(N__5528));
    LocalMux I__1224 (
            .O(N__5545),
            .I(N__5519));
    LocalMux I__1223 (
            .O(N__5542),
            .I(N__5516));
    InMux I__1222 (
            .O(N__5541),
            .I(N__5513));
    InMux I__1221 (
            .O(N__5538),
            .I(N__5510));
    InMux I__1220 (
            .O(N__5535),
            .I(N__5507));
    LocalMux I__1219 (
            .O(N__5528),
            .I(N__5504));
    InMux I__1218 (
            .O(N__5527),
            .I(N__5499));
    InMux I__1217 (
            .O(N__5526),
            .I(N__5499));
    InMux I__1216 (
            .O(N__5525),
            .I(N__5494));
    InMux I__1215 (
            .O(N__5524),
            .I(N__5494));
    InMux I__1214 (
            .O(N__5523),
            .I(N__5491));
    InMux I__1213 (
            .O(N__5522),
            .I(N__5485));
    Span4Mux_v I__1212 (
            .O(N__5519),
            .I(N__5482));
    Span4Mux_v I__1211 (
            .O(N__5516),
            .I(N__5479));
    LocalMux I__1210 (
            .O(N__5513),
            .I(N__5474));
    LocalMux I__1209 (
            .O(N__5510),
            .I(N__5474));
    LocalMux I__1208 (
            .O(N__5507),
            .I(N__5471));
    Span4Mux_h I__1207 (
            .O(N__5504),
            .I(N__5464));
    LocalMux I__1206 (
            .O(N__5499),
            .I(N__5464));
    LocalMux I__1205 (
            .O(N__5494),
            .I(N__5464));
    LocalMux I__1204 (
            .O(N__5491),
            .I(N__5461));
    InMux I__1203 (
            .O(N__5490),
            .I(N__5456));
    InMux I__1202 (
            .O(N__5489),
            .I(N__5456));
    InMux I__1201 (
            .O(N__5488),
            .I(N__5453));
    LocalMux I__1200 (
            .O(N__5485),
            .I(N__5450));
    Span4Mux_v I__1199 (
            .O(N__5482),
            .I(N__5443));
    Span4Mux_h I__1198 (
            .O(N__5479),
            .I(N__5443));
    Span4Mux_v I__1197 (
            .O(N__5474),
            .I(N__5443));
    Span4Mux_v I__1196 (
            .O(N__5471),
            .I(N__5440));
    Span4Mux_v I__1195 (
            .O(N__5464),
            .I(N__5437));
    Span4Mux_h I__1194 (
            .O(N__5461),
            .I(N__5432));
    LocalMux I__1193 (
            .O(N__5456),
            .I(N__5432));
    LocalMux I__1192 (
            .O(N__5453),
            .I(N__5429));
    Span12Mux_s8_v I__1191 (
            .O(N__5450),
            .I(N__5426));
    Span4Mux_h I__1190 (
            .O(N__5443),
            .I(N__5423));
    Span4Mux_h I__1189 (
            .O(N__5440),
            .I(N__5418));
    Span4Mux_h I__1188 (
            .O(N__5437),
            .I(N__5418));
    Span4Mux_v I__1187 (
            .O(N__5432),
            .I(N__5413));
    Span4Mux_v I__1186 (
            .O(N__5429),
            .I(N__5413));
    Odrv12 I__1185 (
            .O(N__5426),
            .I(RESETn_c));
    Odrv4 I__1184 (
            .O(N__5423),
            .I(RESETn_c));
    Odrv4 I__1183 (
            .O(N__5418),
            .I(RESETn_c));
    Odrv4 I__1182 (
            .O(N__5413),
            .I(RESETn_c));
    IoInMux I__1181 (
            .O(N__5404),
            .I(N__5401));
    LocalMux I__1180 (
            .O(N__5401),
            .I(N__5398));
    Odrv12 I__1179 (
            .O(N__5398),
            .I(N_220_3_i));
    InMux I__1178 (
            .O(N__5395),
            .I(N__5392));
    LocalMux I__1177 (
            .O(N__5392),
            .I(N__5389));
    Odrv4 I__1176 (
            .O(N__5389),
            .I(A_c_5));
    CascadeMux I__1175 (
            .O(N__5386),
            .I(N__5383));
    InMux I__1174 (
            .O(N__5383),
            .I(N__5380));
    LocalMux I__1173 (
            .O(N__5380),
            .I(N__5377));
    Span4Mux_v I__1172 (
            .O(N__5377),
            .I(N__5374));
    Odrv4 I__1171 (
            .O(N__5374),
            .I(A_c_13));
    IoInMux I__1170 (
            .O(N__5371),
            .I(N__5368));
    LocalMux I__1169 (
            .O(N__5368),
            .I(N__5365));
    Span12Mux_s3_v I__1168 (
            .O(N__5365),
            .I(N__5362));
    Odrv12 I__1167 (
            .O(N__5362),
            .I(MA_c_3));
    InMux I__1166 (
            .O(N__5359),
            .I(N__5356));
    LocalMux I__1165 (
            .O(N__5356),
            .I(N__5353));
    Span4Mux_h I__1164 (
            .O(N__5353),
            .I(N__5350));
    Odrv4 I__1163 (
            .O(N__5350),
            .I(A_c_3));
    CascadeMux I__1162 (
            .O(N__5347),
            .I(N__5344));
    InMux I__1161 (
            .O(N__5344),
            .I(N__5341));
    LocalMux I__1160 (
            .O(N__5341),
            .I(N__5338));
    Odrv4 I__1159 (
            .O(N__5338),
            .I(A_c_11));
    CascadeMux I__1158 (
            .O(N__5335),
            .I(N__5331));
    InMux I__1157 (
            .O(N__5334),
            .I(N__5328));
    InMux I__1156 (
            .O(N__5331),
            .I(N__5325));
    LocalMux I__1155 (
            .O(N__5328),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__1154 (
            .O(N__5325),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_7 ));
    CEMux I__1153 (
            .O(N__5320),
            .I(N__5316));
    CEMux I__1152 (
            .O(N__5319),
            .I(N__5311));
    LocalMux I__1151 (
            .O(N__5316),
            .I(N__5308));
    CEMux I__1150 (
            .O(N__5315),
            .I(N__5305));
    CEMux I__1149 (
            .O(N__5314),
            .I(N__5302));
    LocalMux I__1148 (
            .O(N__5311),
            .I(N__5299));
    Span4Mux_v I__1147 (
            .O(N__5308),
            .I(N__5294));
    LocalMux I__1146 (
            .O(N__5305),
            .I(N__5294));
    LocalMux I__1145 (
            .O(N__5302),
            .I(N__5291));
    Span4Mux_v I__1144 (
            .O(N__5299),
            .I(N__5286));
    Span4Mux_h I__1143 (
            .O(N__5294),
            .I(N__5286));
    Odrv12 I__1142 (
            .O(N__5291),
            .I(\U400_SDRAM.SDRAM_COUNTERe_0_i ));
    Odrv4 I__1141 (
            .O(N__5286),
            .I(\U400_SDRAM.SDRAM_COUNTERe_0_i ));
    CascadeMux I__1140 (
            .O(N__5281),
            .I(N__5277));
    InMux I__1139 (
            .O(N__5280),
            .I(N__5263));
    InMux I__1138 (
            .O(N__5277),
            .I(N__5260));
    InMux I__1137 (
            .O(N__5276),
            .I(N__5257));
    InMux I__1136 (
            .O(N__5275),
            .I(N__5252));
    InMux I__1135 (
            .O(N__5274),
            .I(N__5252));
    InMux I__1134 (
            .O(N__5273),
            .I(N__5243));
    InMux I__1133 (
            .O(N__5272),
            .I(N__5243));
    InMux I__1132 (
            .O(N__5271),
            .I(N__5243));
    InMux I__1131 (
            .O(N__5270),
            .I(N__5243));
    InMux I__1130 (
            .O(N__5269),
            .I(N__5237));
    InMux I__1129 (
            .O(N__5268),
            .I(N__5233));
    InMux I__1128 (
            .O(N__5267),
            .I(N__5229));
    InMux I__1127 (
            .O(N__5266),
            .I(N__5226));
    LocalMux I__1126 (
            .O(N__5263),
            .I(N__5220));
    LocalMux I__1125 (
            .O(N__5260),
            .I(N__5220));
    LocalMux I__1124 (
            .O(N__5257),
            .I(N__5213));
    LocalMux I__1123 (
            .O(N__5252),
            .I(N__5213));
    LocalMux I__1122 (
            .O(N__5243),
            .I(N__5213));
    InMux I__1121 (
            .O(N__5242),
            .I(N__5210));
    InMux I__1120 (
            .O(N__5241),
            .I(N__5205));
    InMux I__1119 (
            .O(N__5240),
            .I(N__5205));
    LocalMux I__1118 (
            .O(N__5237),
            .I(N__5202));
    InMux I__1117 (
            .O(N__5236),
            .I(N__5199));
    LocalMux I__1116 (
            .O(N__5233),
            .I(N__5196));
    InMux I__1115 (
            .O(N__5232),
            .I(N__5193));
    LocalMux I__1114 (
            .O(N__5229),
            .I(N__5188));
    LocalMux I__1113 (
            .O(N__5226),
            .I(N__5188));
    InMux I__1112 (
            .O(N__5225),
            .I(N__5185));
    Span4Mux_v I__1111 (
            .O(N__5220),
            .I(N__5178));
    Span4Mux_v I__1110 (
            .O(N__5213),
            .I(N__5178));
    LocalMux I__1109 (
            .O(N__5210),
            .I(N__5178));
    LocalMux I__1108 (
            .O(N__5205),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv12 I__1107 (
            .O(N__5202),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1106 (
            .O(N__5199),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1105 (
            .O(N__5196),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1104 (
            .O(N__5193),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv12 I__1103 (
            .O(N__5188),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1102 (
            .O(N__5185),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1101 (
            .O(N__5178),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    CascadeMux I__1100 (
            .O(N__5161),
            .I(N__5156));
    CascadeMux I__1099 (
            .O(N__5160),
            .I(N__5153));
    CascadeMux I__1098 (
            .O(N__5159),
            .I(N__5146));
    InMux I__1097 (
            .O(N__5156),
            .I(N__5143));
    InMux I__1096 (
            .O(N__5153),
            .I(N__5139));
    CascadeMux I__1095 (
            .O(N__5152),
            .I(N__5136));
    CascadeMux I__1094 (
            .O(N__5151),
            .I(N__5132));
    CascadeMux I__1093 (
            .O(N__5150),
            .I(N__5128));
    InMux I__1092 (
            .O(N__5149),
            .I(N__5122));
    InMux I__1091 (
            .O(N__5146),
            .I(N__5122));
    LocalMux I__1090 (
            .O(N__5143),
            .I(N__5119));
    InMux I__1089 (
            .O(N__5142),
            .I(N__5116));
    LocalMux I__1088 (
            .O(N__5139),
            .I(N__5113));
    InMux I__1087 (
            .O(N__5136),
            .I(N__5110));
    InMux I__1086 (
            .O(N__5135),
            .I(N__5103));
    InMux I__1085 (
            .O(N__5132),
            .I(N__5103));
    InMux I__1084 (
            .O(N__5131),
            .I(N__5103));
    InMux I__1083 (
            .O(N__5128),
            .I(N__5098));
    InMux I__1082 (
            .O(N__5127),
            .I(N__5098));
    LocalMux I__1081 (
            .O(N__5122),
            .I(N__5093));
    Span4Mux_v I__1080 (
            .O(N__5119),
            .I(N__5093));
    LocalMux I__1079 (
            .O(N__5116),
            .I(\U400_SDRAM.WRITE_CYCLEZ0 ));
    Odrv4 I__1078 (
            .O(N__5113),
            .I(\U400_SDRAM.WRITE_CYCLEZ0 ));
    LocalMux I__1077 (
            .O(N__5110),
            .I(\U400_SDRAM.WRITE_CYCLEZ0 ));
    LocalMux I__1076 (
            .O(N__5103),
            .I(\U400_SDRAM.WRITE_CYCLEZ0 ));
    LocalMux I__1075 (
            .O(N__5098),
            .I(\U400_SDRAM.WRITE_CYCLEZ0 ));
    Odrv4 I__1074 (
            .O(N__5093),
            .I(\U400_SDRAM.WRITE_CYCLEZ0 ));
    InMux I__1073 (
            .O(N__5080),
            .I(N__5065));
    InMux I__1072 (
            .O(N__5079),
            .I(N__5065));
    InMux I__1071 (
            .O(N__5078),
            .I(N__5065));
    InMux I__1070 (
            .O(N__5077),
            .I(N__5062));
    InMux I__1069 (
            .O(N__5076),
            .I(N__5059));
    CascadeMux I__1068 (
            .O(N__5075),
            .I(N__5056));
    CascadeMux I__1067 (
            .O(N__5074),
            .I(N__5053));
    InMux I__1066 (
            .O(N__5073),
            .I(N__5050));
    InMux I__1065 (
            .O(N__5072),
            .I(N__5047));
    LocalMux I__1064 (
            .O(N__5065),
            .I(N__5044));
    LocalMux I__1063 (
            .O(N__5062),
            .I(N__5033));
    LocalMux I__1062 (
            .O(N__5059),
            .I(N__5033));
    InMux I__1061 (
            .O(N__5056),
            .I(N__5028));
    InMux I__1060 (
            .O(N__5053),
            .I(N__5028));
    LocalMux I__1059 (
            .O(N__5050),
            .I(N__5023));
    LocalMux I__1058 (
            .O(N__5047),
            .I(N__5023));
    Span4Mux_h I__1057 (
            .O(N__5044),
            .I(N__5018));
    InMux I__1056 (
            .O(N__5043),
            .I(N__5013));
    InMux I__1055 (
            .O(N__5042),
            .I(N__5013));
    InMux I__1054 (
            .O(N__5041),
            .I(N__5010));
    InMux I__1053 (
            .O(N__5040),
            .I(N__5007));
    InMux I__1052 (
            .O(N__5039),
            .I(N__5004));
    InMux I__1051 (
            .O(N__5038),
            .I(N__5001));
    Span4Mux_h I__1050 (
            .O(N__5033),
            .I(N__4994));
    LocalMux I__1049 (
            .O(N__5028),
            .I(N__4994));
    Span4Mux_h I__1048 (
            .O(N__5023),
            .I(N__4994));
    InMux I__1047 (
            .O(N__5022),
            .I(N__4989));
    InMux I__1046 (
            .O(N__5021),
            .I(N__4989));
    Odrv4 I__1045 (
            .O(N__5018),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1044 (
            .O(N__5013),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1043 (
            .O(N__5010),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1042 (
            .O(N__5007),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1041 (
            .O(N__5004),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1040 (
            .O(N__5001),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1039 (
            .O(N__4994),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1038 (
            .O(N__4989),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    CascadeMux I__1037 (
            .O(N__4972),
            .I(\U400_SDRAM.N_161_cascade_ ));
    InMux I__1036 (
            .O(N__4969),
            .I(N__4966));
    LocalMux I__1035 (
            .O(N__4966),
            .I(\U400_SDRAM.N_183 ));
    InMux I__1034 (
            .O(N__4963),
            .I(N__4952));
    InMux I__1033 (
            .O(N__4962),
            .I(N__4952));
    InMux I__1032 (
            .O(N__4961),
            .I(N__4952));
    InMux I__1031 (
            .O(N__4960),
            .I(N__4941));
    InMux I__1030 (
            .O(N__4959),
            .I(N__4941));
    LocalMux I__1029 (
            .O(N__4952),
            .I(N__4935));
    InMux I__1028 (
            .O(N__4951),
            .I(N__4930));
    InMux I__1027 (
            .O(N__4950),
            .I(N__4930));
    InMux I__1026 (
            .O(N__4949),
            .I(N__4923));
    InMux I__1025 (
            .O(N__4948),
            .I(N__4920));
    InMux I__1024 (
            .O(N__4947),
            .I(N__4917));
    InMux I__1023 (
            .O(N__4946),
            .I(N__4914));
    LocalMux I__1022 (
            .O(N__4941),
            .I(N__4911));
    InMux I__1021 (
            .O(N__4940),
            .I(N__4908));
    InMux I__1020 (
            .O(N__4939),
            .I(N__4903));
    InMux I__1019 (
            .O(N__4938),
            .I(N__4903));
    Span4Mux_h I__1018 (
            .O(N__4935),
            .I(N__4898));
    LocalMux I__1017 (
            .O(N__4930),
            .I(N__4898));
    InMux I__1016 (
            .O(N__4929),
            .I(N__4895));
    InMux I__1015 (
            .O(N__4928),
            .I(N__4888));
    InMux I__1014 (
            .O(N__4927),
            .I(N__4888));
    InMux I__1013 (
            .O(N__4926),
            .I(N__4888));
    LocalMux I__1012 (
            .O(N__4923),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1011 (
            .O(N__4920),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1010 (
            .O(N__4917),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1009 (
            .O(N__4914),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv12 I__1008 (
            .O(N__4911),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1007 (
            .O(N__4908),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1006 (
            .O(N__4903),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1005 (
            .O(N__4898),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1004 (
            .O(N__4895),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1003 (
            .O(N__4888),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__1002 (
            .O(N__4867),
            .I(N__4863));
    InMux I__1001 (
            .O(N__4866),
            .I(N__4859));
    LocalMux I__1000 (
            .O(N__4863),
            .I(N__4856));
    InMux I__999 (
            .O(N__4862),
            .I(N__4851));
    LocalMux I__998 (
            .O(N__4859),
            .I(N__4848));
    Span4Mux_h I__997 (
            .O(N__4856),
            .I(N__4845));
    InMux I__996 (
            .O(N__4855),
            .I(N__4842));
    InMux I__995 (
            .O(N__4854),
            .I(N__4839));
    LocalMux I__994 (
            .O(N__4851),
            .I(\U400_SDRAM.N_126 ));
    Odrv4 I__993 (
            .O(N__4848),
            .I(\U400_SDRAM.N_126 ));
    Odrv4 I__992 (
            .O(N__4845),
            .I(\U400_SDRAM.N_126 ));
    LocalMux I__991 (
            .O(N__4842),
            .I(\U400_SDRAM.N_126 ));
    LocalMux I__990 (
            .O(N__4839),
            .I(\U400_SDRAM.N_126 ));
    CascadeMux I__989 (
            .O(N__4828),
            .I(N__4821));
    InMux I__988 (
            .O(N__4827),
            .I(N__4818));
    InMux I__987 (
            .O(N__4826),
            .I(N__4815));
    InMux I__986 (
            .O(N__4825),
            .I(N__4812));
    InMux I__985 (
            .O(N__4824),
            .I(N__4809));
    InMux I__984 (
            .O(N__4821),
            .I(N__4806));
    LocalMux I__983 (
            .O(N__4818),
            .I(N__4799));
    LocalMux I__982 (
            .O(N__4815),
            .I(N__4796));
    LocalMux I__981 (
            .O(N__4812),
            .I(N__4789));
    LocalMux I__980 (
            .O(N__4809),
            .I(N__4789));
    LocalMux I__979 (
            .O(N__4806),
            .I(N__4789));
    InMux I__978 (
            .O(N__4805),
            .I(N__4786));
    InMux I__977 (
            .O(N__4804),
            .I(N__4781));
    InMux I__976 (
            .O(N__4803),
            .I(N__4781));
    InMux I__975 (
            .O(N__4802),
            .I(N__4775));
    Span4Mux_h I__974 (
            .O(N__4799),
            .I(N__4772));
    Span4Mux_v I__973 (
            .O(N__4796),
            .I(N__4767));
    Span4Mux_v I__972 (
            .O(N__4789),
            .I(N__4767));
    LocalMux I__971 (
            .O(N__4786),
            .I(N__4762));
    LocalMux I__970 (
            .O(N__4781),
            .I(N__4762));
    InMux I__969 (
            .O(N__4780),
            .I(N__4757));
    InMux I__968 (
            .O(N__4779),
            .I(N__4757));
    InMux I__967 (
            .O(N__4778),
            .I(N__4754));
    LocalMux I__966 (
            .O(N__4775),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__965 (
            .O(N__4772),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__964 (
            .O(N__4767),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__963 (
            .O(N__4762),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__962 (
            .O(N__4757),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__961 (
            .O(N__4754),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__960 (
            .O(N__4741),
            .I(N__4738));
    LocalMux I__959 (
            .O(N__4738),
            .I(N__4735));
    Span4Mux_v I__958 (
            .O(N__4735),
            .I(N__4731));
    InMux I__957 (
            .O(N__4734),
            .I(N__4728));
    Odrv4 I__956 (
            .O(N__4731),
            .I(\U400_SDRAM.N_138 ));
    LocalMux I__955 (
            .O(N__4728),
            .I(\U400_SDRAM.N_138 ));
    CascadeMux I__954 (
            .O(N__4723),
            .I(N__4720));
    InMux I__953 (
            .O(N__4720),
            .I(N__4717));
    LocalMux I__952 (
            .O(N__4717),
            .I(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_a3_1_0_0 ));
    CascadeMux I__951 (
            .O(N__4714),
            .I(N__4703));
    CascadeMux I__950 (
            .O(N__4713),
            .I(N__4700));
    InMux I__949 (
            .O(N__4712),
            .I(N__4697));
    CascadeMux I__948 (
            .O(N__4711),
            .I(N__4694));
    CascadeMux I__947 (
            .O(N__4710),
            .I(N__4691));
    CascadeMux I__946 (
            .O(N__4709),
            .I(N__4688));
    CascadeMux I__945 (
            .O(N__4708),
            .I(N__4685));
    CascadeMux I__944 (
            .O(N__4707),
            .I(N__4681));
    CascadeMux I__943 (
            .O(N__4706),
            .I(N__4677));
    InMux I__942 (
            .O(N__4703),
            .I(N__4674));
    InMux I__941 (
            .O(N__4700),
            .I(N__4671));
    LocalMux I__940 (
            .O(N__4697),
            .I(N__4668));
    InMux I__939 (
            .O(N__4694),
            .I(N__4661));
    InMux I__938 (
            .O(N__4691),
            .I(N__4661));
    InMux I__937 (
            .O(N__4688),
            .I(N__4661));
    InMux I__936 (
            .O(N__4685),
            .I(N__4654));
    InMux I__935 (
            .O(N__4684),
            .I(N__4654));
    InMux I__934 (
            .O(N__4681),
            .I(N__4647));
    InMux I__933 (
            .O(N__4680),
            .I(N__4647));
    InMux I__932 (
            .O(N__4677),
            .I(N__4647));
    LocalMux I__931 (
            .O(N__4674),
            .I(N__4642));
    LocalMux I__930 (
            .O(N__4671),
            .I(N__4642));
    Span4Mux_v I__929 (
            .O(N__4668),
            .I(N__4635));
    LocalMux I__928 (
            .O(N__4661),
            .I(N__4635));
    InMux I__927 (
            .O(N__4660),
            .I(N__4630));
    InMux I__926 (
            .O(N__4659),
            .I(N__4630));
    LocalMux I__925 (
            .O(N__4654),
            .I(N__4622));
    LocalMux I__924 (
            .O(N__4647),
            .I(N__4622));
    Span4Mux_h I__923 (
            .O(N__4642),
            .I(N__4619));
    InMux I__922 (
            .O(N__4641),
            .I(N__4616));
    InMux I__921 (
            .O(N__4640),
            .I(N__4613));
    Span4Mux_h I__920 (
            .O(N__4635),
            .I(N__4608));
    LocalMux I__919 (
            .O(N__4630),
            .I(N__4608));
    InMux I__918 (
            .O(N__4629),
            .I(N__4603));
    InMux I__917 (
            .O(N__4628),
            .I(N__4603));
    InMux I__916 (
            .O(N__4627),
            .I(N__4600));
    Span4Mux_v I__915 (
            .O(N__4622),
            .I(N__4597));
    Odrv4 I__914 (
            .O(N__4619),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__913 (
            .O(N__4616),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__912 (
            .O(N__4613),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__911 (
            .O(N__4608),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__910 (
            .O(N__4603),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__909 (
            .O(N__4600),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__908 (
            .O(N__4597),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    CascadeMux I__907 (
            .O(N__4582),
            .I(N__4578));
    InMux I__906 (
            .O(N__4581),
            .I(N__4573));
    InMux I__905 (
            .O(N__4578),
            .I(N__4570));
    InMux I__904 (
            .O(N__4577),
            .I(N__4567));
    CascadeMux I__903 (
            .O(N__4576),
            .I(N__4562));
    LocalMux I__902 (
            .O(N__4573),
            .I(N__4559));
    LocalMux I__901 (
            .O(N__4570),
            .I(N__4556));
    LocalMux I__900 (
            .O(N__4567),
            .I(N__4553));
    InMux I__899 (
            .O(N__4566),
            .I(N__4548));
    InMux I__898 (
            .O(N__4565),
            .I(N__4548));
    InMux I__897 (
            .O(N__4562),
            .I(N__4545));
    Span4Mux_h I__896 (
            .O(N__4559),
            .I(N__4542));
    Span4Mux_h I__895 (
            .O(N__4556),
            .I(N__4533));
    Span4Mux_h I__894 (
            .O(N__4553),
            .I(N__4533));
    LocalMux I__893 (
            .O(N__4548),
            .I(N__4533));
    LocalMux I__892 (
            .O(N__4545),
            .I(N__4533));
    Odrv4 I__891 (
            .O(N__4542),
            .I(\U400_SDRAM.SDRAM_CONFIGURED_RNIVK7JZ0 ));
    Odrv4 I__890 (
            .O(N__4533),
            .I(\U400_SDRAM.SDRAM_CONFIGURED_RNIVK7JZ0 ));
    InMux I__889 (
            .O(N__4528),
            .I(N__4525));
    LocalMux I__888 (
            .O(N__4525),
            .I(N__4522));
    Span4Mux_s2_v I__887 (
            .O(N__4522),
            .I(N__4519));
    Odrv4 I__886 (
            .O(N__4519),
            .I(A_c_7));
    CascadeMux I__885 (
            .O(N__4516),
            .I(N__4513));
    InMux I__884 (
            .O(N__4513),
            .I(N__4510));
    LocalMux I__883 (
            .O(N__4510),
            .I(N__4507));
    IoSpan4Mux I__882 (
            .O(N__4507),
            .I(N__4504));
    Odrv4 I__881 (
            .O(N__4504),
            .I(A_c_15));
    InMux I__880 (
            .O(N__4501),
            .I(N__4498));
    LocalMux I__879 (
            .O(N__4498),
            .I(\U400_SDRAM.MAc_0_0 ));
    InMux I__878 (
            .O(N__4495),
            .I(N__4492));
    LocalMux I__877 (
            .O(N__4492),
            .I(N__4489));
    Span4Mux_h I__876 (
            .O(N__4489),
            .I(N__4486));
    Odrv4 I__875 (
            .O(N__4486),
            .I(A_c_2));
    CascadeMux I__874 (
            .O(N__4483),
            .I(N__4480));
    InMux I__873 (
            .O(N__4480),
            .I(N__4477));
    LocalMux I__872 (
            .O(N__4477),
            .I(N__4474));
    Span4Mux_s1_v I__871 (
            .O(N__4474),
            .I(N__4471));
    Odrv4 I__870 (
            .O(N__4471),
            .I(A_c_10));
    IoInMux I__869 (
            .O(N__4468),
            .I(N__4465));
    LocalMux I__868 (
            .O(N__4465),
            .I(MA_c_0));
    InMux I__867 (
            .O(N__4462),
            .I(N__4459));
    LocalMux I__866 (
            .O(N__4459),
            .I(N__4456));
    Span12Mux_s10_h I__865 (
            .O(N__4456),
            .I(N__4453));
    Span12Mux_v I__864 (
            .O(N__4453),
            .I(N__4450));
    Odrv12 I__863 (
            .O(N__4450),
            .I(A_c_20));
    InMux I__862 (
            .O(N__4447),
            .I(N__4444));
    LocalMux I__861 (
            .O(N__4444),
            .I(\U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5Z0Z_0 ));
    InMux I__860 (
            .O(N__4441),
            .I(N__4438));
    LocalMux I__859 (
            .O(N__4438),
            .I(N__4435));
    Span4Mux_h I__858 (
            .O(N__4435),
            .I(N__4428));
    InMux I__857 (
            .O(N__4434),
            .I(N__4425));
    InMux I__856 (
            .O(N__4433),
            .I(N__4422));
    InMux I__855 (
            .O(N__4432),
            .I(N__4419));
    InMux I__854 (
            .O(N__4431),
            .I(N__4416));
    Odrv4 I__853 (
            .O(N__4428),
            .I(\U400_SDRAM.N_129 ));
    LocalMux I__852 (
            .O(N__4425),
            .I(\U400_SDRAM.N_129 ));
    LocalMux I__851 (
            .O(N__4422),
            .I(\U400_SDRAM.N_129 ));
    LocalMux I__850 (
            .O(N__4419),
            .I(\U400_SDRAM.N_129 ));
    LocalMux I__849 (
            .O(N__4416),
            .I(\U400_SDRAM.N_129 ));
    InMux I__848 (
            .O(N__4405),
            .I(N__4401));
    InMux I__847 (
            .O(N__4404),
            .I(N__4397));
    LocalMux I__846 (
            .O(N__4401),
            .I(N__4394));
    InMux I__845 (
            .O(N__4400),
            .I(N__4391));
    LocalMux I__844 (
            .O(N__4397),
            .I(\U400_SDRAM.N_260 ));
    Odrv4 I__843 (
            .O(N__4394),
            .I(\U400_SDRAM.N_260 ));
    LocalMux I__842 (
            .O(N__4391),
            .I(\U400_SDRAM.N_260 ));
    InMux I__841 (
            .O(N__4384),
            .I(N__4381));
    LocalMux I__840 (
            .O(N__4381),
            .I(\U400_SDRAM.SDRAM_COUNTER_s_1 ));
    InMux I__839 (
            .O(N__4378),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_0 ));
    InMux I__838 (
            .O(N__4375),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_1 ));
    InMux I__837 (
            .O(N__4372),
            .I(N__4369));
    LocalMux I__836 (
            .O(N__4369),
            .I(\U400_SDRAM.SDRAM_COUNTER_s_3 ));
    InMux I__835 (
            .O(N__4366),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_2 ));
    InMux I__834 (
            .O(N__4363),
            .I(N__4359));
    InMux I__833 (
            .O(N__4362),
            .I(N__4356));
    LocalMux I__832 (
            .O(N__4359),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__831 (
            .O(N__4356),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__830 (
            .O(N__4351),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_3 ));
    InMux I__829 (
            .O(N__4348),
            .I(N__4344));
    InMux I__828 (
            .O(N__4347),
            .I(N__4341));
    LocalMux I__827 (
            .O(N__4344),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__826 (
            .O(N__4341),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_5 ));
    InMux I__825 (
            .O(N__4336),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_4 ));
    InMux I__824 (
            .O(N__4333),
            .I(N__4329));
    InMux I__823 (
            .O(N__4332),
            .I(N__4326));
    LocalMux I__822 (
            .O(N__4329),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__821 (
            .O(N__4326),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__820 (
            .O(N__4321),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_5 ));
    InMux I__819 (
            .O(N__4318),
            .I(N__4307));
    InMux I__818 (
            .O(N__4317),
            .I(N__4307));
    InMux I__817 (
            .O(N__4316),
            .I(N__4307));
    InMux I__816 (
            .O(N__4315),
            .I(N__4301));
    InMux I__815 (
            .O(N__4314),
            .I(N__4298));
    LocalMux I__814 (
            .O(N__4307),
            .I(N__4295));
    InMux I__813 (
            .O(N__4306),
            .I(N__4292));
    InMux I__812 (
            .O(N__4305),
            .I(N__4287));
    InMux I__811 (
            .O(N__4304),
            .I(N__4287));
    LocalMux I__810 (
            .O(N__4301),
            .I(\U400_SDRAM.N_37 ));
    LocalMux I__809 (
            .O(N__4298),
            .I(\U400_SDRAM.N_37 ));
    Odrv4 I__808 (
            .O(N__4295),
            .I(\U400_SDRAM.N_37 ));
    LocalMux I__807 (
            .O(N__4292),
            .I(\U400_SDRAM.N_37 ));
    LocalMux I__806 (
            .O(N__4287),
            .I(\U400_SDRAM.N_37 ));
    InMux I__805 (
            .O(N__4276),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_6 ));
    CascadeMux I__804 (
            .O(N__4273),
            .I(N__4270));
    InMux I__803 (
            .O(N__4270),
            .I(N__4267));
    LocalMux I__802 (
            .O(N__4267),
            .I(N__4264));
    Span12Mux_v I__801 (
            .O(N__4264),
            .I(N__4261));
    Odrv12 I__800 (
            .O(N__4261),
            .I(A_c_25));
    IoInMux I__799 (
            .O(N__4258),
            .I(N__4255));
    LocalMux I__798 (
            .O(N__4255),
            .I(N__4252));
    Span4Mux_s3_v I__797 (
            .O(N__4252),
            .I(N__4249));
    Odrv4 I__796 (
            .O(N__4249),
            .I(MA_c_11));
    InMux I__795 (
            .O(N__4246),
            .I(N__4243));
    LocalMux I__794 (
            .O(N__4243),
            .I(N__4236));
    InMux I__793 (
            .O(N__4242),
            .I(N__4233));
    InMux I__792 (
            .O(N__4241),
            .I(N__4230));
    InMux I__791 (
            .O(N__4240),
            .I(N__4225));
    InMux I__790 (
            .O(N__4239),
            .I(N__4225));
    Odrv4 I__789 (
            .O(N__4236),
            .I(\U400_SDRAM.N_257 ));
    LocalMux I__788 (
            .O(N__4233),
            .I(\U400_SDRAM.N_257 ));
    LocalMux I__787 (
            .O(N__4230),
            .I(\U400_SDRAM.N_257 ));
    LocalMux I__786 (
            .O(N__4225),
            .I(\U400_SDRAM.N_257 ));
    InMux I__785 (
            .O(N__4216),
            .I(N__4213));
    LocalMux I__784 (
            .O(N__4213),
            .I(N__4210));
    Span4Mux_s3_v I__783 (
            .O(N__4210),
            .I(N__4207));
    Span4Mux_h I__782 (
            .O(N__4207),
            .I(N__4204));
    Odrv4 I__781 (
            .O(N__4204),
            .I(A_c_6));
    CascadeMux I__780 (
            .O(N__4201),
            .I(N__4198));
    InMux I__779 (
            .O(N__4198),
            .I(N__4195));
    LocalMux I__778 (
            .O(N__4195),
            .I(N__4192));
    Span4Mux_h I__777 (
            .O(N__4192),
            .I(N__4189));
    Odrv4 I__776 (
            .O(N__4189),
            .I(A_c_14));
    IoInMux I__775 (
            .O(N__4186),
            .I(N__4183));
    LocalMux I__774 (
            .O(N__4183),
            .I(N__4180));
    Span4Mux_s0_v I__773 (
            .O(N__4180),
            .I(N__4177));
    Span4Mux_h I__772 (
            .O(N__4177),
            .I(N__4174));
    Odrv4 I__771 (
            .O(N__4174),
            .I(MA_c_4));
    IoInMux I__770 (
            .O(N__4171),
            .I(N__4168));
    LocalMux I__769 (
            .O(N__4168),
            .I(N__4165));
    IoSpan4Mux I__768 (
            .O(N__4165),
            .I(N__4162));
    Odrv4 I__767 (
            .O(N__4162),
            .I(MA_c_5));
    InMux I__766 (
            .O(N__4159),
            .I(N__4156));
    LocalMux I__765 (
            .O(N__4156),
            .I(N__4153));
    Odrv4 I__764 (
            .O(N__4153),
            .I(\U400_SDRAM.N_150 ));
    CascadeMux I__763 (
            .O(N__4150),
            .I(\U400_SDRAM.N_150_cascade_ ));
    InMux I__762 (
            .O(N__4147),
            .I(N__4143));
    InMux I__761 (
            .O(N__4146),
            .I(N__4140));
    LocalMux I__760 (
            .O(N__4143),
            .I(\U400_SDRAM.N_252 ));
    LocalMux I__759 (
            .O(N__4140),
            .I(\U400_SDRAM.N_252 ));
    CascadeMux I__758 (
            .O(N__4135),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_61_i_i_a3_1_0_cascade_ ));
    InMux I__757 (
            .O(N__4132),
            .I(N__4126));
    InMux I__756 (
            .O(N__4131),
            .I(N__4126));
    LocalMux I__755 (
            .O(N__4126),
            .I(\U400_SDRAM.N_201 ));
    InMux I__754 (
            .O(N__4123),
            .I(N__4120));
    LocalMux I__753 (
            .O(N__4120),
            .I(TA_EN_i_ess));
    IoInMux I__752 (
            .O(N__4117),
            .I(N__4114));
    LocalMux I__751 (
            .O(N__4114),
            .I(N__4111));
    Odrv12 I__750 (
            .O(N__4111),
            .I(N_529_i));
    CascadeMux I__749 (
            .O(N__4108),
            .I(\U400_SDRAM.N_126_cascade_ ));
    CascadeMux I__748 (
            .O(N__4105),
            .I(\U400_SDRAM.N_129_cascade_ ));
    CascadeMux I__747 (
            .O(N__4102),
            .I(\U400_SDRAM.N_257_cascade_ ));
    InMux I__746 (
            .O(N__4099),
            .I(N__4096));
    LocalMux I__745 (
            .O(N__4096),
            .I(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_1_0 ));
    InMux I__744 (
            .O(N__4093),
            .I(N__4088));
    InMux I__743 (
            .O(N__4092),
            .I(N__4083));
    InMux I__742 (
            .O(N__4091),
            .I(N__4083));
    LocalMux I__741 (
            .O(N__4088),
            .I(\U400_SDRAM.N_133 ));
    LocalMux I__740 (
            .O(N__4083),
            .I(\U400_SDRAM.N_133 ));
    CascadeMux I__739 (
            .O(N__4078),
            .I(\U400_SDRAM.N_133_cascade_ ));
    CascadeMux I__738 (
            .O(N__4075),
            .I(N__4070));
    InMux I__737 (
            .O(N__4074),
            .I(N__4060));
    InMux I__736 (
            .O(N__4073),
            .I(N__4060));
    InMux I__735 (
            .O(N__4070),
            .I(N__4055));
    InMux I__734 (
            .O(N__4069),
            .I(N__4055));
    InMux I__733 (
            .O(N__4068),
            .I(N__4052));
    InMux I__732 (
            .O(N__4067),
            .I(N__4047));
    InMux I__731 (
            .O(N__4066),
            .I(N__4047));
    InMux I__730 (
            .O(N__4065),
            .I(N__4044));
    LocalMux I__729 (
            .O(N__4060),
            .I(\U400_SDRAM.N_139 ));
    LocalMux I__728 (
            .O(N__4055),
            .I(\U400_SDRAM.N_139 ));
    LocalMux I__727 (
            .O(N__4052),
            .I(\U400_SDRAM.N_139 ));
    LocalMux I__726 (
            .O(N__4047),
            .I(\U400_SDRAM.N_139 ));
    LocalMux I__725 (
            .O(N__4044),
            .I(\U400_SDRAM.N_139 ));
    CascadeMux I__724 (
            .O(N__4033),
            .I(\U400_SDRAM.N_141_cascade_ ));
    InMux I__723 (
            .O(N__4030),
            .I(N__4023));
    InMux I__722 (
            .O(N__4029),
            .I(N__4023));
    InMux I__721 (
            .O(N__4028),
            .I(N__4020));
    LocalMux I__720 (
            .O(N__4023),
            .I(N__4009));
    LocalMux I__719 (
            .O(N__4020),
            .I(N__4006));
    InMux I__718 (
            .O(N__4019),
            .I(N__4003));
    InMux I__717 (
            .O(N__4018),
            .I(N__3998));
    InMux I__716 (
            .O(N__4017),
            .I(N__3998));
    InMux I__715 (
            .O(N__4016),
            .I(N__3995));
    InMux I__714 (
            .O(N__4015),
            .I(N__3988));
    InMux I__713 (
            .O(N__4014),
            .I(N__3988));
    InMux I__712 (
            .O(N__4013),
            .I(N__3988));
    InMux I__711 (
            .O(N__4012),
            .I(N__3985));
    Span4Mux_h I__710 (
            .O(N__4009),
            .I(N__3976));
    Span4Mux_v I__709 (
            .O(N__4006),
            .I(N__3976));
    LocalMux I__708 (
            .O(N__4003),
            .I(N__3976));
    LocalMux I__707 (
            .O(N__3998),
            .I(N__3976));
    LocalMux I__706 (
            .O(N__3995),
            .I(\U400_SDRAM.REFRESH_COUNTER_RNIVV903Z0Z_8 ));
    LocalMux I__705 (
            .O(N__3988),
            .I(\U400_SDRAM.REFRESH_COUNTER_RNIVV903Z0Z_8 ));
    LocalMux I__704 (
            .O(N__3985),
            .I(\U400_SDRAM.REFRESH_COUNTER_RNIVV903Z0Z_8 ));
    Odrv4 I__703 (
            .O(N__3976),
            .I(\U400_SDRAM.REFRESH_COUNTER_RNIVV903Z0Z_8 ));
    InMux I__702 (
            .O(N__3967),
            .I(N__3960));
    InMux I__701 (
            .O(N__3966),
            .I(N__3960));
    InMux I__700 (
            .O(N__3965),
            .I(N__3955));
    LocalMux I__699 (
            .O(N__3960),
            .I(N__3952));
    CascadeMux I__698 (
            .O(N__3959),
            .I(N__3945));
    InMux I__697 (
            .O(N__3958),
            .I(N__3941));
    LocalMux I__696 (
            .O(N__3955),
            .I(N__3938));
    Span4Mux_h I__695 (
            .O(N__3952),
            .I(N__3935));
    InMux I__694 (
            .O(N__3951),
            .I(N__3930));
    InMux I__693 (
            .O(N__3950),
            .I(N__3930));
    InMux I__692 (
            .O(N__3949),
            .I(N__3927));
    InMux I__691 (
            .O(N__3948),
            .I(N__3924));
    InMux I__690 (
            .O(N__3945),
            .I(N__3919));
    InMux I__689 (
            .O(N__3944),
            .I(N__3919));
    LocalMux I__688 (
            .O(N__3941),
            .I(\U400_SDRAM.RAM_CYCLE_STARTZ0 ));
    Odrv4 I__687 (
            .O(N__3938),
            .I(\U400_SDRAM.RAM_CYCLE_STARTZ0 ));
    Odrv4 I__686 (
            .O(N__3935),
            .I(\U400_SDRAM.RAM_CYCLE_STARTZ0 ));
    LocalMux I__685 (
            .O(N__3930),
            .I(\U400_SDRAM.RAM_CYCLE_STARTZ0 ));
    LocalMux I__684 (
            .O(N__3927),
            .I(\U400_SDRAM.RAM_CYCLE_STARTZ0 ));
    LocalMux I__683 (
            .O(N__3924),
            .I(\U400_SDRAM.RAM_CYCLE_STARTZ0 ));
    LocalMux I__682 (
            .O(N__3919),
            .I(\U400_SDRAM.RAM_CYCLE_STARTZ0 ));
    InMux I__681 (
            .O(N__3904),
            .I(N__3901));
    LocalMux I__680 (
            .O(N__3901),
            .I(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_2_0 ));
    InMux I__679 (
            .O(N__3898),
            .I(N__3895));
    LocalMux I__678 (
            .O(N__3895),
            .I(\U400_SDRAM.SDRAM_COUNTER_s_0 ));
    CascadeMux I__677 (
            .O(N__3892),
            .I(\U400_SDRAM.N_181_cascade_ ));
    CascadeMux I__676 (
            .O(N__3889),
            .I(\U400_SDRAM.N_200_cascade_ ));
    InMux I__675 (
            .O(N__3886),
            .I(N__3883));
    LocalMux I__674 (
            .O(N__3883),
            .I(N__3880));
    Odrv4 I__673 (
            .O(N__3880),
            .I(\U400_SDRAM.N_199 ));
    CascadeMux I__672 (
            .O(N__3877),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_61_i_i_1_cascade_ ));
    InMux I__671 (
            .O(N__3874),
            .I(N__3870));
    InMux I__670 (
            .O(N__3873),
            .I(N__3866));
    LocalMux I__669 (
            .O(N__3870),
            .I(N__3863));
    InMux I__668 (
            .O(N__3869),
            .I(N__3860));
    LocalMux I__667 (
            .O(N__3866),
            .I(\U400_SDRAM.N_17 ));
    Odrv4 I__666 (
            .O(N__3863),
            .I(\U400_SDRAM.N_17 ));
    LocalMux I__665 (
            .O(N__3860),
            .I(\U400_SDRAM.N_17 ));
    InMux I__664 (
            .O(N__3853),
            .I(N__3850));
    LocalMux I__663 (
            .O(N__3850),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_0_1_1 ));
    InMux I__662 (
            .O(N__3847),
            .I(N__3842));
    InMux I__661 (
            .O(N__3846),
            .I(N__3839));
    InMux I__660 (
            .O(N__3845),
            .I(N__3836));
    LocalMux I__659 (
            .O(N__3842),
            .I(\U400_SDRAM.N_228 ));
    LocalMux I__658 (
            .O(N__3839),
            .I(\U400_SDRAM.N_228 ));
    LocalMux I__657 (
            .O(N__3836),
            .I(\U400_SDRAM.N_228 ));
    CascadeMux I__656 (
            .O(N__3829),
            .I(\U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5Z0Z_0_cascade_ ));
    InMux I__655 (
            .O(N__3826),
            .I(N__3823));
    LocalMux I__654 (
            .O(N__3823),
            .I(\U400_SDRAM.N_203 ));
    InMux I__653 (
            .O(N__3820),
            .I(N__3817));
    LocalMux I__652 (
            .O(N__3817),
            .I(\U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_i_0 ));
    CascadeMux I__651 (
            .O(N__3814),
            .I(\U400_SDRAM.N_176_cascade_ ));
    CascadeMux I__650 (
            .O(N__3811),
            .I(N__3808));
    InMux I__649 (
            .O(N__3808),
            .I(N__3805));
    LocalMux I__648 (
            .O(N__3805),
            .I(N__3801));
    InMux I__647 (
            .O(N__3804),
            .I(N__3798));
    Odrv4 I__646 (
            .O(N__3801),
            .I(\U400_SDRAM.CS1_ENZ0 ));
    LocalMux I__645 (
            .O(N__3798),
            .I(\U400_SDRAM.CS1_ENZ0 ));
    IoInMux I__644 (
            .O(N__3793),
            .I(N__3790));
    LocalMux I__643 (
            .O(N__3790),
            .I(N__3787));
    Odrv12 I__642 (
            .O(N__3787),
            .I(CS1n_c));
    CascadeMux I__641 (
            .O(N__3784),
            .I(N__3781));
    InMux I__640 (
            .O(N__3781),
            .I(N__3778));
    LocalMux I__639 (
            .O(N__3778),
            .I(N__3775));
    Span4Mux_h I__638 (
            .O(N__3775),
            .I(N__3772));
    Span4Mux_v I__637 (
            .O(N__3772),
            .I(N__3769));
    Span4Mux_v I__636 (
            .O(N__3769),
            .I(N__3766));
    Odrv4 I__635 (
            .O(N__3766),
            .I(A_c_26));
    IoInMux I__634 (
            .O(N__3763),
            .I(N__3760));
    LocalMux I__633 (
            .O(N__3760),
            .I(N__3757));
    Span12Mux_s0_v I__632 (
            .O(N__3757),
            .I(N__3754));
    Odrv12 I__631 (
            .O(N__3754),
            .I(MA_c_12));
    IoInMux I__630 (
            .O(N__3751),
            .I(N__3748));
    LocalMux I__629 (
            .O(N__3748),
            .I(N__3745));
    IoSpan4Mux I__628 (
            .O(N__3745),
            .I(N__3741));
    InMux I__627 (
            .O(N__3744),
            .I(N__3738));
    Span4Mux_s2_h I__626 (
            .O(N__3741),
            .I(N__3735));
    LocalMux I__625 (
            .O(N__3738),
            .I(N__3732));
    Odrv4 I__624 (
            .O(N__3735),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__623 (
            .O(N__3732),
            .I(CONSTANT_ONE_NET));
    IoInMux I__622 (
            .O(N__3727),
            .I(N__3724));
    LocalMux I__621 (
            .O(N__3724),
            .I(N__3721));
    Odrv12 I__620 (
            .O(N__3721),
            .I(UUBEn_c));
    InMux I__619 (
            .O(N__3718),
            .I(N__3715));
    LocalMux I__618 (
            .O(N__3715),
            .I(N__3709));
    InMux I__617 (
            .O(N__3714),
            .I(N__3706));
    InMux I__616 (
            .O(N__3713),
            .I(N__3701));
    InMux I__615 (
            .O(N__3712),
            .I(N__3701));
    Span4Mux_h I__614 (
            .O(N__3709),
            .I(N__3696));
    LocalMux I__613 (
            .O(N__3706),
            .I(N__3696));
    LocalMux I__612 (
            .O(N__3701),
            .I(\U400_SDRAM.TA_COUNTER23 ));
    Odrv4 I__611 (
            .O(N__3696),
            .I(\U400_SDRAM.TA_COUNTER23 ));
    InMux I__610 (
            .O(N__3691),
            .I(N__3688));
    LocalMux I__609 (
            .O(N__3688),
            .I(N__3682));
    InMux I__608 (
            .O(N__3687),
            .I(N__3676));
    InMux I__607 (
            .O(N__3686),
            .I(N__3676));
    InMux I__606 (
            .O(N__3685),
            .I(N__3672));
    Span4Mux_h I__605 (
            .O(N__3682),
            .I(N__3669));
    InMux I__604 (
            .O(N__3681),
            .I(N__3666));
    LocalMux I__603 (
            .O(N__3676),
            .I(N__3663));
    InMux I__602 (
            .O(N__3675),
            .I(N__3660));
    LocalMux I__601 (
            .O(N__3672),
            .I(\U400_SDRAM.TACKZ0 ));
    Odrv4 I__600 (
            .O(N__3669),
            .I(\U400_SDRAM.TACKZ0 ));
    LocalMux I__599 (
            .O(N__3666),
            .I(\U400_SDRAM.TACKZ0 ));
    Odrv4 I__598 (
            .O(N__3663),
            .I(\U400_SDRAM.TACKZ0 ));
    LocalMux I__597 (
            .O(N__3660),
            .I(\U400_SDRAM.TACKZ0 ));
    ClkMux I__596 (
            .O(N__3649),
            .I(N__3568));
    ClkMux I__595 (
            .O(N__3648),
            .I(N__3568));
    ClkMux I__594 (
            .O(N__3647),
            .I(N__3568));
    ClkMux I__593 (
            .O(N__3646),
            .I(N__3568));
    ClkMux I__592 (
            .O(N__3645),
            .I(N__3568));
    ClkMux I__591 (
            .O(N__3644),
            .I(N__3568));
    ClkMux I__590 (
            .O(N__3643),
            .I(N__3568));
    ClkMux I__589 (
            .O(N__3642),
            .I(N__3568));
    ClkMux I__588 (
            .O(N__3641),
            .I(N__3568));
    ClkMux I__587 (
            .O(N__3640),
            .I(N__3568));
    ClkMux I__586 (
            .O(N__3639),
            .I(N__3568));
    ClkMux I__585 (
            .O(N__3638),
            .I(N__3568));
    ClkMux I__584 (
            .O(N__3637),
            .I(N__3568));
    ClkMux I__583 (
            .O(N__3636),
            .I(N__3568));
    ClkMux I__582 (
            .O(N__3635),
            .I(N__3568));
    ClkMux I__581 (
            .O(N__3634),
            .I(N__3568));
    ClkMux I__580 (
            .O(N__3633),
            .I(N__3568));
    ClkMux I__579 (
            .O(N__3632),
            .I(N__3568));
    ClkMux I__578 (
            .O(N__3631),
            .I(N__3568));
    ClkMux I__577 (
            .O(N__3630),
            .I(N__3568));
    ClkMux I__576 (
            .O(N__3629),
            .I(N__3568));
    ClkMux I__575 (
            .O(N__3628),
            .I(N__3568));
    ClkMux I__574 (
            .O(N__3627),
            .I(N__3568));
    ClkMux I__573 (
            .O(N__3626),
            .I(N__3568));
    ClkMux I__572 (
            .O(N__3625),
            .I(N__3568));
    ClkMux I__571 (
            .O(N__3624),
            .I(N__3568));
    ClkMux I__570 (
            .O(N__3623),
            .I(N__3568));
    GlobalMux I__569 (
            .O(N__3568),
            .I(N__3565));
    gio2CtrlBuf I__568 (
            .O(N__3565),
            .I(CLK40_c_g));
    CEMux I__567 (
            .O(N__3562),
            .I(N__3559));
    LocalMux I__566 (
            .O(N__3559),
            .I(N__3556));
    Odrv12 I__565 (
            .O(N__3556),
            .I(\U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en_0 ));
    CascadeMux I__564 (
            .O(N__3553),
            .I(\U400_SDRAM.N_252_cascade_ ));
    CascadeMux I__563 (
            .O(N__3550),
            .I(N__3547));
    InMux I__562 (
            .O(N__3547),
            .I(N__3543));
    InMux I__561 (
            .O(N__3546),
            .I(N__3540));
    LocalMux I__560 (
            .O(N__3543),
            .I(\U400_SDRAM.RAM_CYCLEZ0 ));
    LocalMux I__559 (
            .O(N__3540),
            .I(\U400_SDRAM.RAM_CYCLEZ0 ));
    CascadeMux I__558 (
            .O(N__3535),
            .I(\U400_SDRAM.N_75_cascade_ ));
    InMux I__557 (
            .O(N__3532),
            .I(N__3529));
    LocalMux I__556 (
            .O(N__3529),
            .I(\U400_SDRAM.CS1_EN_0 ));
    CascadeMux I__555 (
            .O(N__3526),
            .I(\U400_SDRAM.CS1_EN_7_i_0_o3_0_cascade_ ));
    InMux I__554 (
            .O(N__3523),
            .I(N__3520));
    LocalMux I__553 (
            .O(N__3520),
            .I(\U400_SDRAM.N_159 ));
    InMux I__552 (
            .O(N__3517),
            .I(N__3511));
    InMux I__551 (
            .O(N__3516),
            .I(N__3511));
    LocalMux I__550 (
            .O(N__3511),
            .I(N__3508));
    Odrv12 I__549 (
            .O(N__3508),
            .I(A_c_23));
    CascadeMux I__548 (
            .O(N__3505),
            .I(N__3502));
    InMux I__547 (
            .O(N__3502),
            .I(N__3498));
    InMux I__546 (
            .O(N__3501),
            .I(N__3495));
    LocalMux I__545 (
            .O(N__3498),
            .I(\U400_SDRAM.CS0_ENZ0 ));
    LocalMux I__544 (
            .O(N__3495),
            .I(\U400_SDRAM.CS0_ENZ0 ));
    CascadeMux I__543 (
            .O(N__3490),
            .I(\U400_SDRAM.N_159_cascade_ ));
    InMux I__542 (
            .O(N__3487),
            .I(N__3484));
    LocalMux I__541 (
            .O(N__3484),
            .I(\U400_SDRAM.N_75 ));
    InMux I__540 (
            .O(N__3481),
            .I(N__3478));
    LocalMux I__539 (
            .O(N__3478),
            .I(\U400_SDRAM.CS0_EN_0 ));
    InMux I__538 (
            .O(N__3475),
            .I(N__3472));
    LocalMux I__537 (
            .O(N__3472),
            .I(N__3468));
    InMux I__536 (
            .O(N__3471),
            .I(N__3465));
    Odrv12 I__535 (
            .O(N__3468),
            .I(\U400_SDRAM.N_250 ));
    LocalMux I__534 (
            .O(N__3465),
            .I(\U400_SDRAM.N_250 ));
    InMux I__533 (
            .O(N__3460),
            .I(N__3457));
    LocalMux I__532 (
            .O(N__3457),
            .I(\U400_SDRAM.N_189 ));
    CascadeMux I__531 (
            .O(N__3454),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_1_32_i_0_i_1_1_cascade_ ));
    CascadeMux I__530 (
            .O(N__3451),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_1_32_i_0_i_1_cascade_ ));
    CascadeMux I__529 (
            .O(N__3448),
            .I(N__3445));
    InMux I__528 (
            .O(N__3445),
            .I(N__3440));
    InMux I__527 (
            .O(N__3444),
            .I(N__3435));
    InMux I__526 (
            .O(N__3443),
            .I(N__3435));
    LocalMux I__525 (
            .O(N__3440),
            .I(\U400_SDRAM.N_128 ));
    LocalMux I__524 (
            .O(N__3435),
            .I(\U400_SDRAM.N_128 ));
    InMux I__523 (
            .O(N__3430),
            .I(N__3427));
    LocalMux I__522 (
            .O(N__3427),
            .I(\U400_SDRAM.N_185 ));
    SRMux I__521 (
            .O(N__3424),
            .I(N__3420));
    SRMux I__520 (
            .O(N__3423),
            .I(N__3417));
    LocalMux I__519 (
            .O(N__3420),
            .I(N__3412));
    LocalMux I__518 (
            .O(N__3417),
            .I(N__3412));
    Odrv4 I__517 (
            .O(N__3412),
            .I(\U400_SDRAM.SDRAM_COUNTER_RNIJKCA2Z0Z_1 ));
    InMux I__516 (
            .O(N__3409),
            .I(N__3405));
    InMux I__515 (
            .O(N__3408),
            .I(N__3402));
    LocalMux I__514 (
            .O(N__3405),
            .I(N__3399));
    LocalMux I__513 (
            .O(N__3402),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_3 ));
    Odrv4 I__512 (
            .O(N__3399),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__511 (
            .O(N__3394),
            .I(N__3390));
    InMux I__510 (
            .O(N__3393),
            .I(N__3387));
    LocalMux I__509 (
            .O(N__3390),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_2 ));
    LocalMux I__508 (
            .O(N__3387),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_2 ));
    CascadeMux I__507 (
            .O(N__3382),
            .I(N__3378));
    InMux I__506 (
            .O(N__3381),
            .I(N__3375));
    InMux I__505 (
            .O(N__3378),
            .I(N__3372));
    LocalMux I__504 (
            .O(N__3375),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__503 (
            .O(N__3372),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__502 (
            .O(N__3367),
            .I(N__3362));
    InMux I__501 (
            .O(N__3366),
            .I(N__3359));
    InMux I__500 (
            .O(N__3365),
            .I(N__3356));
    LocalMux I__499 (
            .O(N__3362),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__498 (
            .O(N__3359),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__497 (
            .O(N__3356),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_1 ));
    InMux I__496 (
            .O(N__3349),
            .I(N__3346));
    LocalMux I__495 (
            .O(N__3346),
            .I(N__3336));
    InMux I__494 (
            .O(N__3345),
            .I(N__3331));
    InMux I__493 (
            .O(N__3344),
            .I(N__3331));
    InMux I__492 (
            .O(N__3343),
            .I(N__3328));
    InMux I__491 (
            .O(N__3342),
            .I(N__3319));
    InMux I__490 (
            .O(N__3341),
            .I(N__3319));
    InMux I__489 (
            .O(N__3340),
            .I(N__3319));
    InMux I__488 (
            .O(N__3339),
            .I(N__3319));
    Odrv4 I__487 (
            .O(N__3336),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_0 ));
    LocalMux I__486 (
            .O(N__3331),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_0 ));
    LocalMux I__485 (
            .O(N__3328),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_0 ));
    LocalMux I__484 (
            .O(N__3319),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_0 ));
    InMux I__483 (
            .O(N__3310),
            .I(N__3305));
    InMux I__482 (
            .O(N__3309),
            .I(N__3300));
    InMux I__481 (
            .O(N__3308),
            .I(N__3300));
    LocalMux I__480 (
            .O(N__3305),
            .I(\U400_SDRAM.BURSTZ0 ));
    LocalMux I__479 (
            .O(N__3300),
            .I(\U400_SDRAM.BURSTZ0 ));
    InMux I__478 (
            .O(N__3295),
            .I(N__3292));
    LocalMux I__477 (
            .O(N__3292),
            .I(\U400_SDRAM.TA_EN11_m ));
    InMux I__476 (
            .O(N__3289),
            .I(N__3285));
    InMux I__475 (
            .O(N__3288),
            .I(N__3282));
    LocalMux I__474 (
            .O(N__3285),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__473 (
            .O(N__3282),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_6 ));
    CascadeMux I__472 (
            .O(N__3277),
            .I(N__3272));
    InMux I__471 (
            .O(N__3276),
            .I(N__3266));
    InMux I__470 (
            .O(N__3275),
            .I(N__3266));
    InMux I__469 (
            .O(N__3272),
            .I(N__3263));
    InMux I__468 (
            .O(N__3271),
            .I(N__3260));
    LocalMux I__467 (
            .O(N__3266),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_0 ));
    LocalMux I__466 (
            .O(N__3263),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_0 ));
    LocalMux I__465 (
            .O(N__3260),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_0 ));
    CascadeMux I__464 (
            .O(N__3253),
            .I(N__3249));
    InMux I__463 (
            .O(N__3252),
            .I(N__3246));
    InMux I__462 (
            .O(N__3249),
            .I(N__3243));
    LocalMux I__461 (
            .O(N__3246),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__460 (
            .O(N__3243),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__459 (
            .O(N__3238),
            .I(N__3234));
    InMux I__458 (
            .O(N__3237),
            .I(N__3231));
    LocalMux I__457 (
            .O(N__3234),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__456 (
            .O(N__3231),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_5 ));
    CascadeMux I__455 (
            .O(N__3226),
            .I(\U400_SDRAM.N_205_cascade_ ));
    CascadeMux I__454 (
            .O(N__3223),
            .I(N__3220));
    InMux I__453 (
            .O(N__3220),
            .I(N__3217));
    LocalMux I__452 (
            .O(N__3217),
            .I(\U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en ));
    InMux I__451 (
            .O(N__3214),
            .I(N__3211));
    LocalMux I__450 (
            .O(N__3211),
            .I(\U400_SDRAM.un1_REFRESH_COUNTERlto7_4 ));
    InMux I__449 (
            .O(N__3208),
            .I(N__3204));
    InMux I__448 (
            .O(N__3207),
            .I(N__3201));
    LocalMux I__447 (
            .O(N__3204),
            .I(N__3198));
    LocalMux I__446 (
            .O(N__3201),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_8 ));
    Odrv4 I__445 (
            .O(N__3198),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_8 ));
    InMux I__444 (
            .O(N__3193),
            .I(N__3190));
    LocalMux I__443 (
            .O(N__3190),
            .I(\U400_SDRAM.un1_REFRESH_COUNTERlto7_5 ));
    InMux I__442 (
            .O(N__3187),
            .I(N__3183));
    InMux I__441 (
            .O(N__3186),
            .I(N__3180));
    LocalMux I__440 (
            .O(N__3183),
            .I(\U400_SDRAM.N_255 ));
    LocalMux I__439 (
            .O(N__3180),
            .I(\U400_SDRAM.N_255 ));
    CascadeMux I__438 (
            .O(N__3175),
            .I(\U400_SDRAM.TACK_7_iv_i_i_0_cascade_ ));
    InMux I__437 (
            .O(N__3172),
            .I(N__3169));
    LocalMux I__436 (
            .O(N__3169),
            .I(\U400_SDRAM.TACK_7_iv_i_i_1 ));
    InMux I__435 (
            .O(N__3166),
            .I(N__3163));
    LocalMux I__434 (
            .O(N__3163),
            .I(\U400_SDRAM.N_15 ));
    InMux I__433 (
            .O(N__3160),
            .I(N__3157));
    LocalMux I__432 (
            .O(N__3157),
            .I(\U400_SDRAM.RAM_CYCLE_e_1 ));
    InMux I__431 (
            .O(N__3154),
            .I(N__3149));
    InMux I__430 (
            .O(N__3153),
            .I(N__3144));
    InMux I__429 (
            .O(N__3152),
            .I(N__3144));
    LocalMux I__428 (
            .O(N__3149),
            .I(\U400_SDRAM.N_6 ));
    LocalMux I__427 (
            .O(N__3144),
            .I(\U400_SDRAM.N_6 ));
    InMux I__426 (
            .O(N__3139),
            .I(N__3136));
    LocalMux I__425 (
            .O(N__3136),
            .I(N__3133));
    Span4Mux_v I__424 (
            .O(N__3133),
            .I(N__3130));
    Span4Mux_h I__423 (
            .O(N__3130),
            .I(N__3127));
    Odrv4 I__422 (
            .O(N__3127),
            .I(RnW_c));
    IoInMux I__421 (
            .O(N__3124),
            .I(N__3121));
    LocalMux I__420 (
            .O(N__3121),
            .I(N__3118));
    IoSpan4Mux I__419 (
            .O(N__3118),
            .I(N__3115));
    Span4Mux_s3_h I__418 (
            .O(N__3115),
            .I(N__3112));
    Odrv4 I__417 (
            .O(N__3112),
            .I(CS0n_c));
    CascadeMux I__416 (
            .O(N__3109),
            .I(N__3106));
    InMux I__415 (
            .O(N__3106),
            .I(N__3103));
    LocalMux I__414 (
            .O(N__3103),
            .I(N__3100));
    Span4Mux_v I__413 (
            .O(N__3100),
            .I(N__3097));
    Sp12to4 I__412 (
            .O(N__3097),
            .I(N__3094));
    Odrv12 I__411 (
            .O(N__3094),
            .I(A_c_19));
    IoInMux I__410 (
            .O(N__3091),
            .I(N__3088));
    LocalMux I__409 (
            .O(N__3088),
            .I(N__3085));
    Odrv12 I__408 (
            .O(N__3085),
            .I(MA_c_9));
    InMux I__407 (
            .O(N__3082),
            .I(N__3074));
    InMux I__406 (
            .O(N__3081),
            .I(N__3071));
    InMux I__405 (
            .O(N__3080),
            .I(N__3062));
    InMux I__404 (
            .O(N__3079),
            .I(N__3062));
    InMux I__403 (
            .O(N__3078),
            .I(N__3062));
    InMux I__402 (
            .O(N__3077),
            .I(N__3062));
    LocalMux I__401 (
            .O(N__3074),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_1 ));
    LocalMux I__400 (
            .O(N__3071),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_1 ));
    LocalMux I__399 (
            .O(N__3062),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_1 ));
    CascadeMux I__398 (
            .O(N__3055),
            .I(N__3050));
    CascadeMux I__397 (
            .O(N__3054),
            .I(N__3045));
    CascadeMux I__396 (
            .O(N__3053),
            .I(N__3042));
    InMux I__395 (
            .O(N__3050),
            .I(N__3039));
    InMux I__394 (
            .O(N__3049),
            .I(N__3032));
    InMux I__393 (
            .O(N__3048),
            .I(N__3032));
    InMux I__392 (
            .O(N__3045),
            .I(N__3032));
    InMux I__391 (
            .O(N__3042),
            .I(N__3029));
    LocalMux I__390 (
            .O(N__3039),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_3 ));
    LocalMux I__389 (
            .O(N__3032),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_3 ));
    LocalMux I__388 (
            .O(N__3029),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_3 ));
    InMux I__387 (
            .O(N__3022),
            .I(N__3018));
    InMux I__386 (
            .O(N__3021),
            .I(N__3015));
    LocalMux I__385 (
            .O(N__3018),
            .I(\U400_SDRAM.TA_COUNTER_0_sqmuxa ));
    LocalMux I__384 (
            .O(N__3015),
            .I(\U400_SDRAM.TA_COUNTER_0_sqmuxa ));
    InMux I__383 (
            .O(N__3010),
            .I(N__3006));
    InMux I__382 (
            .O(N__3009),
            .I(N__3003));
    LocalMux I__381 (
            .O(N__3006),
            .I(\U400_SDRAM.TA_COUNTER27 ));
    LocalMux I__380 (
            .O(N__3003),
            .I(\U400_SDRAM.TA_COUNTER27 ));
    CascadeMux I__379 (
            .O(N__2998),
            .I(\U400_SDRAM.TA_COUNTER_0_sqmuxa_cascade_ ));
    CascadeMux I__378 (
            .O(N__2995),
            .I(\U400_SDRAM.un1_SDRAM_COUNTER52_2_0_i_1_cascade_ ));
    InMux I__377 (
            .O(N__2992),
            .I(N__2986));
    InMux I__376 (
            .O(N__2991),
            .I(N__2986));
    LocalMux I__375 (
            .O(N__2986),
            .I(\U400_SDRAM.N_23 ));
    InMux I__374 (
            .O(N__2983),
            .I(\U400_SDRAM.un2_REFRESH_COUNTER_cry_1 ));
    InMux I__373 (
            .O(N__2980),
            .I(\U400_SDRAM.un2_REFRESH_COUNTER_cry_2 ));
    InMux I__372 (
            .O(N__2977),
            .I(\U400_SDRAM.un2_REFRESH_COUNTER_cry_3 ));
    InMux I__371 (
            .O(N__2974),
            .I(\U400_SDRAM.un2_REFRESH_COUNTER_cry_4 ));
    InMux I__370 (
            .O(N__2971),
            .I(\U400_SDRAM.un2_REFRESH_COUNTER_cry_5 ));
    InMux I__369 (
            .O(N__2968),
            .I(\U400_SDRAM.un2_REFRESH_COUNTER_cry_6 ));
    InMux I__368 (
            .O(N__2965),
            .I(\U400_SDRAM.un2_REFRESH_COUNTER_cry_7 ));
    CascadeMux I__367 (
            .O(N__2962),
            .I(N__2955));
    InMux I__366 (
            .O(N__2961),
            .I(N__2951));
    InMux I__365 (
            .O(N__2960),
            .I(N__2948));
    InMux I__364 (
            .O(N__2959),
            .I(N__2939));
    InMux I__363 (
            .O(N__2958),
            .I(N__2939));
    InMux I__362 (
            .O(N__2955),
            .I(N__2939));
    InMux I__361 (
            .O(N__2954),
            .I(N__2939));
    LocalMux I__360 (
            .O(N__2951),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_2 ));
    LocalMux I__359 (
            .O(N__2948),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_2 ));
    LocalMux I__358 (
            .O(N__2939),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_2 ));
    InMux I__357 (
            .O(N__2932),
            .I(N__2929));
    LocalMux I__356 (
            .O(N__2929),
            .I(\U400_SDRAM.un1_TA_COUNTER26_2_0 ));
    IoInMux I__355 (
            .O(N__2926),
            .I(N__2923));
    LocalMux I__354 (
            .O(N__2923),
            .I(N__2919));
    CascadeMux I__353 (
            .O(N__2922),
            .I(N__2916));
    Span12Mux_s7_h I__352 (
            .O(N__2919),
            .I(N__2913));
    InMux I__351 (
            .O(N__2916),
            .I(N__2910));
    Odrv12 I__350 (
            .O(N__2913),
            .I(TA_OUT));
    LocalMux I__349 (
            .O(N__2910),
            .I(TA_OUT));
    CascadeMux I__348 (
            .O(N__2905),
            .I(\U400_SDRAM.N_208_cascade_ ));
    CascadeMux I__347 (
            .O(N__2902),
            .I(N__2899));
    InMux I__346 (
            .O(N__2899),
            .I(N__2896));
    LocalMux I__345 (
            .O(N__2896),
            .I(\U400_SDRAM.un1_SDRAM_COUNTER52_4_0_i_2 ));
    IoInMux I__344 (
            .O(N__2893),
            .I(N__2890));
    LocalMux I__343 (
            .O(N__2890),
            .I(N__2887));
    Span4Mux_s3_h I__342 (
            .O(N__2887),
            .I(N__2884));
    Odrv4 I__341 (
            .O(N__2884),
            .I(RASn_c));
    IoInMux I__340 (
            .O(N__2881),
            .I(N__2878));
    LocalMux I__339 (
            .O(N__2878),
            .I(N__2875));
    Odrv12 I__338 (
            .O(N__2875),
            .I(CASn_c));
    IoInMux I__337 (
            .O(N__2872),
            .I(N__2869));
    LocalMux I__336 (
            .O(N__2869),
            .I(N__2866));
    Odrv12 I__335 (
            .O(N__2866),
            .I(WEn_c));
    InMux I__334 (
            .O(N__2863),
            .I(N__2860));
    LocalMux I__333 (
            .O(N__2860),
            .I(N__2857));
    Span4Mux_h I__332 (
            .O(N__2857),
            .I(N__2854));
    Sp12to4 I__331 (
            .O(N__2854),
            .I(N__2851));
    Span12Mux_v I__330 (
            .O(N__2851),
            .I(N__2848));
    Odrv12 I__329 (
            .O(N__2848),
            .I(A_c_24));
    CascadeMux I__328 (
            .O(N__2845),
            .I(N__2842));
    InMux I__327 (
            .O(N__2842),
            .I(N__2839));
    LocalMux I__326 (
            .O(N__2839),
            .I(N__2836));
    Span12Mux_s10_v I__325 (
            .O(N__2836),
            .I(N__2833));
    Odrv12 I__324 (
            .O(N__2833),
            .I(A_c_18));
    IoInMux I__323 (
            .O(N__2830),
            .I(N__2827));
    LocalMux I__322 (
            .O(N__2827),
            .I(N__2824));
    Span4Mux_s1_v I__321 (
            .O(N__2824),
            .I(N__2821));
    Odrv4 I__320 (
            .O(N__2821),
            .I(MA_c_8));
    InMux I__319 (
            .O(N__2818),
            .I(N__2815));
    LocalMux I__318 (
            .O(N__2815),
            .I(N__2812));
    Span4Mux_v I__317 (
            .O(N__2812),
            .I(N__2809));
    Odrv4 I__316 (
            .O(N__2809),
            .I(A_c_17));
    InMux I__315 (
            .O(N__2806),
            .I(N__2803));
    LocalMux I__314 (
            .O(N__2803),
            .I(N__2800));
    Odrv12 I__313 (
            .O(N__2800),
            .I(A_c_9));
    IoInMux I__312 (
            .O(N__2797),
            .I(N__2794));
    LocalMux I__311 (
            .O(N__2794),
            .I(N__2791));
    Odrv12 I__310 (
            .O(N__2791),
            .I(MA_c_7));
    InMux I__309 (
            .O(N__2788),
            .I(N__2785));
    LocalMux I__308 (
            .O(N__2785),
            .I(N__2782));
    Odrv12 I__307 (
            .O(N__2782),
            .I(A_c_8));
    CascadeMux I__306 (
            .O(N__2779),
            .I(N__2776));
    InMux I__305 (
            .O(N__2776),
            .I(N__2773));
    LocalMux I__304 (
            .O(N__2773),
            .I(N__2770));
    Span4Mux_v I__303 (
            .O(N__2770),
            .I(N__2767));
    Span4Mux_v I__302 (
            .O(N__2767),
            .I(N__2764));
    Odrv4 I__301 (
            .O(N__2764),
            .I(A_c_16));
    IoInMux I__300 (
            .O(N__2761),
            .I(N__2758));
    LocalMux I__299 (
            .O(N__2758),
            .I(N__2755));
    Odrv12 I__298 (
            .O(N__2755),
            .I(MA_c_6));
    CascadeMux I__297 (
            .O(N__2752),
            .I(\U400_SDRAM.TA_COUNTER23_cascade_ ));
    InMux I__296 (
            .O(N__2749),
            .I(N__2746));
    LocalMux I__295 (
            .O(N__2746),
            .I(\U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0 ));
    CascadeMux I__294 (
            .O(N__2743),
            .I(\U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0_cascade_ ));
    InMux I__293 (
            .O(N__2740),
            .I(N__2737));
    LocalMux I__292 (
            .O(N__2737),
            .I(\U400_SDRAM.CO1 ));
    CascadeMux I__291 (
            .O(N__2734),
            .I(\U400_SDRAM.CO1_cascade_ ));
    CascadeMux I__290 (
            .O(N__2731),
            .I(N__2728));
    InMux I__289 (
            .O(N__2728),
            .I(N__2725));
    LocalMux I__288 (
            .O(N__2725),
            .I(N__2722));
    Span4Mux_v I__287 (
            .O(N__2722),
            .I(N__2719));
    Odrv4 I__286 (
            .O(N__2719),
            .I(A_c_21));
    IoInMux I__285 (
            .O(N__2716),
            .I(N__2713));
    LocalMux I__284 (
            .O(N__2713),
            .I(N__2710));
    Span4Mux_s3_h I__283 (
            .O(N__2710),
            .I(N__2707));
    Span4Mux_v I__282 (
            .O(N__2707),
            .I(N__2703));
    InMux I__281 (
            .O(N__2706),
            .I(N__2700));
    Odrv4 I__280 (
            .O(N__2703),
            .I(BANK0_c));
    LocalMux I__279 (
            .O(N__2700),
            .I(BANK0_c));
    CascadeMux I__278 (
            .O(N__2695),
            .I(N__2692));
    InMux I__277 (
            .O(N__2692),
            .I(N__2689));
    LocalMux I__276 (
            .O(N__2689),
            .I(N__2686));
    Span4Mux_h I__275 (
            .O(N__2686),
            .I(N__2683));
    Span4Mux_v I__274 (
            .O(N__2683),
            .I(N__2680));
    Odrv4 I__273 (
            .O(N__2680),
            .I(A_c_22));
    IoInMux I__272 (
            .O(N__2677),
            .I(N__2674));
    LocalMux I__271 (
            .O(N__2674),
            .I(N__2671));
    Span4Mux_s3_h I__270 (
            .O(N__2671),
            .I(N__2668));
    Span4Mux_v I__269 (
            .O(N__2668),
            .I(N__2664));
    InMux I__268 (
            .O(N__2667),
            .I(N__2661));
    Odrv4 I__267 (
            .O(N__2664),
            .I(BANK1_c));
    LocalMux I__266 (
            .O(N__2661),
            .I(BANK1_c));
    CascadeMux I__265 (
            .O(N__2656),
            .I(\U400_SDRAM.un1_SDRAM_COUNTER52_4_0_i_a3_0_cascade_ ));
    InMux I__264 (
            .O(N__2653),
            .I(N__2650));
    LocalMux I__263 (
            .O(N__2650),
            .I(\U400_SDRAM.un1_SDRAM_COUNTER52_4_0_i_1 ));
    IoInMux I__262 (
            .O(N__2647),
            .I(N__2644));
    LocalMux I__261 (
            .O(N__2644),
            .I(N__2641));
    Odrv4 I__260 (
            .O(N__2641),
            .I(RESETn_c_i));
    InMux I__259 (
            .O(N__2638),
            .I(N__2635));
    LocalMux I__258 (
            .O(N__2635),
            .I(N__2632));
    Span4Mux_h I__257 (
            .O(N__2632),
            .I(N__2629));
    Odrv4 I__256 (
            .O(N__2629),
            .I(A_c_30));
    InMux I__255 (
            .O(N__2626),
            .I(N__2623));
    LocalMux I__254 (
            .O(N__2623),
            .I(N__2620));
    Span12Mux_s10_h I__253 (
            .O(N__2620),
            .I(N__2617));
    Odrv12 I__252 (
            .O(N__2617),
            .I(A_c_29));
    CascadeMux I__251 (
            .O(N__2614),
            .I(N__2611));
    InMux I__250 (
            .O(N__2611),
            .I(N__2608));
    LocalMux I__249 (
            .O(N__2608),
            .I(A_c_28));
    InMux I__248 (
            .O(N__2605),
            .I(N__2602));
    LocalMux I__247 (
            .O(N__2602),
            .I(N__2599));
    Span4Mux_s1_v I__246 (
            .O(N__2599),
            .I(N__2596));
    Odrv4 I__245 (
            .O(N__2596),
            .I(A_c_27));
    CascadeMux I__244 (
            .O(N__2593),
            .I(\U400_SDRAM.TA_COUNTER_7_f1_0_0_cascade_ ));
    CascadeMux I__243 (
            .O(N__2590),
            .I(\U400_SDRAM.un1_TA_COUNTER26_0_cascade_ ));
    IoInMux I__242 (
            .O(N__2587),
            .I(N__2584));
    LocalMux I__241 (
            .O(N__2584),
            .I(N__2581));
    IoSpan4Mux I__240 (
            .O(N__2581),
            .I(N__2578));
    IoSpan4Mux I__239 (
            .O(N__2578),
            .I(N__2575));
    Span4Mux_s2_h I__238 (
            .O(N__2575),
            .I(N__2572));
    Sp12to4 I__237 (
            .O(N__2572),
            .I(N__2569));
    Odrv12 I__236 (
            .O(N__2569),
            .I(CLK40_ibuf_gb_io_gb_input));
    INV \INVU400_SDRAM.MA_2C  (
            .O(\INVU400_SDRAM.MA_2C_net ),
            .I(N__3649));
    INV \INVU400_SDRAM.MA_3C  (
            .O(\INVU400_SDRAM.MA_3C_net ),
            .I(N__3646));
    INV \INVU400_SDRAM.MA_0C  (
            .O(\INVU400_SDRAM.MA_0C_net ),
            .I(N__3648));
    INV \INVU400_SDRAM.SDRAM_COUNTER_2C  (
            .O(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .I(N__3638));
    INV \INVU400_SDRAM.SDRAM_COUNTER_1C  (
            .O(\INVU400_SDRAM.SDRAM_COUNTER_1C_net ),
            .I(N__3642));
    INV \INVU400_SDRAM.MA_4C  (
            .O(\INVU400_SDRAM.MA_4C_net ),
            .I(N__3647));
    INV \INVU400_SDRAM.MA_11C  (
            .O(\INVU400_SDRAM.MA_11C_net ),
            .I(N__3632));
    INV \INVU400_SDRAM.SDRAM_COUNTER_0C  (
            .O(\INVU400_SDRAM.SDRAM_COUNTER_0C_net ),
            .I(N__3625));
    INV \INVU400_SDRAM.SDRAM_COUNTER_3C  (
            .O(\INVU400_SDRAM.SDRAM_COUNTER_3C_net ),
            .I(N__3637));
    INV \INVU400_SDRAM.SDRAM_CMD_2C  (
            .O(\INVU400_SDRAM.SDRAM_CMD_2C_net ),
            .I(N__3641));
    INV \INVU400_SDRAM.CS1nC  (
            .O(\INVU400_SDRAM.CS1nC_net ),
            .I(N__3629));
    INV \INVU400_SDRAM.SDRAM_CMD_0C  (
            .O(\INVU400_SDRAM.SDRAM_CMD_0C_net ),
            .I(N__3636));
    INV \INVU400_SDRAM.SDRAM_CMD_1C  (
            .O(\INVU400_SDRAM.SDRAM_CMD_1C_net ),
            .I(N__3640));
    INV \INVU400_SDRAM.REFRESH_COUNTER_0C  (
            .O(\INVU400_SDRAM.REFRESH_COUNTER_0C_net ),
            .I(N__3645));
    INV \INVU400_SDRAM.CS0_ENC  (
            .O(\INVU400_SDRAM.CS0_ENC_net ),
            .I(N__3624));
    INV \INVU400_SDRAM.RAM_CYCLEC  (
            .O(\INVU400_SDRAM.RAM_CYCLEC_net ),
            .I(N__3628));
    INV \INVU400_SDRAM.BURSTC  (
            .O(\INVU400_SDRAM.BURSTC_net ),
            .I(N__3635));
    INV \INVU400_SDRAM.REFRESH_COUNTER_2C  (
            .O(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .I(N__3643));
    INV \INVU400_SDRAM.MA_6C  (
            .O(\INVU400_SDRAM.MA_6C_net ),
            .I(N__3633));
    INV \INVU400_SDRAM.MA_8C  (
            .O(\INVU400_SDRAM.MA_8C_net ),
            .I(N__3626));
    INV \INVU400_SDRAM.RASnC  (
            .O(\INVU400_SDRAM.RASnC_net ),
            .I(N__3623));
    INV \INVU400_SDRAM.BANK0C  (
            .O(\INVU400_SDRAM.BANK0C_net ),
            .I(N__3627));
    defparam IN_MUX_bfv_5_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_3_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_8_0_));
    ICE_GB CLK40_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__2587),
            .GLOBALBUFFEROUTPUT(CLK40_c_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__2647),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_2_8_5.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_2_8_5.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_2_8_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_2_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5555),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_0_a3_3_LC_4_1_3 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_0_a3_3_LC_4_1_3 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_0_a3_3_LC_4_1_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U400_ADDRESS_DECODE.RAM_SPACE_0_a3_3_LC_4_1_3  (
            .in0(N__2638),
            .in1(N__2626),
            .in2(N__2614),
            .in3(N__2605),
            .lcout(U400_ADDRESS_DECODE_RAM_SPACE_0_a3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_4_4_1 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_4_4_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_4_4_1 .LUT_INIT=16'b0010001001100110;
    LogicCell40 \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_4_4_1  (
            .in0(N__3345),
            .in1(N__3712),
            .in2(_gnd_net_),
            .in3(N__3686),
            .lcout(),
            .ltout(\U400_SDRAM.TA_COUNTER_7_f1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_0_LC_4_4_2 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_0_LC_4_4_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_0_LC_4_4_2 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \U400_SDRAM.TA_COUNTER_0_LC_4_4_2  (
            .in0(N__5522),
            .in1(_gnd_net_),
            .in2(N__2593),
            .in3(N__3022),
            .lcout(\U400_SDRAM.TA_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3634),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_OUT_RNO_2_LC_4_4_6 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_OUT_RNO_2_LC_4_4_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_OUT_RNO_2_LC_4_4_6 .LUT_INIT=16'b1111111011110100;
    LogicCell40 \U400_SDRAM.TA_OUT_RNO_2_LC_4_4_6  (
            .in0(N__2960),
            .in1(N__3082),
            .in2(N__3055),
            .in3(N__3344),
            .lcout(),
            .ltout(\U400_SDRAM.un1_TA_COUNTER26_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_OUT_RNO_1_LC_4_4_7 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_OUT_RNO_1_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_OUT_RNO_1_LC_4_4_7 .LUT_INIT=16'b0000111100000011;
    LogicCell40 \U400_SDRAM.TA_OUT_RNO_1_LC_4_4_7  (
            .in0(_gnd_net_),
            .in1(N__3713),
            .in2(N__2590),
            .in3(N__3687),
            .lcout(\U400_SDRAM.un1_TA_COUNTER26_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_RNIAJGG1_3_LC_4_5_0 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_RNIAJGG1_3_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_COUNTER_RNIAJGG1_3_LC_4_5_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_RNIAJGG1_3_LC_4_5_0  (
            .in0(N__3339),
            .in1(N__2954),
            .in2(N__3054),
            .in3(N__3077),
            .lcout(\U400_SDRAM.TA_COUNTER27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_1_LC_4_5_2 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_1_LC_4_5_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_1_LC_4_5_2 .LUT_INIT=16'b0110000000000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_1_LC_4_5_2  (
            .in0(N__3342),
            .in1(N__3080),
            .in2(N__5557),
            .in3(N__2749),
            .lcout(\U400_SDRAM.TA_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3630),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_RNIAJGG1_0_3_LC_4_5_3 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_RNIAJGG1_0_3_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_COUNTER_RNIAJGG1_0_3_LC_4_5_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U400_SDRAM.TA_COUNTER_RNIAJGG1_0_3_LC_4_5_3  (
            .in0(N__3078),
            .in1(N__3048),
            .in2(N__2962),
            .in3(N__3340),
            .lcout(\U400_SDRAM.TA_COUNTER23 ),
            .ltout(\U400_SDRAM.TA_COUNTER23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNI0LUG4_LC_4_5_4 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNI0LUG4_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNI0LUG4_LC_4_5_4 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \U400_SDRAM.TACK_RNI0LUG4_LC_4_5_4  (
            .in0(N__3010),
            .in1(N__3681),
            .in2(N__2752),
            .in3(N__3021),
            .lcout(\U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0 ),
            .ltout(\U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_2_LC_4_5_5 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_2_LC_4_5_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_2_LC_4_5_5 .LUT_INIT=16'b0100000010000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_2_LC_4_5_5  (
            .in0(N__2958),
            .in1(N__5551),
            .in2(N__2743),
            .in3(N__2740),
            .lcout(\U400_SDRAM.TA_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3630),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_RNIJ78O_1_LC_4_5_6 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_RNIJ78O_1_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_COUNTER_RNIJ78O_1_LC_4_5_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_RNIJ78O_1_LC_4_5_6  (
            .in0(N__3341),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3079),
            .lcout(\U400_SDRAM.CO1 ),
            .ltout(\U400_SDRAM.CO1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_3_LC_4_5_7 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_3_LC_4_5_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_3_LC_4_5_7 .LUT_INIT=16'b0100110010000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_3_LC_4_5_7  (
            .in0(N__2959),
            .in1(N__5552),
            .in2(N__2734),
            .in3(N__3049),
            .lcout(\U400_SDRAM.TA_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3630),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.BANK0_LC_4_6_0 .C_ON=1'b0;
    defparam \U400_SDRAM.BANK0_LC_4_6_0 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.BANK0_LC_4_6_0 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \U400_SDRAM.BANK0_LC_4_6_0  (
            .in0(N__2991),
            .in1(N__2706),
            .in2(N__2731),
            .in3(N__3967),
            .lcout(BANK0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.BANK0C_net ),
            .ce(),
            .sr(N__5922));
    defparam \U400_SDRAM.BANK1_LC_4_6_1 .C_ON=1'b0;
    defparam \U400_SDRAM.BANK1_LC_4_6_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.BANK1_LC_4_6_1 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \U400_SDRAM.BANK1_LC_4_6_1  (
            .in0(N__3966),
            .in1(N__2667),
            .in2(N__2695),
            .in3(N__2992),
            .lcout(BANK1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.BANK0C_net ),
            .ce(),
            .sr(N__5922));
    defparam \U400_SDRAM.TACK_LC_4_6_2 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_LC_4_6_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TACK_LC_4_6_2 .LUT_INIT=16'b1111110100000001;
    LogicCell40 \U400_SDRAM.TACK_LC_4_6_2  (
            .in0(N__3166),
            .in1(N__2653),
            .in2(N__2902),
            .in3(N__3685),
            .lcout(\U400_SDRAM.TACKZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.BANK0C_net ),
            .ce(),
            .sr(N__5922));
    defparam \U400_SDRAM.TACK_RNO_6_LC_4_7_0 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_6_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_6_LC_4_7_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U400_SDRAM.TACK_RNO_6_LC_4_7_0  (
            .in0(N__5079),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4959),
            .lcout(),
            .ltout(\U400_SDRAM.un1_SDRAM_COUNTER52_4_0_i_a3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_1_LC_4_7_1 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_1_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_1_LC_4_7_1 .LUT_INIT=16'b1111111101100000;
    LogicCell40 \U400_SDRAM.TACK_RNO_1_LC_4_7_1  (
            .in0(N__5149),
            .in1(N__5269),
            .in2(N__2656),
            .in3(N__4741),
            .lcout(\U400_SDRAM.un1_SDRAM_COUNTER52_4_0_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_7_LC_4_7_3 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_7_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_7_LC_4_7_3 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \U400_SDRAM.TACK_RNO_7_LC_4_7_3  (
            .in0(N__4960),
            .in1(N__5078),
            .in2(N__5159),
            .in3(N__4827),
            .lcout(),
            .ltout(\U400_SDRAM.N_208_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_2_LC_4_7_4 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_2_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_2_LC_4_7_4 .LUT_INIT=16'b1111010011111111;
    LogicCell40 \U400_SDRAM.TACK_RNO_2_LC_4_7_4  (
            .in0(N__5080),
            .in1(N__3187),
            .in2(N__2905),
            .in3(N__4712),
            .lcout(\U400_SDRAM.un1_SDRAM_COUNTER52_4_0_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RASn_LC_4_9_2 .C_ON=1'b0;
    defparam \U400_SDRAM.RASn_LC_4_9_2 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.RASn_LC_4_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U400_SDRAM.RASn_LC_4_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6049),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.RASnC_net ),
            .ce(),
            .sr(N__5921));
    defparam \U400_SDRAM.CASn_LC_4_9_6 .C_ON=1'b0;
    defparam \U400_SDRAM.CASn_LC_4_9_6 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.CASn_LC_4_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U400_SDRAM.CASn_LC_4_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6299),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.RASnC_net ),
            .ce(),
            .sr(N__5921));
    defparam \U400_SDRAM.WEn_LC_4_9_7 .C_ON=1'b0;
    defparam \U400_SDRAM.WEn_LC_4_9_7 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.WEn_LC_4_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U400_SDRAM.WEn_LC_4_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6198),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.RASnC_net ),
            .ce(),
            .sr(N__5921));
    defparam \U400_SDRAM.MA_8_LC_4_12_3 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_8_LC_4_12_3 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_8_LC_4_12_3 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \U400_SDRAM.MA_8_LC_4_12_3  (
            .in0(N__2863),
            .in1(N__6113),
            .in2(N__2845),
            .in3(N__6360),
            .lcout(MA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_8C_net ),
            .ce(),
            .sr(N__5924));
    defparam \U400_SDRAM.MA_7_LC_4_12_7 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_7_LC_4_12_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_7_LC_4_12_7 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \U400_SDRAM.MA_7_LC_4_12_7  (
            .in0(N__2818),
            .in1(N__2806),
            .in2(N__6115),
            .in3(N__6359),
            .lcout(MA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_8C_net ),
            .ce(),
            .sr(N__5924));
    defparam \U400_SDRAM.MA_6_LC_4_14_0 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_6_LC_4_14_0 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_6_LC_4_14_0 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \U400_SDRAM.MA_6_LC_4_14_0  (
            .in0(N__2788),
            .in1(N__6109),
            .in2(N__2779),
            .in3(N__6376),
            .lcout(MA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_6C_net ),
            .ce(),
            .sr(N__5932));
    defparam \U400_SDRAM.un2_REFRESH_COUNTER_cry_1_c_LC_5_3_0 .C_ON=1'b1;
    defparam \U400_SDRAM.un2_REFRESH_COUNTER_cry_1_c_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.un2_REFRESH_COUNTER_cry_1_c_LC_5_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U400_SDRAM.un2_REFRESH_COUNTER_cry_1_c_LC_5_3_0  (
            .in0(_gnd_net_),
            .in1(N__3366),
            .in2(N__3277),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_3_0_),
            .carryout(\U400_SDRAM.un2_REFRESH_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_2_LC_5_3_1 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_2_LC_5_3_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_2_LC_5_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_2_LC_5_3_1  (
            .in0(_gnd_net_),
            .in1(N__3394),
            .in2(_gnd_net_),
            .in3(N__2983),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U400_SDRAM.un2_REFRESH_COUNTER_cry_1 ),
            .carryout(\U400_SDRAM.un2_REFRESH_COUNTER_cry_2 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3424));
    defparam \U400_SDRAM.REFRESH_COUNTER_3_LC_5_3_2 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_3_LC_5_3_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_3_LC_5_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_3_LC_5_3_2  (
            .in0(_gnd_net_),
            .in1(N__3408),
            .in2(_gnd_net_),
            .in3(N__2980),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U400_SDRAM.un2_REFRESH_COUNTER_cry_2 ),
            .carryout(\U400_SDRAM.un2_REFRESH_COUNTER_cry_3 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3424));
    defparam \U400_SDRAM.REFRESH_COUNTER_4_LC_5_3_3 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_4_LC_5_3_3 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_4_LC_5_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_4_LC_5_3_3  (
            .in0(_gnd_net_),
            .in1(N__3381),
            .in2(_gnd_net_),
            .in3(N__2977),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U400_SDRAM.un2_REFRESH_COUNTER_cry_3 ),
            .carryout(\U400_SDRAM.un2_REFRESH_COUNTER_cry_4 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3424));
    defparam \U400_SDRAM.REFRESH_COUNTER_5_LC_5_3_4 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_5_LC_5_3_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_5_LC_5_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_5_LC_5_3_4  (
            .in0(_gnd_net_),
            .in1(N__3238),
            .in2(_gnd_net_),
            .in3(N__2974),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U400_SDRAM.un2_REFRESH_COUNTER_cry_4 ),
            .carryout(\U400_SDRAM.un2_REFRESH_COUNTER_cry_5 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3424));
    defparam \U400_SDRAM.REFRESH_COUNTER_6_LC_5_3_5 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_6_LC_5_3_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_6_LC_5_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_6_LC_5_3_5  (
            .in0(_gnd_net_),
            .in1(N__3289),
            .in2(_gnd_net_),
            .in3(N__2971),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U400_SDRAM.un2_REFRESH_COUNTER_cry_5 ),
            .carryout(\U400_SDRAM.un2_REFRESH_COUNTER_cry_6 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3424));
    defparam \U400_SDRAM.REFRESH_COUNTER_7_LC_5_3_6 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_7_LC_5_3_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_7_LC_5_3_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_7_LC_5_3_6  (
            .in0(_gnd_net_),
            .in1(N__3252),
            .in2(_gnd_net_),
            .in3(N__2968),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(\U400_SDRAM.un2_REFRESH_COUNTER_cry_6 ),
            .carryout(\U400_SDRAM.un2_REFRESH_COUNTER_cry_7 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3424));
    defparam \U400_SDRAM.REFRESH_COUNTER_8_LC_5_3_7 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_8_LC_5_3_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_8_LC_5_3_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_8_LC_5_3_7  (
            .in0(_gnd_net_),
            .in1(N__3207),
            .in2(_gnd_net_),
            .in3(N__2965),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3424));
    defparam \U400_SDRAM.TA_OUT_LC_5_4_2 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_OUT_LC_5_4_2 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.TA_OUT_LC_5_4_2 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \U400_SDRAM.TA_OUT_LC_5_4_2  (
            .in0(N__2961),
            .in1(N__2932),
            .in2(N__2922),
            .in3(N__3295),
            .lcout(TA_OUT),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3639),
            .ce(),
            .sr(N__5927));
    defparam \U400_SDRAM.BURST_RNISKH51_LC_5_5_0 .C_ON=1'b0;
    defparam \U400_SDRAM.BURST_RNISKH51_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.BURST_RNISKH51_LC_5_5_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U400_SDRAM.BURST_RNISKH51_LC_5_5_0  (
            .in0(N__3081),
            .in1(N__3343),
            .in2(N__3053),
            .in3(N__3308),
            .lcout(\U400_SDRAM.TA_COUNTER_0_sqmuxa ),
            .ltout(\U400_SDRAM.TA_COUNTER_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_EN_i_ess_RNO_1_LC_5_5_1 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_EN_i_ess_RNO_1_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_EN_i_ess_RNO_1_LC_5_5_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \U400_SDRAM.TA_EN_i_ess_RNO_1_LC_5_5_1  (
            .in0(N__3714),
            .in1(N__3009),
            .in2(N__2998),
            .in3(N__3675),
            .lcout(\U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.BURST_LC_5_5_3 .C_ON=1'b0;
    defparam \U400_SDRAM.BURST_LC_5_5_3 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.BURST_LC_5_5_3 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \U400_SDRAM.BURST_LC_5_5_3  (
            .in0(N__3309),
            .in1(N__5751),
            .in2(N__5686),
            .in3(N__3154),
            .lcout(\U400_SDRAM.BURSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.BURSTC_net ),
            .ce(),
            .sr(N__5925));
    defparam \U400_SDRAM.RAM_CYCLE_RNO_1_LC_5_6_0 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_1_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_1_LC_5_6_0 .LUT_INIT=16'b1011111111001111;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_RNO_1_LC_5_6_0  (
            .in0(N__4963),
            .in1(N__5272),
            .in2(N__4709),
            .in3(N__5077),
            .lcout(),
            .ltout(\U400_SDRAM.un1_SDRAM_COUNTER52_2_0_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_RNO_0_LC_5_6_1 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_0_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_0_LC_5_6_1 .LUT_INIT=16'b0000111000001100;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_RNO_0_LC_5_6_1  (
            .in0(N__4015),
            .in1(N__3444),
            .in2(N__2995),
            .in3(N__3950),
            .lcout(\U400_SDRAM.RAM_CYCLE_e_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNISAQQ4_LC_5_6_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNISAQQ4_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNISAQQ4_LC_5_6_2 .LUT_INIT=16'b1111111100111111;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNISAQQ4_LC_5_6_2  (
            .in0(_gnd_net_),
            .in1(N__4014),
            .in2(N__4711),
            .in3(N__4067),
            .lcout(\U400_SDRAM.N_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_5_LC_5_6_3 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_5_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_5_LC_5_6_3 .LUT_INIT=16'b1111111100110001;
    LogicCell40 \U400_SDRAM.TACK_RNO_5_LC_5_6_3  (
            .in0(N__5271),
            .in1(N__3443),
            .in2(N__5152),
            .in3(N__4867),
            .lcout(\U400_SDRAM.TACK_7_iv_i_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_RNI58I35_LC_5_6_4 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNI58I35_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNI58I35_LC_5_6_4 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_RNI58I35_LC_5_6_4  (
            .in0(N__3951),
            .in1(N__4066),
            .in2(N__4710),
            .in3(N__4013),
            .lcout(\U400_SDRAM.N_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.WRITE_CYCLE_RNI18LH_LC_5_6_5 .C_ON=1'b0;
    defparam \U400_SDRAM.WRITE_CYCLE_RNI18LH_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.WRITE_CYCLE_RNI18LH_LC_5_6_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U400_SDRAM.WRITE_CYCLE_RNI18LH_LC_5_6_5  (
            .in0(N__5270),
            .in1(N__5127),
            .in2(_gnd_net_),
            .in3(N__4961),
            .lcout(\U400_SDRAM.N_255 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_4_LC_5_6_6 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_4_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_4_LC_5_6_6 .LUT_INIT=16'b1110110011011100;
    LogicCell40 \U400_SDRAM.TACK_RNO_4_LC_5_6_6  (
            .in0(N__4962),
            .in1(N__4159),
            .in2(N__5150),
            .in3(N__5273),
            .lcout(),
            .ltout(\U400_SDRAM.TACK_7_iv_i_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_0_LC_5_6_7 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_0_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_0_LC_5_6_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U400_SDRAM.TACK_RNO_0_LC_5_6_7  (
            .in0(N__3186),
            .in1(N__3460),
            .in2(N__3175),
            .in3(N__3172),
            .lcout(\U400_SDRAM.N_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_LC_5_7_1 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_LC_5_7_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.RAM_CYCLE_LC_5_7_1 .LUT_INIT=16'b1111000001110010;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_LC_5_7_1  (
            .in0(N__3160),
            .in1(N__3152),
            .in2(N__3550),
            .in3(N__4441),
            .lcout(\U400_SDRAM.RAM_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.RAM_CYCLEC_net ),
            .ce(),
            .sr(N__5923));
    defparam \U400_SDRAM.WRITE_CYCLE_LC_5_7_2 .C_ON=1'b0;
    defparam \U400_SDRAM.WRITE_CYCLE_LC_5_7_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.WRITE_CYCLE_LC_5_7_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \U400_SDRAM.WRITE_CYCLE_LC_5_7_2  (
            .in0(N__3153),
            .in1(N__3139),
            .in2(_gnd_net_),
            .in3(N__5142),
            .lcout(\U400_SDRAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.RAM_CYCLEC_net ),
            .ce(),
            .sr(N__5923));
    defparam \U400_SDRAM.CS0_EN_LC_5_8_0 .C_ON=1'b0;
    defparam \U400_SDRAM.CS0_EN_LC_5_8_0 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.CS0_EN_LC_5_8_0 .LUT_INIT=16'b1111111100010011;
    LogicCell40 \U400_SDRAM.CS0_EN_LC_5_8_0  (
            .in0(N__4029),
            .in1(N__4073),
            .in2(N__4713),
            .in3(N__3481),
            .lcout(\U400_SDRAM.CS0_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS0_ENC_net ),
            .ce(),
            .sr(N__5920));
    defparam \U400_SDRAM.CS0n_LC_5_8_1 .C_ON=1'b0;
    defparam \U400_SDRAM.CS0n_LC_5_8_1 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.CS0n_LC_5_8_1 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \U400_SDRAM.CS0n_LC_5_8_1  (
            .in0(N__6297),
            .in1(N__6055),
            .in2(N__3505),
            .in3(N__6188),
            .lcout(CS0n_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS0_ENC_net ),
            .ce(),
            .sr(N__5920));
    defparam \U400_SDRAM.MA_9_LC_5_8_2 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_9_LC_5_8_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_9_LC_5_8_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U400_SDRAM.MA_9_LC_5_8_2  (
            .in0(N__6189),
            .in1(N__6056),
            .in2(N__3109),
            .in3(N__6298),
            .lcout(MA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS0_ENC_net ),
            .ce(),
            .sr(N__5920));
    defparam \U400_SDRAM.CS1_EN_LC_5_8_7 .C_ON=1'b0;
    defparam \U400_SDRAM.CS1_EN_LC_5_8_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.CS1_EN_LC_5_8_7 .LUT_INIT=16'b1111111100010101;
    LogicCell40 \U400_SDRAM.CS1_EN_LC_5_8_7  (
            .in0(N__4074),
            .in1(N__4030),
            .in2(N__4714),
            .in3(N__3532),
            .lcout(\U400_SDRAM.CS1_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS0_ENC_net ),
            .ce(),
            .sr(N__5920));
    defparam \U400_SDRAM.REFRESH_COUNTER_0_LC_6_3_1 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_0_LC_6_3_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_0_LC_6_3_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_0_LC_6_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3275),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_0C_net ),
            .ce(),
            .sr(N__3423));
    defparam \U400_SDRAM.REFRESH_COUNTER_1_LC_6_3_2 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_1_LC_6_3_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_1_LC_6_3_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_1_LC_6_3_2  (
            .in0(N__3276),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3367),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_0C_net ),
            .ce(),
            .sr(N__3423));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2_1_LC_6_4_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2_1_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2_1_LC_6_4_0 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2_1_LC_6_4_0  (
            .in0(N__5556),
            .in1(N__5276),
            .in2(_gnd_net_),
            .in3(N__3475),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_RNIJKCA2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIMIPA1_1_LC_6_4_1 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIMIPA1_1_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIMIPA1_1_LC_6_4_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_RNIMIPA1_1_LC_6_4_1  (
            .in0(N__3409),
            .in1(N__3393),
            .in2(N__3382),
            .in3(N__3365),
            .lcout(\U400_SDRAM.un1_REFRESH_COUNTERlto7_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_OUT_RNO_0_LC_6_4_3 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_OUT_RNO_0_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_OUT_RNO_0_LC_6_4_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U400_SDRAM.TA_OUT_RNO_0_LC_6_4_3  (
            .in0(_gnd_net_),
            .in1(N__3349),
            .in2(_gnd_net_),
            .in3(N__3310),
            .lcout(\U400_SDRAM.TA_EN11_m ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIUQPA1_5_LC_6_4_4 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIUQPA1_5_LC_6_4_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIUQPA1_5_LC_6_4_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_RNIUQPA1_5_LC_6_4_4  (
            .in0(N__3288),
            .in1(N__3271),
            .in2(N__3253),
            .in3(N__3237),
            .lcout(\U400_SDRAM.un1_REFRESH_COUNTERlto7_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_6_5_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_6_5_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_6_5_0  (
            .in0(N__3846),
            .in1(N__4016),
            .in2(_gnd_net_),
            .in3(N__4825),
            .lcout(),
            .ltout(\U400_SDRAM.N_205_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_1_LC_6_5_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_1_LC_6_5_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CMD_1_LC_6_5_1 .LUT_INIT=16'b1000100010001011;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_1_LC_6_5_1  (
            .in0(N__6255),
            .in1(N__3874),
            .in2(N__3226),
            .in3(N__3853),
            .lcout(\U400_SDRAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_CMD_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_EN_i_ess_RNO_0_LC_6_5_4 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_EN_i_ess_RNO_0_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_EN_i_ess_RNO_0_LC_6_5_4 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U400_SDRAM.TA_EN_i_ess_RNO_0_LC_6_5_4  (
            .in0(N__5941),
            .in1(_gnd_net_),
            .in2(N__3223),
            .in3(_gnd_net_),
            .lcout(\U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIVV903_8_LC_6_5_5 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIVV903_8_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIVV903_8_LC_6_5_5 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_RNIVV903_8_LC_6_5_5  (
            .in0(N__3214),
            .in1(N__3208),
            .in2(_gnd_net_),
            .in3(N__3193),
            .lcout(\U400_SDRAM.REFRESH_COUNTER_RNIVV903Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_6_6_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_6_6_0 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_6_6_0  (
            .in0(N__4012),
            .in1(N__4577),
            .in2(N__3448),
            .in3(N__3949),
            .lcout(\U400_SDRAM.N_199 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_3_LC_6_6_1 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_3_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_3_LC_6_6_1 .LUT_INIT=16'b0000000010001100;
    LogicCell40 \U400_SDRAM.TACK_RNO_3_LC_6_6_1  (
            .in0(N__5274),
            .in1(N__5076),
            .in2(N__4828),
            .in3(N__5131),
            .lcout(\U400_SDRAM.N_189 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_0_LC_6_6_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_0_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_0_LC_6_6_4 .LUT_INIT=16'b0011011101110111;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_2_0_LC_6_6_4  (
            .in0(N__4824),
            .in1(N__3845),
            .in2(N__5151),
            .in3(N__4947),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_0_1_32_i_0_i_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_0_LC_6_6_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_0_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_0_LC_6_6_5 .LUT_INIT=16'b0010111100001111;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_1_0_LC_6_6_5  (
            .in0(N__5275),
            .in1(N__4581),
            .in2(N__3454),
            .in3(N__5135),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_0_1_32_i_0_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_0_LC_6_6_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_0_LC_6_6_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CMD_0_LC_6_6_6 .LUT_INIT=16'b1000100010001011;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_0_LC_6_6_6  (
            .in0(N__6161),
            .in1(N__3869),
            .in2(N__3451),
            .in3(N__3430),
            .lcout(\U400_SDRAM.SDRAM_CMDZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_CMD_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIP3PD_0_LC_6_7_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIP3PD_0_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIP3PD_0_LC_6_7_0 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIP3PD_0_LC_6_7_0  (
            .in0(N__4939),
            .in1(_gnd_net_),
            .in2(N__5075),
            .in3(_gnd_net_),
            .lcout(\U400_SDRAM.N_128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNITTDH4_0_LC_6_7_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNITTDH4_0_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNITTDH4_0_LC_6_7_1 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNITTDH4_0_LC_6_7_1  (
            .in0(N__5541),
            .in1(N__3820),
            .in2(_gnd_net_),
            .in3(N__4242),
            .lcout(\U400_SDRAM.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_0_LC_6_7_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_0_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_0_LC_6_7_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_0_LC_6_7_4  (
            .in0(N__4938),
            .in1(N__5242),
            .in2(N__5074),
            .in3(N__4433),
            .lcout(\U400_SDRAM.N_139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_0_LC_6_7_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_0_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_0_LC_6_7_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_0_0_LC_6_7_5  (
            .in0(_gnd_net_),
            .in1(N__4147),
            .in2(_gnd_net_),
            .in3(N__4093),
            .lcout(\U400_SDRAM.N_185 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_LC_6_7_6 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_LC_6_7_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.RAM_CYCLE_START_LC_6_7_6 .LUT_INIT=16'b1011000010100000;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_LC_6_7_6  (
            .in0(N__5764),
            .in1(N__3546),
            .in2(N__5554),
            .in3(N__3958),
            .lcout(\U400_SDRAM.RAM_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3631),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIPOT15_LC_6_8_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIPOT15_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIPOT15_LC_6_8_1 .LUT_INIT=16'b0011101111111011;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNIPOT15_LC_6_8_1  (
            .in0(N__4240),
            .in1(N__4065),
            .in2(N__4707),
            .in3(N__4092),
            .lcout(\U400_SDRAM.N_75 ),
            .ltout(\U400_SDRAM.N_75_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.CS1_EN_RNO_0_LC_6_8_2 .C_ON=1'b0;
    defparam \U400_SDRAM.CS1_EN_RNO_0_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.CS1_EN_RNO_0_LC_6_8_2 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \U400_SDRAM.CS1_EN_RNO_0_LC_6_8_2  (
            .in0(N__3517),
            .in1(N__3804),
            .in2(N__3535),
            .in3(N__3523),
            .lcout(\U400_SDRAM.CS1_EN_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIHALH3_LC_6_8_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIHALH3_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIHALH3_LC_6_8_4 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNIHALH3_LC_6_8_4  (
            .in0(N__4091),
            .in1(N__4680),
            .in2(N__5281),
            .in3(N__4239),
            .lcout(),
            .ltout(\U400_SDRAM.CS1_EN_7_i_0_o3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIA1BE8_LC_6_8_5 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIA1BE8_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIA1BE8_LC_6_8_5 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_RNIA1BE8_LC_6_8_5  (
            .in0(N__4019),
            .in1(N__3471),
            .in2(N__3526),
            .in3(N__3948),
            .lcout(\U400_SDRAM.N_159 ),
            .ltout(\U400_SDRAM.N_159_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.CS0_EN_RNO_0_LC_6_8_6 .C_ON=1'b0;
    defparam \U400_SDRAM.CS0_EN_RNO_0_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.CS0_EN_RNO_0_LC_6_8_6 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \U400_SDRAM.CS0_EN_RNO_0_LC_6_8_6  (
            .in0(N__3516),
            .in1(N__3501),
            .in2(N__3490),
            .in3(N__3487),
            .lcout(\U400_SDRAM.CS0_EN_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIHPJJ1_LC_6_8_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIHPJJ1_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIHPJJ1_LC_6_8_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNIHPJJ1_LC_6_8_7  (
            .in0(N__5039),
            .in1(N__4940),
            .in2(N__4706),
            .in3(N__4434),
            .lcout(\U400_SDRAM.N_250 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_6_9_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_6_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_6_9_1  (
            .in0(N__5043),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3744),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_6_9_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_6_9_6 .LUT_INIT=16'b0110001000100010;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_6_9_6  (
            .in0(N__5280),
            .in1(N__5042),
            .in2(N__5160),
            .in3(N__4826),
            .lcout(),
            .ltout(\U400_SDRAM.N_176_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_6_9_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_6_9_7 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_6_9_7  (
            .in0(N__4640),
            .in1(N__4862),
            .in2(N__3814),
            .in3(N__4099),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.CS1n_LC_6_10_2 .C_ON=1'b0;
    defparam \U400_SDRAM.CS1n_LC_6_10_2 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.CS1n_LC_6_10_2 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \U400_SDRAM.CS1n_LC_6_10_2  (
            .in0(N__6047),
            .in1(N__6190),
            .in2(N__3811),
            .in3(N__6301),
            .lcout(CS1n_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS1nC_net ),
            .ce(),
            .sr(N__5926));
    defparam \U400_SDRAM.MA_12_LC_6_10_6 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_12_LC_6_10_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_12_LC_6_10_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U400_SDRAM.MA_12_LC_6_10_6  (
            .in0(N__6048),
            .in1(N__6191),
            .in2(N__3784),
            .in3(N__6302),
            .lcout(MA_c_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS1nC_net ),
            .ce(),
            .sr(N__5926));
    defparam \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_6_12_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_6_12_2 .LUT_INIT=16'b1011101101010101;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_6_12_2  (
            .in0(N__6042),
            .in1(N__6162),
            .in2(_gnd_net_),
            .in3(N__6256),
            .lcout(\U400_SDRAM.MAc_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_6_12_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_6_12_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_6_12_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_6_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_BYTE_ENABLE.un1_UUBEn_0_a3_LC_7_3_6 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_UUBEn_0_a3_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_UUBEn_0_a3_LC_7_3_6 .LUT_INIT=16'b0000111011100000;
    LogicCell40 \U400_BYTE_ENABLE.un1_UUBEn_0_a3_LC_7_3_6  (
            .in0(N__5841),
            .in1(N__5812),
            .in2(N__5752),
            .in3(N__5685),
            .lcout(UUBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_EN_i_ess_LC_7_5_5 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_EN_i_ess_LC_7_5_5 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.TA_EN_i_ess_LC_7_5_5 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U400_SDRAM.TA_EN_i_ess_LC_7_5_5  (
            .in0(N__5523),
            .in1(N__3718),
            .in2(_gnd_net_),
            .in3(N__3691),
            .lcout(TA_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3644),
            .ce(N__3562),
            .sr(N__5933));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7J_0_LC_7_6_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7J_0_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7J_0_LC_7_6_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7J_0_LC_7_6_0  (
            .in0(N__5527),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4684),
            .lcout(\U400_SDRAM.N_252 ),
            .ltout(\U400_SDRAM.N_252_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_7_6_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_7_6_1 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_7_6_1  (
            .in0(N__5241),
            .in1(N__4405),
            .in2(N__3553),
            .in3(N__4948),
            .lcout(),
            .ltout(\U400_SDRAM.N_200_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_7_6_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_7_6_2 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_7_6_2  (
            .in0(N__4132),
            .in1(N__3847),
            .in2(N__3889),
            .in3(N__4805),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_0_61_i_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_2_LC_7_6_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_2_LC_7_6_3 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CMD_2_LC_7_6_3 .LUT_INIT=16'b1010101000000011;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_2_LC_7_6_3  (
            .in0(N__6029),
            .in1(N__3886),
            .in2(N__3877),
            .in3(N__3873),
            .lcout(\U400_SDRAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_CMD_2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_7_6_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_7_6_4 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_7_6_4  (
            .in0(N__4131),
            .in1(N__5240),
            .in2(N__4582),
            .in3(N__3826),
            .lcout(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIA54Q_LC_7_6_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIA54Q_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIA54Q_LC_7_6_7 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNIA54Q_LC_7_6_7  (
            .in0(N__5073),
            .in1(_gnd_net_),
            .in2(N__4708),
            .in3(N__5526),
            .lcout(\U400_SDRAM.N_228 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_LC_7_7_0 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_LC_7_7_0 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_LC_7_7_0  (
            .in0(N__4565),
            .in1(N__3944),
            .in2(N__4075),
            .in3(N__4017),
            .lcout(\U400_SDRAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_0_LC_7_7_1 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_0_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_0_LC_7_7_1 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_0_LC_7_7_1  (
            .in0(N__4018),
            .in1(N__4069),
            .in2(N__3959),
            .in3(N__4566),
            .lcout(\U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5Z0Z_0 ),
            .ltout(\U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_3_LC_7_7_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_3_LC_7_7_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_3_LC_7_7_2 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_3_LC_7_7_2  (
            .in0(N__5617),
            .in1(N__4372),
            .in2(N__3829),
            .in3(N__4314),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_3C_net ),
            .ce(N__5315),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_7_7_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_7_7_7 .LUT_INIT=16'b0110000000000000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_7_7_7  (
            .in0(N__5236),
            .in1(N__4946),
            .in2(N__5553),
            .in3(N__4400),
            .lcout(\U400_SDRAM.N_203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2_0_LC_7_8_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2_0_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2_0_LC_7_8_0 .LUT_INIT=16'b0000101000001110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2_0_LC_7_8_0  (
            .in0(N__4734),
            .in1(N__5232),
            .in2(N__4576),
            .in3(N__5041),
            .lcout(\U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_7_8_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_7_8_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_7_8_1  (
            .in0(N__4332),
            .in1(N__4347),
            .in2(N__5335),
            .in3(N__4362),
            .lcout(\U400_SDRAM.N_126 ),
            .ltout(\U400_SDRAM.N_126_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIFAF21_2_LC_7_8_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIFAF21_2_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIFAF21_2_LC_7_8_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIFAF21_2_LC_7_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4108),
            .in3(N__4778),
            .lcout(\U400_SDRAM.N_129 ),
            .ltout(\U400_SDRAM.N_129_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_0_0_LC_7_8_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_0_0_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_0_0_LC_7_8_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_0_0_LC_7_8_3  (
            .in0(N__4927),
            .in1(N__5225),
            .in2(N__4105),
            .in3(N__5021),
            .lcout(\U400_SDRAM.N_257 ),
            .ltout(\U400_SDRAM.N_257_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_5_0_LC_7_8_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_5_0_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_5_0_LC_7_8_4 .LUT_INIT=16'b1111110111110101;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_5_0_LC_7_8_4  (
            .in0(N__5525),
            .in1(N__4660),
            .in2(N__4102),
            .in3(N__4928),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_0_LC_7_8_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_0_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_0_LC_7_8_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_0_LC_7_8_5  (
            .in0(N__4926),
            .in1(N__5022),
            .in2(_gnd_net_),
            .in3(N__4431),
            .lcout(\U400_SDRAM.N_133 ),
            .ltout(\U400_SDRAM.N_133_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3_LC_7_8_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3_LC_7_8_6 .LUT_INIT=16'b0011111100001100;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3_LC_7_8_6  (
            .in0(_gnd_net_),
            .in1(N__4659),
            .in2(N__4078),
            .in3(N__4241),
            .lcout(),
            .ltout(\U400_SDRAM.N_141_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIJG6G7_LC_7_8_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIJG6G7_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIJG6G7_LC_7_8_7 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNIJG6G7_LC_7_8_7  (
            .in0(N__4068),
            .in1(N__5524),
            .in2(N__4033),
            .in3(N__4969),
            .lcout(\U400_SDRAM.N_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_7_9_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_7_9_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_7_9_6  (
            .in0(N__4028),
            .in1(N__4404),
            .in2(N__4723),
            .in3(N__3965),
            .lcout(),
            .ltout(\U400_SDRAM.N_181_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_0_LC_7_9_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_0_LC_7_9_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_0_LC_7_9_7 .LUT_INIT=16'b0000010111001100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_0_LC_7_9_7  (
            .in0(N__3904),
            .in1(N__3898),
            .in2(N__3892),
            .in3(N__4306),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_0C_net ),
            .ce(N__5319),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_11_LC_7_10_4 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_11_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_11_LC_7_10_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U400_SDRAM.MA_11_LC_7_10_4  (
            .in0(N__6046),
            .in1(N__6203),
            .in2(N__4273),
            .in3(N__6300),
            .lcout(MA_c_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_11C_net ),
            .ce(),
            .sr(N__5928));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_LC_7_10_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_LC_7_10_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_LC_7_10_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_LC_7_10_5  (
            .in0(_gnd_net_),
            .in1(N__4641),
            .in2(_gnd_net_),
            .in3(N__4246),
            .lcout(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_11C_net ),
            .ce(),
            .sr(N__5928));
    defparam \U400_SDRAM.MA_4_LC_7_16_3 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_4_LC_7_16_3 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_4_LC_7_16_3 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \U400_SDRAM.MA_4_LC_7_16_3  (
            .in0(N__4216),
            .in1(N__6090),
            .in2(N__4201),
            .in3(N__6384),
            .lcout(MA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_4C_net ),
            .ce(),
            .sr(N__5935));
    defparam \U400_SDRAM.MA_5_LC_7_16_4 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_5_LC_7_16_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_5_LC_7_16_4 .LUT_INIT=16'b0000001000110001;
    LogicCell40 \U400_SDRAM.MA_5_LC_7_16_4  (
            .in0(N__6204),
            .in1(N__4501),
            .in2(N__6108),
            .in3(N__6318),
            .lcout(MA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_4C_net ),
            .ce(),
            .sr(N__5935));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI6MLK_2_LC_8_6_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI6MLK_2_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI6MLK_2_LC_8_6_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI6MLK_2_LC_8_6_3  (
            .in0(N__5072),
            .in1(N__4929),
            .in2(_gnd_net_),
            .in3(N__4803),
            .lcout(\U400_SDRAM.N_150 ),
            .ltout(\U400_SDRAM.N_150_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIVPE21_2_LC_8_6_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIVPE21_2_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIVPE21_2_LC_8_6_4 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIVPE21_2_LC_8_6_4  (
            .in0(N__4804),
            .in1(_gnd_net_),
            .in2(N__4150),
            .in3(N__5268),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_0_61_i_i_a3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI079H2_2_LC_8_6_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI079H2_2_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI079H2_2_LC_8_6_5 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI079H2_2_LC_8_6_5  (
            .in0(_gnd_net_),
            .in1(N__4146),
            .in2(N__4135),
            .in3(N__4866),
            .lcout(\U400_SDRAM.N_201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TAn_obuft_RNO_LC_8_6_6.C_ON=1'b0;
    defparam TAn_obuft_RNO_LC_8_6_6.SEQ_MODE=4'b0000;
    defparam TAn_obuft_RNO_LC_8_6_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 TAn_obuft_RNO_LC_8_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4123),
            .lcout(N_529_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_1_LC_8_7_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_1_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_1_LC_8_7_5 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_1_LC_8_7_5  (
            .in0(N__4384),
            .in1(N__4447),
            .in2(N__5613),
            .in3(N__4315),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_1C_net ),
            .ce(N__5314),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIQQB91_0_LC_8_8_0 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIQQB91_0_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIQQB91_0_LC_8_8_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIQQB91_0_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__5040),
            .in2(_gnd_net_),
            .in3(N__4432),
            .lcout(\U400_SDRAM.N_260 ),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_8_8_1 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_8_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__5267),
            .in2(_gnd_net_),
            .in3(N__4378),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_s_1 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_2_LC_8_8_2 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_2_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_2_LC_8_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_2_LC_8_8_2  (
            .in0(N__4316),
            .in1(N__4802),
            .in2(_gnd_net_),
            .in3(N__4375),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_2 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__5320),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_8_8_3 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_8_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(N__4949),
            .in2(_gnd_net_),
            .in3(N__4366),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_s_3 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_4_LC_8_8_4 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_4_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_4_LC_8_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_4_LC_8_8_4  (
            .in0(N__4317),
            .in1(N__4363),
            .in2(_gnd_net_),
            .in3(N__4351),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_4 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__5320),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_5_LC_8_8_5 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_5_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_5_LC_8_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_5_LC_8_8_5  (
            .in0(N__4304),
            .in1(N__4348),
            .in2(_gnd_net_),
            .in3(N__4336),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_5 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__5320),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_6_LC_8_8_6 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_6_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_6_LC_8_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_6_LC_8_8_6  (
            .in0(N__4318),
            .in1(N__4333),
            .in2(_gnd_net_),
            .in3(N__4321),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_6 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__5320),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_7_LC_8_8_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_7_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_7_LC_8_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_7_LC_8_8_7  (
            .in0(N__4305),
            .in1(N__5334),
            .in2(_gnd_net_),
            .in3(N__4276),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__5320),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.WRITE_CYCLE_RNICOHO_LC_8_9_0 .C_ON=1'b0;
    defparam \U400_SDRAM.WRITE_CYCLE_RNICOHO_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.WRITE_CYCLE_RNICOHO_LC_8_9_0 .LUT_INIT=16'b0111011001100110;
    LogicCell40 \U400_SDRAM.WRITE_CYCLE_RNICOHO_LC_8_9_0  (
            .in0(N__4951),
            .in1(N__5266),
            .in2(N__5161),
            .in3(N__5038),
            .lcout(),
            .ltout(\U400_SDRAM.N_161_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI4ECU1_2_LC_8_9_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI4ECU1_2_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI4ECU1_2_LC_8_9_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI4ECU1_2_LC_8_9_1  (
            .in0(N__4780),
            .in1(N__4628),
            .in2(N__4972),
            .in3(N__4855),
            .lcout(\U400_SDRAM.N_183 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNITTB91_2_LC_8_9_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNITTB91_2_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNITTB91_2_LC_8_9_2 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNITTB91_2_LC_8_9_2  (
            .in0(N__4950),
            .in1(N__4854),
            .in2(_gnd_net_),
            .in3(N__4779),
            .lcout(\U400_SDRAM.N_138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_8_9_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_8_9_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_8_9_6  (
            .in0(N__4629),
            .in1(N__5741),
            .in2(_gnd_net_),
            .in3(N__5675),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_a3_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7J_LC_8_10_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7J_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7J_LC_8_10_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7J_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__5488),
            .in2(_gnd_net_),
            .in3(N__4627),
            .lcout(\U400_SDRAM.SDRAM_CONFIGURED_RNIVK7JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_RNO_0_5_LC_8_15_7 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_RNO_0_5_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.MA_RNO_0_5_LC_8_15_7 .LUT_INIT=16'b0100111101000100;
    LogicCell40 \U400_SDRAM.MA_RNO_0_5_LC_8_15_7  (
            .in0(N__4528),
            .in1(N__6087),
            .in2(N__4516),
            .in3(N__6303),
            .lcout(\U400_SDRAM.MAc_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_0_LC_8_16_1 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_0_LC_8_16_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_0_LC_8_16_1 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \U400_SDRAM.MA_0_LC_8_16_1  (
            .in0(N__4495),
            .in1(N__6089),
            .in2(N__4483),
            .in3(N__6385),
            .lcout(MA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_0C_net ),
            .ce(),
            .sr(N__5936));
    defparam \U400_SDRAM.MA_10_LC_8_16_2 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_10_LC_8_16_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_10_LC_8_16_2 .LUT_INIT=16'b0101101000011010;
    LogicCell40 \U400_SDRAM.MA_10_LC_8_16_2  (
            .in0(N__6088),
            .in1(N__6199),
            .in2(N__6319),
            .in3(N__4462),
            .lcout(MA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_0C_net ),
            .ce(),
            .sr(N__5936));
    defparam \U400_BYTE_ENABLE.un1_UMBEn_0_LC_9_3_0 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_UMBEn_0_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_UMBEn_0_LC_9_3_0 .LUT_INIT=16'b0110000001100100;
    LogicCell40 \U400_BYTE_ENABLE.un1_UMBEn_0_LC_9_3_0  (
            .in0(N__5744),
            .in1(N__5681),
            .in2(N__5857),
            .in3(N__5817),
            .lcout(UMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_BYTE_ENABLE.un1_LLBEn_0_LC_9_3_1 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_LLBEn_0_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_LLBEn_0_LC_9_3_1 .LUT_INIT=16'b0001000100101010;
    LogicCell40 \U400_BYTE_ENABLE.un1_LLBEn_0_LC_9_3_1  (
            .in0(N__5679),
            .in1(N__5849),
            .in2(N__5818),
            .in3(N__5742),
            .lcout(LLBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_BYTE_ENABLE.un1_LMBEn_0_a3_LC_9_3_4 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_LMBEn_0_a3_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_LMBEn_0_a3_LC_9_3_4 .LUT_INIT=16'b0110011000000110;
    LogicCell40 \U400_BYTE_ENABLE.un1_LMBEn_0_a3_LC_9_3_4  (
            .in0(N__5743),
            .in1(N__5680),
            .in2(N__5856),
            .in3(N__5816),
            .lcout(LMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_9_6_0 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_9_6_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_9_6_0  (
            .in0(N__5490),
            .in1(N__5596),
            .in2(N__5575),
            .in3(N__5776),
            .lcout(\U400_SDRAM.N_220 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.BURST8_0_a2_LC_9_6_2 .C_ON=1'b0;
    defparam \U400_SDRAM.BURST8_0_a2_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.BURST8_0_a2_LC_9_6_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U400_SDRAM.BURST8_0_a2_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(N__5724),
            .in2(_gnd_net_),
            .in3(N__5664),
            .lcout(\U400_SDRAM.BURST8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.N_220_3_i_LC_9_6_5 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.N_220_3_i_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.N_220_3_i_LC_9_6_5 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \U400_ADDRESS_DECODE.N_220_3_i_LC_9_6_5  (
            .in0(N__5595),
            .in1(N__5571),
            .in2(_gnd_net_),
            .in3(N__5489),
            .lcout(N_220_3_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_3_LC_9_13_4 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_3_LC_9_13_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_3_LC_9_13_4 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \U400_SDRAM.MA_3_LC_9_13_4  (
            .in0(N__5395),
            .in1(N__6078),
            .in2(N__5386),
            .in3(N__6375),
            .lcout(MA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_3C_net ),
            .ce(),
            .sr(N__5934));
    defparam \U400_SDRAM.MA_RNO_0_1_LC_9_15_4 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_RNO_0_1_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.MA_RNO_0_1_LC_9_15_4 .LUT_INIT=16'b0100111101000100;
    LogicCell40 \U400_SDRAM.MA_RNO_0_1_LC_9_15_4  (
            .in0(N__5359),
            .in1(N__6103),
            .in2(N__5347),
            .in3(N__6304),
            .lcout(\U400_SDRAM.MAc_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_2_LC_9_16_2 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_2_LC_9_16_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_2_LC_9_16_2 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \U400_SDRAM.MA_2_LC_9_16_2  (
            .in0(N__6104),
            .in1(N__6409),
            .in2(N__6394),
            .in3(N__6383),
            .lcout(MA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_2C_net ),
            .ce(),
            .sr(N__5937));
    defparam \U400_SDRAM.MA_1_LC_9_16_4 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_1_LC_9_16_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_1_LC_9_16_4 .LUT_INIT=16'b0000000001011001;
    LogicCell40 \U400_SDRAM.MA_1_LC_9_16_4  (
            .in0(N__6314),
            .in1(N__6208),
            .in2(N__6114),
            .in3(N__5953),
            .lcout(MA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_2C_net ),
            .ce(),
            .sr(N__5937));
endmodule // U400_TOP

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 12 2025 17:26:36

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U400_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U400_TOP
entity U400_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    MA : out std_logic_vector(12 downto 0);
    A : in std_logic_vector(31 downto 0);
    LBENn : out std_logic;
    CS0n : out std_logic;
    UUBEn : out std_logic;
    TAn : out std_logic;
    CLK40 : in std_logic;
    RnW : in std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    WEn : out std_logic;
    LLBEn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    RASn : out std_logic;
    CS1n : out std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic);
end U400_TOP;

-- Architecture of U400_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U400_TOP is

signal \N__7469\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3859\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3723\ : std_logic;
signal \N__3720\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3548\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3510\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3439\ : std_logic;
signal \N__3436\ : std_logic;
signal \N__3433\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3307\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3216\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2874\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2862\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2854\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2850\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2836\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2827\ : std_logic;
signal \N__2824\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2799\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2767\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2749\ : std_logic;
signal \CLK40_ibuf_gb_io_gb_input\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \INVU400_SDRAM.REFRESH_COUNTER_0C_net\ : std_logic;
signal \A_c_31\ : std_logic;
signal \A_c_27\ : std_logic;
signal \INVU400_SDRAM.REFRESH_COUNTER_1C_net\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_0\ : std_logic;
signal \bfn_2_4_0_\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_1\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_2\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_3\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_4\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_5\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_6\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_7\ : std_logic;
signal \INVU400_SDRAM.REFRESH_COUNTER_2C_net\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_8\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U400_SDRAM.un1_REFRESH_COUNTERlt7_0_cascade_\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \CASn_c\ : std_logic;
signal \WEn_c\ : std_logic;
signal \INVU400_SDRAM.CASnC_net\ : std_logic;
signal \RASn_c\ : std_logic;
signal \INVU400_SDRAM.RASnC_net\ : std_logic;
signal \A_c_30\ : std_logic;
signal \A_c_29\ : std_logic;
signal \A_c_28\ : std_logic;
signal \U400_ADDRESS_DECODE.m2Z0Z_1\ : std_logic;
signal \INVU400_SDRAM.SDRAM_COUNTER_1C_net\ : std_logic;
signal \INVU400_SDRAM.RAM_CYCLEC_net\ : std_logic;
signal \U400_ADDRESS_DECODE.N_185_cascade_\ : std_logic;
signal \U400_ADDRESS_DECODE.m84_amZ0_cascade_\ : std_logic;
signal \U400_ADDRESS_DECODE.m84_bmZ0\ : std_logic;
signal \N_85_0\ : std_logic;
signal \U400_ADDRESS_DECODE.N_46_0\ : std_logic;
signal \U400_ADDRESS_DECODE.N_47_0_cascade_\ : std_logic;
signal \U400_ADDRESS_DECODE.m71_amZ0Z_1\ : std_logic;
signal \U400_ADDRESS_DECODE.m71_amZ0_cascade_\ : std_logic;
signal \U400_ADDRESS_DECODE.m71_bmZ0\ : std_logic;
signal \U400_ADDRESS_DECODE.N_72_0_cascade_\ : std_logic;
signal \N_73_0_cascade_\ : std_logic;
signal \INVU400_SDRAM.SDRAM_CMD_2C_net\ : std_logic;
signal \U400_ADDRESS_DECODE.m56_amZ0\ : std_logic;
signal \N_57_0\ : std_logic;
signal \U400_ADDRESS_DECODE.N_7_0_cascade_\ : std_logic;
signal \INVU400_SDRAM.SDRAM_CMD_0C_net\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_17\ : std_logic;
signal \MA_c_7\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_24\ : std_logic;
signal \MA_c_8\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_7C_net\ : std_logic;
signal \A_c_8\ : std_logic;
signal \A_c_16\ : std_logic;
signal \MA_c_6\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_6C_net\ : std_logic;
signal \bfn_5_3_0_\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_s_1\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_s_3\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \INVU400_SDRAM.SDRAM_COUNTER_2C_net\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \N_60_cascade_\ : std_logic;
signal \U400_ADDRESS_DECODE.N_98_0_cascade_\ : std_logic;
signal \U400_SDRAM_SDRAM_CMD_5_sqmuxa\ : std_logic;
signal \U400_ADDRESS_DECODE.m41_amZ0_cascade_\ : std_logic;
signal \U400_ADDRESS_DECODE.m41_bmZ0\ : std_logic;
signal \U400_ADDRESS_DECODE.m54Z0Z_0_cascade_\ : std_logic;
signal \U400_ADDRESS_DECODE.m56_bmZ0\ : std_logic;
signal \U400_ADDRESS_DECODE.N_185\ : std_logic;
signal \U400_ADDRESS_DECODE.N_185_mux_cascade_\ : std_logic;
signal \U400_ADDRESS_DECODE.N_42_0\ : std_logic;
signal \U400_ADDRESS_DECODE.m43_bmZ0_cascade_\ : std_logic;
signal \N_44_0\ : std_logic;
signal \U400_ADDRESS_DECODE.N_33_0\ : std_logic;
signal \U400_ADDRESS_DECODE.m43_amZ0\ : std_logic;
signal \U400_ADDRESS_DECODE.m87_nsZ0Z_1\ : std_logic;
signal \U400_ADDRESS_DECODE.N_88_0_cascade_\ : std_logic;
signal \N_96_0_cascade_\ : std_logic;
signal \N_73_0\ : std_logic;
signal \INVU400_SDRAM.SDRAM_CMD_1C_net\ : std_logic;
signal \U400_ADDRESS_DECODE.m63_nsZ0Z_1\ : std_logic;
signal \U400_ADDRESS_DECODE.N_139_0_cascade_\ : std_logic;
signal \U400_ADDRESS_DECODE.m133Z0Z_0\ : std_logic;
signal \U400_ADDRESS_DECODE.N_47_0\ : std_logic;
signal \U400_ADDRESS_DECODE.N_62_0\ : std_logic;
signal \U400_ADDRESS_DECODE.N_62_0_cascade_\ : std_logic;
signal \U400_ADDRESS_DECODE.m141_bmZ0_cascade_\ : std_logic;
signal \U400_ADDRESS_DECODE.m141_amZ0\ : std_logic;
signal \U400_SDRAM.CS0_ENZ0\ : std_logic;
signal \CS0n_c\ : std_logic;
signal \INVU400_SDRAM.CS0_ENC_net\ : std_logic;
signal \A_c_26\ : std_logic;
signal \MA_c_12\ : std_logic;
signal \A_c_19\ : std_logic;
signal \MA_c_9\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_12C_net\ : std_logic;
signal \U400_SDRAM_RAM_CYCLE\ : std_logic;
signal \U400_SDRAM_RAM_CYCLE_START_2_0\ : std_logic;
signal \U400_ADDRESS_DECODE.N_8_0_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_CONFIGURED_RNIJKCAZ0Z2\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U400_ADDRESS_DECODE.m165_nsZ0Z_1\ : std_logic;
signal \N_13_0_cascade_\ : std_logic;
signal \U400_ADDRESS_DECODE.N_10_0\ : std_logic;
signal \U400_ADDRESS_DECODE.N_8_0\ : std_logic;
signal \U400_ADDRESS_DECODE.N_179_mux_cascade_\ : std_logic;
signal \U400_ADDRESS_DECODE.m94_amZ0Z_1\ : std_logic;
signal \U400_ADDRESS_DECODE.m94_amZ0_cascade_\ : std_logic;
signal \U400_ADDRESS_DECODE.N_95_0\ : std_logic;
signal \U400_SDRAM_RAM_CYCLE_START\ : std_logic;
signal \U400_ADDRESS_DECODE.N_15_0\ : std_logic;
signal \N_13_0\ : std_logic;
signal \U400_SDRAM_SDRAM_CMD11\ : std_logic;
signal \U400_ADDRESS_DECODE.m20_amZ0_cascade_\ : std_logic;
signal \U400_SDRAM_SDRAM_COUNTER_3\ : std_logic;
signal \U400_ADDRESS_DECODE.N_6_0\ : std_logic;
signal \U400_ADDRESS_DECODE.m94_bmZ0\ : std_logic;
signal \U400_SDRAM_SDRAM_COUNTER_1\ : std_logic;
signal \U400_ADDRESS_DECODE.m20_bmZ0\ : std_logic;
signal \U400_ADDRESS_DECODE.N_20_0\ : std_logic;
signal \U400_ADDRESS_DECODE.N_179_mux\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U400_SDRAM_WRITE_CYCLE\ : std_logic;
signal \N_48\ : std_logic;
signal \N_142_0\ : std_logic;
signal \INVU400_SDRAM.WRITE_CYCLEC_net\ : std_logic;
signal \U400_ADDRESS_DECODE.N_12_0\ : std_logic;
signal \U400_ADDRESS_DECODE.N_21_0\ : std_logic;
signal \A_c_23\ : std_logic;
signal \N_137_0\ : std_logic;
signal \N_190_mux\ : std_logic;
signal \N_138_0\ : std_logic;
signal \N_23_0\ : std_logic;
signal \U400_SDRAM.CS1_ENZ0\ : std_logic;
signal \CS1n_c\ : std_logic;
signal \INVU400_SDRAM.CS1_ENC_net\ : std_logic;
signal \U400_SDRAM_TA_COUNTER_4\ : std_logic;
signal \U400_SDRAM_TA_COUNTER_1\ : std_logic;
signal \U400_ADDRESS_DECODE.N_177_mux_cascade_\ : std_logic;
signal \U400_SDRAM_TA_COUNTER_0\ : std_logic;
signal \U400_SDRAM_TACK\ : std_logic;
signal \U400_SDRAM_TA_COUNTER_5\ : std_logic;
signal \U400_SDRAM.N_252_0_0_cascade_\ : std_logic;
signal \U400_SDRAM_TA_COUNTER_2\ : std_logic;
signal \U400_SDRAM_TA_COUNTER_3\ : std_logic;
signal \A_c_22\ : std_logic;
signal \BANK1_c\ : std_logic;
signal \A_c_21\ : std_logic;
signal \U400_SDRAM_un1_SDRAM_COUNTER59_2_0\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \U400_SDRAM_SDRAM_CMD_1_sqmuxa_1\ : std_logic;
signal \INVU400_SDRAM.BANK1C_net\ : std_logic;
signal \U400_SDRAM_SDRAM_COUNTER_2\ : std_logic;
signal \N_60\ : std_logic;
signal \U400_ADDRESS_DECODE.m145_nsZ0Z_1\ : std_logic;
signal \N_100_0_i\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U400_SDRAM_SDRAM_COUNTER_0\ : std_logic;
signal \INVU400_SDRAM.SDRAM_COUNTER_0C_net\ : std_logic;
signal \U400_SDRAM_SDRAM_COUNTERe_0_i\ : std_logic;
signal \U400_ADDRESS_DECODE.N_135_0\ : std_logic;
signal \U400_ADDRESS_DECODE.N_146_0\ : std_logic;
signal \N_14_i\ : std_logic;
signal \U400_ADDRESS_DECODE.N_147_0_cascade_\ : std_logic;
signal \U400_ADDRESS_DECODE.N_136_0\ : std_logic;
signal \N_43\ : std_logic;
signal \A_c_20\ : std_logic;
signal \MA_c_10\ : std_logic;
signal \A_c_25\ : std_logic;
signal \MA_c_11\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_10C_net\ : std_logic;
signal \U400_ADDRESS_DECODE.N_4_0_cascade_\ : std_logic;
signal \N_124_0\ : std_logic;
signal \U400_SDRAM.N_252_0_0\ : std_logic;
signal \U400_SDRAM.N_252_0_0_en\ : std_logic;
signal \N_174\ : std_logic;
signal \U400_SDRAM_TA_OUT_5_0\ : std_logic;
signal \U400_SDRAM_N_252_0\ : std_logic;
signal \TA_OUT\ : std_logic;
signal \CLK40_c_g\ : std_logic;
signal \U400_SDRAM_BURST\ : std_logic;
signal \U400_ADDRESS_DECODE.N_114_0\ : std_logic;
signal \N_65_0\ : std_logic;
signal \U400_SDRAM_SDRAM_CONFIGURED\ : std_logic;
signal \INVU400_SDRAM.SDRAM_CONFIGUREDC_net\ : std_logic;
signal \N_129_0\ : std_logic;
signal \N_127_0\ : std_logic;
signal \A_c_1\ : std_logic;
signal \N_128_0\ : std_logic;
signal \U400_ADDRESS_DECODE.N_122_0\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \A_c_0\ : std_logic;
signal \U400_ADDRESS_DECODE.N_4_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \U400_ADDRESS_DECODE.N_186_mux\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U400_SDRAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U400_SDRAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U400_SDRAM.MA_5_iv_0_1\ : std_logic;
signal \MA_c_1\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U400_SDRAM.MA_5_iv_0_5\ : std_logic;
signal \MA_c_5\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_13\ : std_logic;
signal \MA_c_3\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_1C_net\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_12\ : std_logic;
signal \MA_c_2\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_14\ : std_logic;
signal \MA_c_4\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U400_SDRAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U400_SDRAM.MA19\ : std_logic;
signal \MA_c_0\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_2C_net\ : std_logic;
signal \U400_SDRAM.un1_MA20_0_i_0\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \U400_ADDRESS_DECODE.N_170_mux\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \N_4_0_i\ : std_logic;
signal \TA_EN_i\ : std_logic;
signal \N_304_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \MA_wire\ : std_logic_vector(12 downto 0);
signal \A_wire\ : std_logic_vector(31 downto 0);
signal \CASn_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \UUBEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \LLBEn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \TAn_wire\ : std_logic;
signal \LBENn_wire\ : std_logic;
signal \CS1n_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CS0n_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CLK40_wire\ : std_logic;

begin
    MA <= \MA_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    BANK1 <= \BANK1_wire\;
    UUBEn <= \UUBEn_wire\;
    \SIZ_wire\ <= SIZ;
    LLBEn <= \LLBEn_wire\;
    \TSn_wire\ <= TSn;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    \RESETn_wire\ <= RESETn;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    TAn <= \TAn_wire\;
    LBENn <= \LBENn_wire\;
    CS1n <= \CS1n_wire\;
    WEn <= \WEn_wire\;
    \RnW_wire\ <= RnW;
    CS0n <= \CS0n_wire\;
    LMBEn <= \LMBEn_wire\;
    \CLK40_wire\ <= CLK40;

    \MA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7469\,
            DIN => \N__7468\,
            DOUT => \N__7467\,
            PACKAGEPIN => \MA_wire\(7)
        );

    \MA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7469\,
            PADOUT => \N__7468\,
            PADIN => \N__7467\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3037\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7460\,
            DIN => \N__7459\,
            DOUT => \N__7458\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7460\,
            PADOUT => \N__7459\,
            PADIN => \N__7458\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7451\,
            DIN => \N__7450\,
            DOUT => \N__7449\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7451\,
            PADOUT => \N__7450\,
            PADIN => \N__7449\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2839\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7442\,
            DIN => \N__7441\,
            DOUT => \N__7440\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7442\,
            PADOUT => \N__7441\,
            PADIN => \N__7440\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5104\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7433\,
            DIN => \N__7432\,
            DOUT => \N__7431\,
            PACKAGEPIN => \MA_wire\(8)
        );

    \MA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7433\,
            PADOUT => \N__7432\,
            PADIN => \N__7431\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3175\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7424\,
            DIN => \N__7423\,
            DOUT => \N__7422\,
            PACKAGEPIN => \MA_wire\(10)
        );

    \MA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7424\,
            PADOUT => \N__7423\,
            PADIN => \N__7422\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5356\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7415\,
            DIN => \N__7414\,
            DOUT => \N__7413\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7415\,
            PADOUT => \N__7414\,
            PADIN => \N__7413\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7406\,
            DIN => \N__7405\,
            DOUT => \N__7404\,
            PACKAGEPIN => \MA_wire\(2)
        );

    \MA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7406\,
            PADOUT => \N__7405\,
            PADIN => \N__7404\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6097\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7397\,
            DIN => \N__7396\,
            DOUT => \N__7395\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7397\,
            PADOUT => \N__7396\,
            PADIN => \N__7395\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7388\,
            DIN => \N__7387\,
            DOUT => \N__7386\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7388\,
            PADOUT => \N__7387\,
            PADIN => \N__7386\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7379\,
            DIN => \N__7378\,
            DOUT => \N__7377\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7379\,
            PADOUT => \N__7378\,
            PADIN => \N__7377\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5317\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7370\,
            DIN => \N__7369\,
            DOUT => \N__7368\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7370\,
            PADOUT => \N__7369\,
            PADIN => \N__7368\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7361\,
            DIN => \N__7360\,
            DOUT => \N__7359\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7361\,
            PADOUT => \N__7360\,
            PADIN => \N__7359\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7352\,
            DIN => \N__7351\,
            DOUT => \N__7350\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7352\,
            PADOUT => \N__7351\,
            PADIN => \N__7350\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7343\,
            DIN => \N__7342\,
            DOUT => \N__7341\,
            PACKAGEPIN => \MA_wire\(12)
        );

    \MA_obuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7343\,
            PADOUT => \N__7342\,
            PADIN => \N__7341\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3469\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7334\,
            DIN => \N__7333\,
            DOUT => \N__7332\,
            PACKAGEPIN => \MA_wire\(1)
        );

    \MA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7334\,
            PADOUT => \N__7333\,
            PADIN => \N__7332\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6208\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7325\,
            DIN => \N__7324\,
            DOUT => \N__7323\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7325\,
            PADOUT => \N__7324\,
            PADIN => \N__7323\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7316\,
            DIN => \N__7315\,
            DOUT => \N__7314\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7316\,
            PADOUT => \N__7315\,
            PADIN => \N__7314\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7307\,
            DIN => \N__7306\,
            DOUT => \N__7305\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7307\,
            PADOUT => \N__7306\,
            PADIN => \N__7305\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7298\,
            DIN => \N__7297\,
            DOUT => \N__7296\,
            PACKAGEPIN => \MA_wire\(4)
        );

    \MA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7298\,
            PADOUT => \N__7297\,
            PADIN => \N__7296\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6064\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7289\,
            DIN => \N__7288\,
            DOUT => \N__7287\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7289\,
            PADOUT => \N__7288\,
            PADIN => \N__7287\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7280\,
            DIN => \N__7279\,
            DOUT => \N__7278\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7280\,
            PADOUT => \N__7279\,
            PADIN => \N__7278\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7271\,
            DIN => \N__7270\,
            DOUT => \N__7269\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7271\,
            PADOUT => \N__7270\,
            PADIN => \N__7269\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5668\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7262\,
            DIN => \N__7261\,
            DOUT => \N__7260\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7262\,
            PADOUT => \N__7261\,
            PADIN => \N__7260\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7253\,
            DIN => \N__7252\,
            DOUT => \N__7251\,
            PACKAGEPIN => \MA_wire\(9)
        );

    \MA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7253\,
            PADOUT => \N__7252\,
            PADIN => \N__7251\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3442\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7244\,
            DIN => \N__7243\,
            DOUT => \N__7242\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7244\,
            PADOUT => \N__7243\,
            PADIN => \N__7242\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5659\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7235\,
            DIN => \N__7234\,
            DOUT => \N__7233\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7235\,
            PADOUT => \N__7234\,
            PADIN => \N__7233\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7226\,
            DIN => \N__7225\,
            DOUT => \N__7224\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7226\,
            PADOUT => \N__7225\,
            PADIN => \N__7224\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7217\,
            DIN => \N__7216\,
            DOUT => \N__7215\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7217\,
            PADOUT => \N__7216\,
            PADIN => \N__7215\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4687\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7208\,
            DIN => \N__7207\,
            DOUT => \N__7206\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7208\,
            PADOUT => \N__7207\,
            PADIN => \N__7206\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7199\,
            DIN => \N__7198\,
            DOUT => \N__7197\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7199\,
            PADOUT => \N__7198\,
            PADIN => \N__7197\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7190\,
            DIN => \N__7189\,
            DOUT => \N__7188\,
            PACKAGEPIN => \MA_wire\(3)
        );

    \MA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7190\,
            PADOUT => \N__7189\,
            PADIN => \N__7188\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6139\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7181\,
            DIN => \N__7180\,
            DOUT => \N__7179\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7181\,
            PADOUT => \N__7180\,
            PADIN => \N__7179\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7172\,
            DIN => \N__7171\,
            DOUT => \N__7170\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7172\,
            PADOUT => \N__7171\,
            PADIN => \N__7170\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7163\,
            DIN => \N__7162\,
            DOUT => \N__7161\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7163\,
            PADOUT => \N__7162\,
            PADIN => \N__7161\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7154\,
            DIN => \N__7153\,
            DOUT => \N__7152\,
            PACKAGEPIN => \MA_wire\(6)
        );

    \MA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7154\,
            PADOUT => \N__7153\,
            PADIN => \N__7152\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3136\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7145\,
            DIN => \N__7144\,
            DOUT => \N__7143\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7145\,
            PADOUT => \N__7144\,
            PADIN => \N__7143\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7136\,
            DIN => \N__7135\,
            DOUT => \N__7134\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7136\,
            PADOUT => \N__7135\,
            PADIN => \N__7134\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7127\,
            DIN => \N__7126\,
            DOUT => \N__7125\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7127\,
            PADOUT => \N__7126\,
            PADIN => \N__7125\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7118\,
            DIN => \N__7117\,
            DOUT => \N__7116\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7118\,
            PADOUT => \N__7117\,
            PADIN => \N__7116\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2986\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7109\,
            DIN => \N__7108\,
            DOUT => \N__7107\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7109\,
            PADOUT => \N__7108\,
            PADIN => \N__7107\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7100\,
            DIN => \N__7099\,
            DOUT => \N__7098\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7100\,
            PADOUT => \N__7099\,
            PADIN => \N__7098\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5053\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7091\,
            DIN => \N__7090\,
            DOUT => \N__7089\,
            PACKAGEPIN => \MA_wire\(11)
        );

    \MA_obuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7091\,
            PADOUT => \N__7090\,
            PADIN => \N__7089\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5329\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TAn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7082\,
            DIN => \N__7081\,
            DOUT => \N__7080\,
            PACKAGEPIN => \TAn_wire\
        );

    \TAn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7082\,
            PADOUT => \N__7081\,
            PADIN => \N__7080\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6427\,
            DIN0 => OPEN,
            DOUT0 => \N__5269\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7073\,
            DIN => \N__7072\,
            DOUT => \N__7071\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7073\,
            PADOUT => \N__7072\,
            PADIN => \N__7071\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7064\,
            DIN => \N__7063\,
            DOUT => \N__7062\,
            PACKAGEPIN => \MA_wire\(5)
        );

    \MA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7064\,
            PADOUT => \N__7063\,
            PADIN => \N__7062\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6184\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7055\,
            DIN => \N__7054\,
            DOUT => \N__7053\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7055\,
            PADOUT => \N__7054\,
            PADIN => \N__7053\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7046\,
            DIN => \N__7045\,
            DOUT => \N__7044\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7046\,
            PADOUT => \N__7045\,
            PADIN => \N__7044\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LBENn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7037\,
            DIN => \N__7036\,
            DOUT => \N__7035\,
            PACKAGEPIN => \LBENn_wire\
        );

    \LBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7037\,
            PADOUT => \N__7036\,
            PADIN => \N__7035\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6454\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7028\,
            DIN => \N__7027\,
            DOUT => \N__7026\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7028\,
            PADOUT => \N__7027\,
            PADIN => \N__7026\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CS1n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7019\,
            DIN => \N__7018\,
            DOUT => \N__7017\,
            PACKAGEPIN => \CS1n_wire\
        );

    \CS1n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7019\,
            PADOUT => \N__7018\,
            PADIN => \N__7017\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4174\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7010\,
            DIN => \N__7009\,
            DOUT => \N__7008\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7010\,
            PADOUT => \N__7009\,
            PADIN => \N__7008\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7001\,
            DIN => \N__7000\,
            DOUT => \N__6999\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7001\,
            PADOUT => \N__7000\,
            PADIN => \N__6999\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6992\,
            DIN => \N__6991\,
            DOUT => \N__6990\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6992\,
            PADOUT => \N__6991\,
            PADIN => \N__6990\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6983\,
            DIN => \N__6982\,
            DOUT => \N__6981\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6983\,
            PADOUT => \N__6982\,
            PADIN => \N__6981\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6974\,
            DIN => \N__6973\,
            DOUT => \N__6972\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6974\,
            PADOUT => \N__6973\,
            PADIN => \N__6972\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2995\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6965\,
            DIN => \N__6964\,
            DOUT => \N__6963\,
            PACKAGEPIN => \MA_wire\(0)
        );

    \MA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6965\,
            PADOUT => \N__6964\,
            PADIN => \N__6963\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6808\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6956\,
            DIN => \N__6955\,
            DOUT => \N__6954\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6956\,
            PADOUT => \N__6955\,
            PADIN => \N__6954\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6947\,
            DIN => \N__6946\,
            DOUT => \N__6945\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6947\,
            PADOUT => \N__6946\,
            PADIN => \N__6945\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6938\,
            DIN => \N__6937\,
            DOUT => \N__6936\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6938\,
            PADOUT => \N__6937\,
            PADIN => \N__6936\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CS0n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6929\,
            DIN => \N__6928\,
            DOUT => \N__6927\,
            PACKAGEPIN => \CS0n_wire\
        );

    \CS0n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6929\,
            PADOUT => \N__6928\,
            PADIN => \N__6927\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3505\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6920\,
            DIN => \N__6919\,
            DOUT => \N__6918\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6920\,
            PADOUT => \N__6919\,
            PADIN => \N__6918\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6911\,
            DIN => \N__6910\,
            DOUT => \N__6909\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6911\,
            PADOUT => \N__6910\,
            PADIN => \N__6909\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5614\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6902\,
            DIN => \N__6901\,
            DOUT => \N__6900\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6902\,
            PADOUT => \N__6901\,
            PADIN => \N__6900\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6893\,
            DIN => \N__6892\,
            DOUT => \N__6891\,
            PACKAGEPIN => \CLK40_wire\
        );

    \CLK40_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6893\,
            PADOUT => \N__6892\,
            PADIN => \N__6891\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_ibuf_gb_io_gb_input\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__6874\,
            I => \N__6871\
        );

    \I__1626\ : InMux
    port map (
            O => \N__6871\,
            I => \N__6868\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__6868\,
            I => \N__6865\
        );

    \I__1624\ : Span4Mux_s1_v
    port map (
            O => \N__6865\,
            I => \N__6862\
        );

    \I__1623\ : Odrv4
    port map (
            O => \N__6862\,
            I => \A_c_10\
        );

    \I__1622\ : InMux
    port map (
            O => \N__6859\,
            I => \N__6853\
        );

    \I__1621\ : InMux
    port map (
            O => \N__6858\,
            I => \N__6853\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__6853\,
            I => \N__6846\
        );

    \I__1619\ : InMux
    port map (
            O => \N__6852\,
            I => \N__6843\
        );

    \I__1618\ : InMux
    port map (
            O => \N__6851\,
            I => \N__6836\
        );

    \I__1617\ : InMux
    port map (
            O => \N__6850\,
            I => \N__6836\
        );

    \I__1616\ : InMux
    port map (
            O => \N__6849\,
            I => \N__6836\
        );

    \I__1615\ : Span4Mux_h
    port map (
            O => \N__6846\,
            I => \N__6830\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__6843\,
            I => \N__6827\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__6836\,
            I => \N__6824\
        );

    \I__1612\ : InMux
    port map (
            O => \N__6835\,
            I => \N__6817\
        );

    \I__1611\ : InMux
    port map (
            O => \N__6834\,
            I => \N__6817\
        );

    \I__1610\ : InMux
    port map (
            O => \N__6833\,
            I => \N__6817\
        );

    \I__1609\ : Odrv4
    port map (
            O => \N__6830\,
            I => \U400_SDRAM.MA19\
        );

    \I__1608\ : Odrv12
    port map (
            O => \N__6827\,
            I => \U400_SDRAM.MA19\
        );

    \I__1607\ : Odrv4
    port map (
            O => \N__6824\,
            I => \U400_SDRAM.MA19\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__6817\,
            I => \U400_SDRAM.MA19\
        );

    \I__1605\ : IoInMux
    port map (
            O => \N__6808\,
            I => \N__6805\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__6805\,
            I => \MA_c_0\
        );

    \I__1603\ : CEMux
    port map (
            O => \N__6802\,
            I => \N__6797\
        );

    \I__1602\ : CEMux
    port map (
            O => \N__6801\,
            I => \N__6794\
        );

    \I__1601\ : CEMux
    port map (
            O => \N__6800\,
            I => \N__6791\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__6797\,
            I => \N__6787\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__6794\,
            I => \N__6784\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__6791\,
            I => \N__6781\
        );

    \I__1597\ : CEMux
    port map (
            O => \N__6790\,
            I => \N__6778\
        );

    \I__1596\ : Span4Mux_v
    port map (
            O => \N__6787\,
            I => \N__6767\
        );

    \I__1595\ : Span4Mux_h
    port map (
            O => \N__6784\,
            I => \N__6767\
        );

    \I__1594\ : Span4Mux_s2_v
    port map (
            O => \N__6781\,
            I => \N__6767\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__6778\,
            I => \N__6767\
        );

    \I__1592\ : CEMux
    port map (
            O => \N__6777\,
            I => \N__6764\
        );

    \I__1591\ : CEMux
    port map (
            O => \N__6776\,
            I => \N__6761\
        );

    \I__1590\ : Odrv4
    port map (
            O => \N__6767\,
            I => \U400_SDRAM.un1_MA20_0_i_0\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__6764\,
            I => \U400_SDRAM.un1_MA20_0_i_0\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__6761\,
            I => \U400_SDRAM.un1_MA20_0_i_0\
        );

    \I__1587\ : CascadeMux
    port map (
            O => \N__6754\,
            I => \N__6751\
        );

    \I__1586\ : InMux
    port map (
            O => \N__6751\,
            I => \N__6748\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__6748\,
            I => \N__6743\
        );

    \I__1584\ : SRMux
    port map (
            O => \N__6747\,
            I => \N__6697\
        );

    \I__1583\ : SRMux
    port map (
            O => \N__6746\,
            I => \N__6697\
        );

    \I__1582\ : Glb2LocalMux
    port map (
            O => \N__6743\,
            I => \N__6697\
        );

    \I__1581\ : SRMux
    port map (
            O => \N__6742\,
            I => \N__6697\
        );

    \I__1580\ : SRMux
    port map (
            O => \N__6741\,
            I => \N__6697\
        );

    \I__1579\ : SRMux
    port map (
            O => \N__6740\,
            I => \N__6697\
        );

    \I__1578\ : SRMux
    port map (
            O => \N__6739\,
            I => \N__6697\
        );

    \I__1577\ : SRMux
    port map (
            O => \N__6738\,
            I => \N__6697\
        );

    \I__1576\ : SRMux
    port map (
            O => \N__6737\,
            I => \N__6697\
        );

    \I__1575\ : SRMux
    port map (
            O => \N__6736\,
            I => \N__6697\
        );

    \I__1574\ : SRMux
    port map (
            O => \N__6735\,
            I => \N__6697\
        );

    \I__1573\ : SRMux
    port map (
            O => \N__6734\,
            I => \N__6697\
        );

    \I__1572\ : SRMux
    port map (
            O => \N__6733\,
            I => \N__6697\
        );

    \I__1571\ : SRMux
    port map (
            O => \N__6732\,
            I => \N__6697\
        );

    \I__1570\ : SRMux
    port map (
            O => \N__6731\,
            I => \N__6697\
        );

    \I__1569\ : SRMux
    port map (
            O => \N__6730\,
            I => \N__6697\
        );

    \I__1568\ : GlobalMux
    port map (
            O => \N__6697\,
            I => \N__6694\
        );

    \I__1567\ : gio2CtrlBuf
    port map (
            O => \N__6694\,
            I => \RESETn_c_i_g\
        );

    \I__1566\ : CascadeMux
    port map (
            O => \N__6691\,
            I => \N__6688\
        );

    \I__1565\ : InMux
    port map (
            O => \N__6688\,
            I => \N__6682\
        );

    \I__1564\ : CascadeMux
    port map (
            O => \N__6687\,
            I => \N__6679\
        );

    \I__1563\ : InMux
    port map (
            O => \N__6686\,
            I => \N__6676\
        );

    \I__1562\ : InMux
    port map (
            O => \N__6685\,
            I => \N__6673\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__6682\,
            I => \N__6670\
        );

    \I__1560\ : InMux
    port map (
            O => \N__6679\,
            I => \N__6667\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__6676\,
            I => \N__6664\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__6673\,
            I => \N__6661\
        );

    \I__1557\ : Span4Mux_h
    port map (
            O => \N__6670\,
            I => \N__6656\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__6667\,
            I => \N__6656\
        );

    \I__1555\ : Span12Mux_s8_h
    port map (
            O => \N__6664\,
            I => \N__6653\
        );

    \I__1554\ : Span4Mux_v
    port map (
            O => \N__6661\,
            I => \N__6650\
        );

    \I__1553\ : Span4Mux_v
    port map (
            O => \N__6656\,
            I => \N__6647\
        );

    \I__1552\ : Odrv12
    port map (
            O => \N__6653\,
            I => \U400_ADDRESS_DECODE.N_170_mux\
        );

    \I__1551\ : Odrv4
    port map (
            O => \N__6650\,
            I => \U400_ADDRESS_DECODE.N_170_mux\
        );

    \I__1550\ : Odrv4
    port map (
            O => \N__6647\,
            I => \U400_ADDRESS_DECODE.N_170_mux\
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__6640\,
            I => \N__6636\
        );

    \I__1548\ : InMux
    port map (
            O => \N__6639\,
            I => \N__6632\
        );

    \I__1547\ : InMux
    port map (
            O => \N__6636\,
            I => \N__6627\
        );

    \I__1546\ : InMux
    port map (
            O => \N__6635\,
            I => \N__6627\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__6632\,
            I => \N__6621\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__6627\,
            I => \N__6618\
        );

    \I__1543\ : InMux
    port map (
            O => \N__6626\,
            I => \N__6613\
        );

    \I__1542\ : InMux
    port map (
            O => \N__6625\,
            I => \N__6613\
        );

    \I__1541\ : CascadeMux
    port map (
            O => \N__6624\,
            I => \N__6599\
        );

    \I__1540\ : Span4Mux_s3_v
    port map (
            O => \N__6621\,
            I => \N__6591\
        );

    \I__1539\ : Span4Mux_h
    port map (
            O => \N__6618\,
            I => \N__6591\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__6613\,
            I => \N__6591\
        );

    \I__1537\ : InMux
    port map (
            O => \N__6612\,
            I => \N__6588\
        );

    \I__1536\ : InMux
    port map (
            O => \N__6611\,
            I => \N__6585\
        );

    \I__1535\ : CascadeMux
    port map (
            O => \N__6610\,
            I => \N__6582\
        );

    \I__1534\ : InMux
    port map (
            O => \N__6609\,
            I => \N__6575\
        );

    \I__1533\ : InMux
    port map (
            O => \N__6608\,
            I => \N__6575\
        );

    \I__1532\ : InMux
    port map (
            O => \N__6607\,
            I => \N__6572\
        );

    \I__1531\ : InMux
    port map (
            O => \N__6606\,
            I => \N__6569\
        );

    \I__1530\ : InMux
    port map (
            O => \N__6605\,
            I => \N__6562\
        );

    \I__1529\ : InMux
    port map (
            O => \N__6604\,
            I => \N__6562\
        );

    \I__1528\ : InMux
    port map (
            O => \N__6603\,
            I => \N__6562\
        );

    \I__1527\ : InMux
    port map (
            O => \N__6602\,
            I => \N__6557\
        );

    \I__1526\ : InMux
    port map (
            O => \N__6599\,
            I => \N__6557\
        );

    \I__1525\ : CascadeMux
    port map (
            O => \N__6598\,
            I => \N__6552\
        );

    \I__1524\ : Span4Mux_h
    port map (
            O => \N__6591\,
            I => \N__6547\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__6588\,
            I => \N__6547\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__6585\,
            I => \N__6544\
        );

    \I__1521\ : InMux
    port map (
            O => \N__6582\,
            I => \N__6541\
        );

    \I__1520\ : InMux
    port map (
            O => \N__6581\,
            I => \N__6538\
        );

    \I__1519\ : InMux
    port map (
            O => \N__6580\,
            I => \N__6535\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__6575\,
            I => \N__6530\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__6572\,
            I => \N__6530\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__6569\,
            I => \N__6523\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__6562\,
            I => \N__6523\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__6557\,
            I => \N__6523\
        );

    \I__1513\ : InMux
    port map (
            O => \N__6556\,
            I => \N__6520\
        );

    \I__1512\ : InMux
    port map (
            O => \N__6555\,
            I => \N__6516\
        );

    \I__1511\ : InMux
    port map (
            O => \N__6552\,
            I => \N__6513\
        );

    \I__1510\ : Span4Mux_v
    port map (
            O => \N__6547\,
            I => \N__6510\
        );

    \I__1509\ : Span4Mux_h
    port map (
            O => \N__6544\,
            I => \N__6505\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__6541\,
            I => \N__6505\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__6538\,
            I => \N__6500\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__6535\,
            I => \N__6500\
        );

    \I__1505\ : Span4Mux_v
    port map (
            O => \N__6530\,
            I => \N__6493\
        );

    \I__1504\ : Span4Mux_h
    port map (
            O => \N__6523\,
            I => \N__6493\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__6520\,
            I => \N__6493\
        );

    \I__1502\ : InMux
    port map (
            O => \N__6519\,
            I => \N__6490\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__6516\,
            I => \N__6485\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__6513\,
            I => \N__6485\
        );

    \I__1499\ : Span4Mux_h
    port map (
            O => \N__6510\,
            I => \N__6480\
        );

    \I__1498\ : Span4Mux_h
    port map (
            O => \N__6505\,
            I => \N__6480\
        );

    \I__1497\ : Span4Mux_v
    port map (
            O => \N__6500\,
            I => \N__6477\
        );

    \I__1496\ : Span4Mux_h
    port map (
            O => \N__6493\,
            I => \N__6472\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__6490\,
            I => \N__6472\
        );

    \I__1494\ : Span12Mux_s8_v
    port map (
            O => \N__6485\,
            I => \N__6469\
        );

    \I__1493\ : IoSpan4Mux
    port map (
            O => \N__6480\,
            I => \N__6466\
        );

    \I__1492\ : Span4Mux_h
    port map (
            O => \N__6477\,
            I => \N__6461\
        );

    \I__1491\ : Span4Mux_v
    port map (
            O => \N__6472\,
            I => \N__6461\
        );

    \I__1490\ : Odrv12
    port map (
            O => \N__6469\,
            I => \RESETn_c\
        );

    \I__1489\ : Odrv4
    port map (
            O => \N__6466\,
            I => \RESETn_c\
        );

    \I__1488\ : Odrv4
    port map (
            O => \N__6461\,
            I => \RESETn_c\
        );

    \I__1487\ : IoInMux
    port map (
            O => \N__6454\,
            I => \N__6451\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__6451\,
            I => \N__6448\
        );

    \I__1485\ : Odrv4
    port map (
            O => \N__6448\,
            I => \N_4_0_i\
        );

    \I__1484\ : InMux
    port map (
            O => \N__6445\,
            I => \N__6442\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__6442\,
            I => \N__6439\
        );

    \I__1482\ : Span4Mux_v
    port map (
            O => \N__6439\,
            I => \N__6435\
        );

    \I__1481\ : InMux
    port map (
            O => \N__6438\,
            I => \N__6432\
        );

    \I__1480\ : Odrv4
    port map (
            O => \N__6435\,
            I => \TA_EN_i\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__6432\,
            I => \TA_EN_i\
        );

    \I__1478\ : IoInMux
    port map (
            O => \N__6427\,
            I => \N__6424\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__6424\,
            I => \N__6421\
        );

    \I__1476\ : Odrv4
    port map (
            O => \N__6421\,
            I => \N_304_i\
        );

    \I__1475\ : InMux
    port map (
            O => \N__6418\,
            I => \N__6415\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__6415\,
            I => \N__6412\
        );

    \I__1473\ : Odrv4
    port map (
            O => \N__6412\,
            I => \A_c_7\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__6409\,
            I => \N__6404\
        );

    \I__1471\ : InMux
    port map (
            O => \N__6408\,
            I => \N__6396\
        );

    \I__1470\ : InMux
    port map (
            O => \N__6407\,
            I => \N__6396\
        );

    \I__1469\ : InMux
    port map (
            O => \N__6404\,
            I => \N__6391\
        );

    \I__1468\ : InMux
    port map (
            O => \N__6403\,
            I => \N__6391\
        );

    \I__1467\ : InMux
    port map (
            O => \N__6402\,
            I => \N__6383\
        );

    \I__1466\ : InMux
    port map (
            O => \N__6401\,
            I => \N__6383\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__6396\,
            I => \N__6380\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__6391\,
            I => \N__6377\
        );

    \I__1463\ : InMux
    port map (
            O => \N__6390\,
            I => \N__6372\
        );

    \I__1462\ : InMux
    port map (
            O => \N__6389\,
            I => \N__6372\
        );

    \I__1461\ : InMux
    port map (
            O => \N__6388\,
            I => \N__6368\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__6383\,
            I => \N__6358\
        );

    \I__1459\ : Span4Mux_h
    port map (
            O => \N__6380\,
            I => \N__6358\
        );

    \I__1458\ : Span4Mux_h
    port map (
            O => \N__6377\,
            I => \N__6358\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__6372\,
            I => \N__6358\
        );

    \I__1456\ : InMux
    port map (
            O => \N__6371\,
            I => \N__6354\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__6368\,
            I => \N__6351\
        );

    \I__1454\ : InMux
    port map (
            O => \N__6367\,
            I => \N__6348\
        );

    \I__1453\ : Span4Mux_v
    port map (
            O => \N__6358\,
            I => \N__6345\
        );

    \I__1452\ : InMux
    port map (
            O => \N__6357\,
            I => \N__6342\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__6354\,
            I => \N__6339\
        );

    \I__1450\ : Span4Mux_h
    port map (
            O => \N__6351\,
            I => \N__6334\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__6348\,
            I => \N__6334\
        );

    \I__1448\ : Span4Mux_v
    port map (
            O => \N__6345\,
            I => \N__6331\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__6342\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_1\
        );

    \I__1446\ : Odrv4
    port map (
            O => \N__6339\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_1\
        );

    \I__1445\ : Odrv4
    port map (
            O => \N__6334\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_1\
        );

    \I__1444\ : Odrv4
    port map (
            O => \N__6331\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_1\
        );

    \I__1443\ : CascadeMux
    port map (
            O => \N__6322\,
            I => \N__6319\
        );

    \I__1442\ : InMux
    port map (
            O => \N__6319\,
            I => \N__6316\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__6316\,
            I => \N__6313\
        );

    \I__1440\ : IoSpan4Mux
    port map (
            O => \N__6313\,
            I => \N__6310\
        );

    \I__1439\ : Odrv4
    port map (
            O => \N__6310\,
            I => \A_c_3\
        );

    \I__1438\ : InMux
    port map (
            O => \N__6307\,
            I => \N__6299\
        );

    \I__1437\ : InMux
    port map (
            O => \N__6306\,
            I => \N__6299\
        );

    \I__1436\ : InMux
    port map (
            O => \N__6305\,
            I => \N__6292\
        );

    \I__1435\ : InMux
    port map (
            O => \N__6304\,
            I => \N__6292\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__6299\,
            I => \N__6285\
        );

    \I__1433\ : InMux
    port map (
            O => \N__6298\,
            I => \N__6280\
        );

    \I__1432\ : InMux
    port map (
            O => \N__6297\,
            I => \N__6280\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__6292\,
            I => \N__6277\
        );

    \I__1430\ : InMux
    port map (
            O => \N__6291\,
            I => \N__6272\
        );

    \I__1429\ : InMux
    port map (
            O => \N__6290\,
            I => \N__6272\
        );

    \I__1428\ : InMux
    port map (
            O => \N__6289\,
            I => \N__6269\
        );

    \I__1427\ : InMux
    port map (
            O => \N__6288\,
            I => \N__6266\
        );

    \I__1426\ : Span4Mux_h
    port map (
            O => \N__6285\,
            I => \N__6257\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__6280\,
            I => \N__6257\
        );

    \I__1424\ : Span4Mux_h
    port map (
            O => \N__6277\,
            I => \N__6257\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__6272\,
            I => \N__6257\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__6269\,
            I => \N__6253\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__6266\,
            I => \N__6250\
        );

    \I__1420\ : Span4Mux_v
    port map (
            O => \N__6257\,
            I => \N__6246\
        );

    \I__1419\ : InMux
    port map (
            O => \N__6256\,
            I => \N__6243\
        );

    \I__1418\ : Span4Mux_s3_h
    port map (
            O => \N__6253\,
            I => \N__6238\
        );

    \I__1417\ : Span4Mux_h
    port map (
            O => \N__6250\,
            I => \N__6238\
        );

    \I__1416\ : InMux
    port map (
            O => \N__6249\,
            I => \N__6235\
        );

    \I__1415\ : Span4Mux_h
    port map (
            O => \N__6246\,
            I => \N__6232\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__6243\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_0\
        );

    \I__1413\ : Odrv4
    port map (
            O => \N__6238\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_0\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__6235\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_0\
        );

    \I__1411\ : Odrv4
    port map (
            O => \N__6232\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_0\
        );

    \I__1410\ : InMux
    port map (
            O => \N__6223\,
            I => \N__6220\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__6220\,
            I => \N__6217\
        );

    \I__1408\ : Odrv4
    port map (
            O => \N__6217\,
            I => \A_c_11\
        );

    \I__1407\ : InMux
    port map (
            O => \N__6214\,
            I => \N__6211\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__6211\,
            I => \U400_SDRAM.MA_5_iv_0_1\
        );

    \I__1405\ : IoInMux
    port map (
            O => \N__6208\,
            I => \N__6205\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__6205\,
            I => \N__6202\
        );

    \I__1403\ : Odrv4
    port map (
            O => \N__6202\,
            I => \MA_c_1\
        );

    \I__1402\ : InMux
    port map (
            O => \N__6199\,
            I => \N__6196\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__6196\,
            I => \N__6193\
        );

    \I__1400\ : Odrv4
    port map (
            O => \N__6193\,
            I => \A_c_15\
        );

    \I__1399\ : InMux
    port map (
            O => \N__6190\,
            I => \N__6187\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__6187\,
            I => \U400_SDRAM.MA_5_iv_0_5\
        );

    \I__1397\ : IoInMux
    port map (
            O => \N__6184\,
            I => \N__6181\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__6181\,
            I => \N__6178\
        );

    \I__1395\ : IoSpan4Mux
    port map (
            O => \N__6178\,
            I => \N__6175\
        );

    \I__1394\ : Span4Mux_s1_v
    port map (
            O => \N__6175\,
            I => \N__6172\
        );

    \I__1393\ : Span4Mux_h
    port map (
            O => \N__6172\,
            I => \N__6169\
        );

    \I__1392\ : Odrv4
    port map (
            O => \N__6169\,
            I => \MA_c_5\
        );

    \I__1391\ : InMux
    port map (
            O => \N__6166\,
            I => \N__6163\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__6163\,
            I => \N__6160\
        );

    \I__1389\ : Span4Mux_s3_v
    port map (
            O => \N__6160\,
            I => \N__6157\
        );

    \I__1388\ : Odrv4
    port map (
            O => \N__6157\,
            I => \A_c_5\
        );

    \I__1387\ : CascadeMux
    port map (
            O => \N__6154\,
            I => \N__6151\
        );

    \I__1386\ : InMux
    port map (
            O => \N__6151\,
            I => \N__6148\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__6148\,
            I => \N__6145\
        );

    \I__1384\ : Span4Mux_v
    port map (
            O => \N__6145\,
            I => \N__6142\
        );

    \I__1383\ : Odrv4
    port map (
            O => \N__6142\,
            I => \A_c_13\
        );

    \I__1382\ : IoInMux
    port map (
            O => \N__6139\,
            I => \N__6136\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__6136\,
            I => \N__6133\
        );

    \I__1380\ : IoSpan4Mux
    port map (
            O => \N__6133\,
            I => \N__6130\
        );

    \I__1379\ : Span4Mux_s3_h
    port map (
            O => \N__6130\,
            I => \N__6127\
        );

    \I__1378\ : Span4Mux_h
    port map (
            O => \N__6127\,
            I => \N__6124\
        );

    \I__1377\ : Odrv4
    port map (
            O => \N__6124\,
            I => \MA_c_3\
        );

    \I__1376\ : InMux
    port map (
            O => \N__6121\,
            I => \N__6118\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__6118\,
            I => \N__6115\
        );

    \I__1374\ : Span4Mux_s2_v
    port map (
            O => \N__6115\,
            I => \N__6112\
        );

    \I__1373\ : IoSpan4Mux
    port map (
            O => \N__6112\,
            I => \N__6109\
        );

    \I__1372\ : Odrv4
    port map (
            O => \N__6109\,
            I => \A_c_4\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__6106\,
            I => \N__6103\
        );

    \I__1370\ : InMux
    port map (
            O => \N__6103\,
            I => \N__6100\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__6100\,
            I => \A_c_12\
        );

    \I__1368\ : IoInMux
    port map (
            O => \N__6097\,
            I => \N__6094\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__6094\,
            I => \MA_c_2\
        );

    \I__1366\ : InMux
    port map (
            O => \N__6091\,
            I => \N__6088\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__6088\,
            I => \N__6085\
        );

    \I__1364\ : Span4Mux_s3_v
    port map (
            O => \N__6085\,
            I => \N__6082\
        );

    \I__1363\ : Odrv4
    port map (
            O => \N__6082\,
            I => \A_c_6\
        );

    \I__1362\ : CascadeMux
    port map (
            O => \N__6079\,
            I => \N__6076\
        );

    \I__1361\ : InMux
    port map (
            O => \N__6076\,
            I => \N__6073\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__6073\,
            I => \N__6070\
        );

    \I__1359\ : Span4Mux_h
    port map (
            O => \N__6070\,
            I => \N__6067\
        );

    \I__1358\ : Odrv4
    port map (
            O => \N__6067\,
            I => \A_c_14\
        );

    \I__1357\ : IoInMux
    port map (
            O => \N__6064\,
            I => \N__6061\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__6061\,
            I => \N__6058\
        );

    \I__1355\ : IoSpan4Mux
    port map (
            O => \N__6058\,
            I => \N__6055\
        );

    \I__1354\ : IoSpan4Mux
    port map (
            O => \N__6055\,
            I => \N__6052\
        );

    \I__1353\ : Odrv4
    port map (
            O => \N__6052\,
            I => \MA_c_4\
        );

    \I__1352\ : InMux
    port map (
            O => \N__6049\,
            I => \N__6046\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__6046\,
            I => \N__6043\
        );

    \I__1350\ : Span4Mux_h
    port map (
            O => \N__6043\,
            I => \N__6040\
        );

    \I__1349\ : Odrv4
    port map (
            O => \N__6040\,
            I => \A_c_2\
        );

    \I__1348\ : CascadeMux
    port map (
            O => \N__6037\,
            I => \N__6028\
        );

    \I__1347\ : InMux
    port map (
            O => \N__6036\,
            I => \N__6020\
        );

    \I__1346\ : InMux
    port map (
            O => \N__6035\,
            I => \N__6017\
        );

    \I__1345\ : InMux
    port map (
            O => \N__6034\,
            I => \N__6012\
        );

    \I__1344\ : InMux
    port map (
            O => \N__6033\,
            I => \N__6012\
        );

    \I__1343\ : InMux
    port map (
            O => \N__6032\,
            I => \N__6007\
        );

    \I__1342\ : InMux
    port map (
            O => \N__6031\,
            I => \N__6007\
        );

    \I__1341\ : InMux
    port map (
            O => \N__6028\,
            I => \N__6001\
        );

    \I__1340\ : InMux
    port map (
            O => \N__6027\,
            I => \N__6001\
        );

    \I__1339\ : InMux
    port map (
            O => \N__6026\,
            I => \N__5996\
        );

    \I__1338\ : InMux
    port map (
            O => \N__6025\,
            I => \N__5996\
        );

    \I__1337\ : InMux
    port map (
            O => \N__6024\,
            I => \N__5989\
        );

    \I__1336\ : InMux
    port map (
            O => \N__6023\,
            I => \N__5989\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__6020\,
            I => \N__5980\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__6017\,
            I => \N__5980\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__6012\,
            I => \N__5980\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__6007\,
            I => \N__5980\
        );

    \I__1331\ : InMux
    port map (
            O => \N__6006\,
            I => \N__5975\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__6001\,
            I => \N__5972\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__5996\,
            I => \N__5969\
        );

    \I__1328\ : InMux
    port map (
            O => \N__5995\,
            I => \N__5966\
        );

    \I__1327\ : InMux
    port map (
            O => \N__5994\,
            I => \N__5962\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__5989\,
            I => \N__5959\
        );

    \I__1325\ : Span4Mux_s3_v
    port map (
            O => \N__5980\,
            I => \N__5956\
        );

    \I__1324\ : InMux
    port map (
            O => \N__5979\,
            I => \N__5953\
        );

    \I__1323\ : InMux
    port map (
            O => \N__5978\,
            I => \N__5950\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__5975\,
            I => \N__5947\
        );

    \I__1321\ : Span4Mux_s3_v
    port map (
            O => \N__5972\,
            I => \N__5942\
        );

    \I__1320\ : Span4Mux_s3_v
    port map (
            O => \N__5969\,
            I => \N__5942\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__5966\,
            I => \N__5938\
        );

    \I__1318\ : InMux
    port map (
            O => \N__5965\,
            I => \N__5935\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__5962\,
            I => \N__5928\
        );

    \I__1316\ : Span4Mux_s3_v
    port map (
            O => \N__5959\,
            I => \N__5928\
        );

    \I__1315\ : Span4Mux_h
    port map (
            O => \N__5956\,
            I => \N__5928\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__5953\,
            I => \N__5925\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__5950\,
            I => \N__5918\
        );

    \I__1312\ : Span4Mux_s3_v
    port map (
            O => \N__5947\,
            I => \N__5918\
        );

    \I__1311\ : Span4Mux_h
    port map (
            O => \N__5942\,
            I => \N__5918\
        );

    \I__1310\ : InMux
    port map (
            O => \N__5941\,
            I => \N__5915\
        );

    \I__1309\ : Span4Mux_v
    port map (
            O => \N__5938\,
            I => \N__5912\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__5935\,
            I => \N__5907\
        );

    \I__1307\ : Span4Mux_v
    port map (
            O => \N__5928\,
            I => \N__5907\
        );

    \I__1306\ : Span4Mux_h
    port map (
            O => \N__5925\,
            I => \N__5902\
        );

    \I__1305\ : Span4Mux_v
    port map (
            O => \N__5918\,
            I => \N__5902\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__5915\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1303\ : Odrv4
    port map (
            O => \N__5912\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1302\ : Odrv4
    port map (
            O => \N__5907\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1301\ : Odrv4
    port map (
            O => \N__5902\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1300\ : InMux
    port map (
            O => \N__5893\,
            I => \N__5889\
        );

    \I__1299\ : InMux
    port map (
            O => \N__5892\,
            I => \N__5883\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__5889\,
            I => \N__5880\
        );

    \I__1297\ : InMux
    port map (
            O => \N__5888\,
            I => \N__5875\
        );

    \I__1296\ : InMux
    port map (
            O => \N__5887\,
            I => \N__5875\
        );

    \I__1295\ : InMux
    port map (
            O => \N__5886\,
            I => \N__5872\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__5883\,
            I => \U400_SDRAM_BURST\
        );

    \I__1293\ : Odrv4
    port map (
            O => \N__5880\,
            I => \U400_SDRAM_BURST\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__5875\,
            I => \U400_SDRAM_BURST\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__5872\,
            I => \U400_SDRAM_BURST\
        );

    \I__1290\ : InMux
    port map (
            O => \N__5863\,
            I => \N__5860\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5860\,
            I => \U400_ADDRESS_DECODE.N_114_0\
        );

    \I__1288\ : InMux
    port map (
            O => \N__5857\,
            I => \N__5853\
        );

    \I__1287\ : InMux
    port map (
            O => \N__5856\,
            I => \N__5848\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__5853\,
            I => \N__5843\
        );

    \I__1285\ : InMux
    port map (
            O => \N__5852\,
            I => \N__5838\
        );

    \I__1284\ : InMux
    port map (
            O => \N__5851\,
            I => \N__5838\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__5848\,
            I => \N__5835\
        );

    \I__1282\ : InMux
    port map (
            O => \N__5847\,
            I => \N__5830\
        );

    \I__1281\ : InMux
    port map (
            O => \N__5846\,
            I => \N__5830\
        );

    \I__1280\ : Span12Mux_s6_h
    port map (
            O => \N__5843\,
            I => \N__5827\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__5838\,
            I => \N__5824\
        );

    \I__1278\ : Span4Mux_h
    port map (
            O => \N__5835\,
            I => \N__5821\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__5830\,
            I => \N__5818\
        );

    \I__1276\ : Odrv12
    port map (
            O => \N__5827\,
            I => \N_65_0\
        );

    \I__1275\ : Odrv4
    port map (
            O => \N__5824\,
            I => \N_65_0\
        );

    \I__1274\ : Odrv4
    port map (
            O => \N__5821\,
            I => \N_65_0\
        );

    \I__1273\ : Odrv4
    port map (
            O => \N__5818\,
            I => \N_65_0\
        );

    \I__1272\ : InMux
    port map (
            O => \N__5809\,
            I => \N__5797\
        );

    \I__1271\ : InMux
    port map (
            O => \N__5808\,
            I => \N__5792\
        );

    \I__1270\ : InMux
    port map (
            O => \N__5807\,
            I => \N__5792\
        );

    \I__1269\ : InMux
    port map (
            O => \N__5806\,
            I => \N__5789\
        );

    \I__1268\ : CascadeMux
    port map (
            O => \N__5805\,
            I => \N__5779\
        );

    \I__1267\ : InMux
    port map (
            O => \N__5804\,
            I => \N__5776\
        );

    \I__1266\ : InMux
    port map (
            O => \N__5803\,
            I => \N__5773\
        );

    \I__1265\ : InMux
    port map (
            O => \N__5802\,
            I => \N__5768\
        );

    \I__1264\ : InMux
    port map (
            O => \N__5801\,
            I => \N__5768\
        );

    \I__1263\ : InMux
    port map (
            O => \N__5800\,
            I => \N__5765\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__5797\,
            I => \N__5758\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__5792\,
            I => \N__5758\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__5789\,
            I => \N__5758\
        );

    \I__1259\ : CascadeMux
    port map (
            O => \N__5788\,
            I => \N__5755\
        );

    \I__1258\ : InMux
    port map (
            O => \N__5787\,
            I => \N__5752\
        );

    \I__1257\ : InMux
    port map (
            O => \N__5786\,
            I => \N__5747\
        );

    \I__1256\ : InMux
    port map (
            O => \N__5785\,
            I => \N__5747\
        );

    \I__1255\ : InMux
    port map (
            O => \N__5784\,
            I => \N__5742\
        );

    \I__1254\ : InMux
    port map (
            O => \N__5783\,
            I => \N__5742\
        );

    \I__1253\ : InMux
    port map (
            O => \N__5782\,
            I => \N__5739\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5779\,
            I => \N__5736\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__5776\,
            I => \N__5733\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__5773\,
            I => \N__5728\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__5768\,
            I => \N__5728\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__5765\,
            I => \N__5720\
        );

    \I__1247\ : Span4Mux_v
    port map (
            O => \N__5758\,
            I => \N__5720\
        );

    \I__1246\ : InMux
    port map (
            O => \N__5755\,
            I => \N__5717\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__5752\,
            I => \N__5714\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__5747\,
            I => \N__5711\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__5742\,
            I => \N__5704\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__5739\,
            I => \N__5704\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__5736\,
            I => \N__5704\
        );

    \I__1240\ : Span4Mux_v
    port map (
            O => \N__5733\,
            I => \N__5699\
        );

    \I__1239\ : Span4Mux_v
    port map (
            O => \N__5728\,
            I => \N__5699\
        );

    \I__1238\ : InMux
    port map (
            O => \N__5727\,
            I => \N__5696\
        );

    \I__1237\ : InMux
    port map (
            O => \N__5726\,
            I => \N__5691\
        );

    \I__1236\ : InMux
    port map (
            O => \N__5725\,
            I => \N__5691\
        );

    \I__1235\ : Span4Mux_h
    port map (
            O => \N__5720\,
            I => \N__5688\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__5717\,
            I => \N__5677\
        );

    \I__1233\ : Span4Mux_v
    port map (
            O => \N__5714\,
            I => \N__5677\
        );

    \I__1232\ : Span4Mux_v
    port map (
            O => \N__5711\,
            I => \N__5677\
        );

    \I__1231\ : Span4Mux_v
    port map (
            O => \N__5704\,
            I => \N__5677\
        );

    \I__1230\ : Span4Mux_h
    port map (
            O => \N__5699\,
            I => \N__5677\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__5696\,
            I => \U400_SDRAM_SDRAM_CONFIGURED\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__5691\,
            I => \U400_SDRAM_SDRAM_CONFIGURED\
        );

    \I__1227\ : Odrv4
    port map (
            O => \N__5688\,
            I => \U400_SDRAM_SDRAM_CONFIGURED\
        );

    \I__1226\ : Odrv4
    port map (
            O => \N__5677\,
            I => \U400_SDRAM_SDRAM_CONFIGURED\
        );

    \I__1225\ : IoInMux
    port map (
            O => \N__5668\,
            I => \N__5665\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__5665\,
            I => \N__5662\
        );

    \I__1223\ : Odrv4
    port map (
            O => \N__5662\,
            I => \N_129_0\
        );

    \I__1222\ : IoInMux
    port map (
            O => \N__5659\,
            I => \N__5656\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__5656\,
            I => \N__5653\
        );

    \I__1220\ : Odrv12
    port map (
            O => \N__5653\,
            I => \N_127_0\
        );

    \I__1219\ : InMux
    port map (
            O => \N__5650\,
            I => \N__5641\
        );

    \I__1218\ : InMux
    port map (
            O => \N__5649\,
            I => \N__5641\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5648\,
            I => \N__5641\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__5641\,
            I => \N__5638\
        );

    \I__1215\ : Span4Mux_v
    port map (
            O => \N__5638\,
            I => \N__5635\
        );

    \I__1214\ : Span4Mux_v
    port map (
            O => \N__5635\,
            I => \N__5631\
        );

    \I__1213\ : InMux
    port map (
            O => \N__5634\,
            I => \N__5628\
        );

    \I__1212\ : Span4Mux_v
    port map (
            O => \N__5631\,
            I => \N__5625\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__5628\,
            I => \N__5622\
        );

    \I__1210\ : Sp12to4
    port map (
            O => \N__5625\,
            I => \N__5617\
        );

    \I__1209\ : Span12Mux_v
    port map (
            O => \N__5622\,
            I => \N__5617\
        );

    \I__1208\ : Odrv12
    port map (
            O => \N__5617\,
            I => \A_c_1\
        );

    \I__1207\ : IoInMux
    port map (
            O => \N__5614\,
            I => \N__5611\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__5611\,
            I => \N__5608\
        );

    \I__1205\ : Odrv4
    port map (
            O => \N__5608\,
            I => \N_128_0\
        );

    \I__1204\ : CascadeMux
    port map (
            O => \N__5605\,
            I => \N__5600\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__5604\,
            I => \N__5597\
        );

    \I__1202\ : InMux
    port map (
            O => \N__5603\,
            I => \N__5593\
        );

    \I__1201\ : InMux
    port map (
            O => \N__5600\,
            I => \N__5586\
        );

    \I__1200\ : InMux
    port map (
            O => \N__5597\,
            I => \N__5586\
        );

    \I__1199\ : InMux
    port map (
            O => \N__5596\,
            I => \N__5586\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__5593\,
            I => \U400_ADDRESS_DECODE.N_122_0\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__5586\,
            I => \U400_ADDRESS_DECODE.N_122_0\
        );

    \I__1196\ : CascadeMux
    port map (
            O => \N__5581\,
            I => \N__5578\
        );

    \I__1195\ : InMux
    port map (
            O => \N__5578\,
            I => \N__5573\
        );

    \I__1194\ : InMux
    port map (
            O => \N__5577\,
            I => \N__5568\
        );

    \I__1193\ : InMux
    port map (
            O => \N__5576\,
            I => \N__5568\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__5573\,
            I => \N__5565\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__5568\,
            I => \N__5561\
        );

    \I__1190\ : Span4Mux_v
    port map (
            O => \N__5565\,
            I => \N__5558\
        );

    \I__1189\ : InMux
    port map (
            O => \N__5564\,
            I => \N__5555\
        );

    \I__1188\ : Span4Mux_v
    port map (
            O => \N__5561\,
            I => \N__5552\
        );

    \I__1187\ : Sp12to4
    port map (
            O => \N__5558\,
            I => \N__5547\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__5555\,
            I => \N__5547\
        );

    \I__1185\ : Odrv4
    port map (
            O => \N__5552\,
            I => \SIZ_c_0\
        );

    \I__1184\ : Odrv12
    port map (
            O => \N__5547\,
            I => \SIZ_c_0\
        );

    \I__1183\ : InMux
    port map (
            O => \N__5542\,
            I => \N__5538\
        );

    \I__1182\ : InMux
    port map (
            O => \N__5541\,
            I => \N__5535\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__5538\,
            I => \N__5531\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__5535\,
            I => \N__5528\
        );

    \I__1179\ : InMux
    port map (
            O => \N__5534\,
            I => \N__5525\
        );

    \I__1178\ : Span4Mux_h
    port map (
            O => \N__5531\,
            I => \N__5520\
        );

    \I__1177\ : Span4Mux_v
    port map (
            O => \N__5528\,
            I => \N__5520\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__5525\,
            I => \N__5517\
        );

    \I__1175\ : Span4Mux_v
    port map (
            O => \N__5520\,
            I => \N__5514\
        );

    \I__1174\ : Sp12to4
    port map (
            O => \N__5517\,
            I => \N__5511\
        );

    \I__1173\ : Span4Mux_v
    port map (
            O => \N__5514\,
            I => \N__5508\
        );

    \I__1172\ : Span12Mux_v
    port map (
            O => \N__5511\,
            I => \N__5505\
        );

    \I__1171\ : Span4Mux_h
    port map (
            O => \N__5508\,
            I => \N__5502\
        );

    \I__1170\ : Odrv12
    port map (
            O => \N__5505\,
            I => \A_c_0\
        );

    \I__1169\ : Odrv4
    port map (
            O => \N__5502\,
            I => \A_c_0\
        );

    \I__1168\ : CascadeMux
    port map (
            O => \N__5497\,
            I => \N__5493\
        );

    \I__1167\ : InMux
    port map (
            O => \N__5496\,
            I => \N__5490\
        );

    \I__1166\ : InMux
    port map (
            O => \N__5493\,
            I => \N__5486\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__5490\,
            I => \N__5483\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5489\,
            I => \N__5480\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__5486\,
            I => \U400_ADDRESS_DECODE.N_4_0\
        );

    \I__1162\ : Odrv12
    port map (
            O => \N__5483\,
            I => \U400_ADDRESS_DECODE.N_4_0\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__5480\,
            I => \U400_ADDRESS_DECODE.N_4_0\
        );

    \I__1160\ : InMux
    port map (
            O => \N__5473\,
            I => \N__5470\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__5470\,
            I => \N__5466\
        );

    \I__1158\ : InMux
    port map (
            O => \N__5469\,
            I => \N__5463\
        );

    \I__1157\ : Span4Mux_v
    port map (
            O => \N__5466\,
            I => \N__5456\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__5463\,
            I => \N__5456\
        );

    \I__1155\ : InMux
    port map (
            O => \N__5462\,
            I => \N__5451\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5461\,
            I => \N__5451\
        );

    \I__1153\ : Span4Mux_v
    port map (
            O => \N__5456\,
            I => \N__5448\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__5451\,
            I => \N__5445\
        );

    \I__1151\ : Span4Mux_h
    port map (
            O => \N__5448\,
            I => \N__5442\
        );

    \I__1150\ : Span4Mux_v
    port map (
            O => \N__5445\,
            I => \N__5439\
        );

    \I__1149\ : Odrv4
    port map (
            O => \N__5442\,
            I => \SIZ_c_1\
        );

    \I__1148\ : Odrv4
    port map (
            O => \N__5439\,
            I => \SIZ_c_1\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5434\,
            I => \N__5428\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5433\,
            I => \N__5428\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__5428\,
            I => \U400_ADDRESS_DECODE.N_186_mux\
        );

    \I__1144\ : InMux
    port map (
            O => \N__5425\,
            I => \N__5422\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__5422\,
            I => \U400_ADDRESS_DECODE.N_146_0\
        );

    \I__1142\ : CascadeMux
    port map (
            O => \N__5419\,
            I => \N__5415\
        );

    \I__1141\ : CascadeMux
    port map (
            O => \N__5418\,
            I => \N__5412\
        );

    \I__1140\ : InMux
    port map (
            O => \N__5415\,
            I => \N__5407\
        );

    \I__1139\ : InMux
    port map (
            O => \N__5412\,
            I => \N__5407\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__5407\,
            I => \N__5404\
        );

    \I__1137\ : Span4Mux_h
    port map (
            O => \N__5404\,
            I => \N__5401\
        );

    \I__1136\ : Span4Mux_v
    port map (
            O => \N__5401\,
            I => \N__5397\
        );

    \I__1135\ : InMux
    port map (
            O => \N__5400\,
            I => \N__5394\
        );

    \I__1134\ : Odrv4
    port map (
            O => \N__5397\,
            I => \N_14_i\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__5394\,
            I => \N_14_i\
        );

    \I__1132\ : CascadeMux
    port map (
            O => \N__5389\,
            I => \U400_ADDRESS_DECODE.N_147_0_cascade_\
        );

    \I__1131\ : InMux
    port map (
            O => \N__5386\,
            I => \N__5383\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__5383\,
            I => \U400_ADDRESS_DECODE.N_136_0\
        );

    \I__1129\ : InMux
    port map (
            O => \N__5380\,
            I => \N__5377\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__5377\,
            I => \N_43\
        );

    \I__1127\ : InMux
    port map (
            O => \N__5374\,
            I => \N__5371\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__5371\,
            I => \N__5368\
        );

    \I__1125\ : Span4Mux_h
    port map (
            O => \N__5368\,
            I => \N__5365\
        );

    \I__1124\ : Sp12to4
    port map (
            O => \N__5365\,
            I => \N__5362\
        );

    \I__1123\ : Span12Mux_v
    port map (
            O => \N__5362\,
            I => \N__5359\
        );

    \I__1122\ : Odrv12
    port map (
            O => \N__5359\,
            I => \A_c_20\
        );

    \I__1121\ : IoInMux
    port map (
            O => \N__5356\,
            I => \N__5353\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__5353\,
            I => \N__5350\
        );

    \I__1119\ : Span4Mux_s0_v
    port map (
            O => \N__5350\,
            I => \N__5347\
        );

    \I__1118\ : Odrv4
    port map (
            O => \N__5347\,
            I => \MA_c_10\
        );

    \I__1117\ : CascadeMux
    port map (
            O => \N__5344\,
            I => \N__5341\
        );

    \I__1116\ : InMux
    port map (
            O => \N__5341\,
            I => \N__5338\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__5338\,
            I => \N__5335\
        );

    \I__1114\ : Span12Mux_s11_v
    port map (
            O => \N__5335\,
            I => \N__5332\
        );

    \I__1113\ : Odrv12
    port map (
            O => \N__5332\,
            I => \A_c_25\
        );

    \I__1112\ : IoInMux
    port map (
            O => \N__5329\,
            I => \N__5326\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__5326\,
            I => \N__5323\
        );

    \I__1110\ : Odrv4
    port map (
            O => \N__5323\,
            I => \MA_c_11\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__5320\,
            I => \U400_ADDRESS_DECODE.N_4_0_cascade_\
        );

    \I__1108\ : IoInMux
    port map (
            O => \N__5317\,
            I => \N__5314\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__5314\,
            I => \N__5311\
        );

    \I__1106\ : Span12Mux_s3_v
    port map (
            O => \N__5311\,
            I => \N__5308\
        );

    \I__1105\ : Odrv12
    port map (
            O => \N__5308\,
            I => \N_124_0\
        );

    \I__1104\ : InMux
    port map (
            O => \N__5305\,
            I => \N__5302\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5302\,
            I => \U400_SDRAM.N_252_0_0\
        );

    \I__1102\ : InMux
    port map (
            O => \N__5299\,
            I => \N__5296\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__5296\,
            I => \U400_SDRAM.N_252_0_0_en\
        );

    \I__1100\ : InMux
    port map (
            O => \N__5293\,
            I => \N__5289\
        );

    \I__1099\ : InMux
    port map (
            O => \N__5292\,
            I => \N__5286\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__5289\,
            I => \N_174\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__5286\,
            I => \N_174\
        );

    \I__1096\ : InMux
    port map (
            O => \N__5281\,
            I => \N__5278\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__5278\,
            I => \U400_SDRAM_TA_OUT_5_0\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5275\,
            I => \N__5272\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__5272\,
            I => \U400_SDRAM_N_252_0\
        );

    \I__1092\ : IoInMux
    port map (
            O => \N__5269\,
            I => \N__5266\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__5266\,
            I => \N__5262\
        );

    \I__1090\ : CascadeMux
    port map (
            O => \N__5265\,
            I => \N__5259\
        );

    \I__1089\ : Span4Mux_s3_h
    port map (
            O => \N__5262\,
            I => \N__5256\
        );

    \I__1088\ : InMux
    port map (
            O => \N__5259\,
            I => \N__5253\
        );

    \I__1087\ : Odrv4
    port map (
            O => \N__5256\,
            I => \TA_OUT\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__5253\,
            I => \TA_OUT\
        );

    \I__1085\ : ClkMux
    port map (
            O => \N__5248\,
            I => \N__5167\
        );

    \I__1084\ : ClkMux
    port map (
            O => \N__5247\,
            I => \N__5167\
        );

    \I__1083\ : ClkMux
    port map (
            O => \N__5246\,
            I => \N__5167\
        );

    \I__1082\ : ClkMux
    port map (
            O => \N__5245\,
            I => \N__5167\
        );

    \I__1081\ : ClkMux
    port map (
            O => \N__5244\,
            I => \N__5167\
        );

    \I__1080\ : ClkMux
    port map (
            O => \N__5243\,
            I => \N__5167\
        );

    \I__1079\ : ClkMux
    port map (
            O => \N__5242\,
            I => \N__5167\
        );

    \I__1078\ : ClkMux
    port map (
            O => \N__5241\,
            I => \N__5167\
        );

    \I__1077\ : ClkMux
    port map (
            O => \N__5240\,
            I => \N__5167\
        );

    \I__1076\ : ClkMux
    port map (
            O => \N__5239\,
            I => \N__5167\
        );

    \I__1075\ : ClkMux
    port map (
            O => \N__5238\,
            I => \N__5167\
        );

    \I__1074\ : ClkMux
    port map (
            O => \N__5237\,
            I => \N__5167\
        );

    \I__1073\ : ClkMux
    port map (
            O => \N__5236\,
            I => \N__5167\
        );

    \I__1072\ : ClkMux
    port map (
            O => \N__5235\,
            I => \N__5167\
        );

    \I__1071\ : ClkMux
    port map (
            O => \N__5234\,
            I => \N__5167\
        );

    \I__1070\ : ClkMux
    port map (
            O => \N__5233\,
            I => \N__5167\
        );

    \I__1069\ : ClkMux
    port map (
            O => \N__5232\,
            I => \N__5167\
        );

    \I__1068\ : ClkMux
    port map (
            O => \N__5231\,
            I => \N__5167\
        );

    \I__1067\ : ClkMux
    port map (
            O => \N__5230\,
            I => \N__5167\
        );

    \I__1066\ : ClkMux
    port map (
            O => \N__5229\,
            I => \N__5167\
        );

    \I__1065\ : ClkMux
    port map (
            O => \N__5228\,
            I => \N__5167\
        );

    \I__1064\ : ClkMux
    port map (
            O => \N__5227\,
            I => \N__5167\
        );

    \I__1063\ : ClkMux
    port map (
            O => \N__5226\,
            I => \N__5167\
        );

    \I__1062\ : ClkMux
    port map (
            O => \N__5225\,
            I => \N__5167\
        );

    \I__1061\ : ClkMux
    port map (
            O => \N__5224\,
            I => \N__5167\
        );

    \I__1060\ : ClkMux
    port map (
            O => \N__5223\,
            I => \N__5167\
        );

    \I__1059\ : ClkMux
    port map (
            O => \N__5222\,
            I => \N__5167\
        );

    \I__1058\ : GlobalMux
    port map (
            O => \N__5167\,
            I => \N__5164\
        );

    \I__1057\ : gio2CtrlBuf
    port map (
            O => \N__5164\,
            I => \CLK40_c_g\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5161\,
            I => \N__5155\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5160\,
            I => \N__5155\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__5155\,
            I => \U400_SDRAM_TA_COUNTER_5\
        );

    \I__1053\ : CascadeMux
    port map (
            O => \N__5152\,
            I => \U400_SDRAM.N_252_0_0_cascade_\
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__5149\,
            I => \N__5145\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5148\,
            I => \N__5137\
        );

    \I__1050\ : InMux
    port map (
            O => \N__5145\,
            I => \N__5137\
        );

    \I__1049\ : InMux
    port map (
            O => \N__5144\,
            I => \N__5137\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__5137\,
            I => \U400_SDRAM_TA_COUNTER_2\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5134\,
            I => \N__5130\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5133\,
            I => \N__5127\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__5130\,
            I => \U400_SDRAM_TA_COUNTER_3\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__5127\,
            I => \U400_SDRAM_TA_COUNTER_3\
        );

    \I__1043\ : CascadeMux
    port map (
            O => \N__5122\,
            I => \N__5119\
        );

    \I__1042\ : InMux
    port map (
            O => \N__5119\,
            I => \N__5116\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__5116\,
            I => \N__5113\
        );

    \I__1040\ : Span4Mux_v
    port map (
            O => \N__5113\,
            I => \N__5110\
        );

    \I__1039\ : Span4Mux_h
    port map (
            O => \N__5110\,
            I => \N__5107\
        );

    \I__1038\ : Odrv4
    port map (
            O => \N__5107\,
            I => \A_c_22\
        );

    \I__1037\ : IoInMux
    port map (
            O => \N__5104\,
            I => \N__5101\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__5101\,
            I => \N__5098\
        );

    \I__1035\ : Span4Mux_s2_h
    port map (
            O => \N__5098\,
            I => \N__5095\
        );

    \I__1034\ : Span4Mux_h
    port map (
            O => \N__5095\,
            I => \N__5092\
        );

    \I__1033\ : Span4Mux_v
    port map (
            O => \N__5092\,
            I => \N__5088\
        );

    \I__1032\ : InMux
    port map (
            O => \N__5091\,
            I => \N__5085\
        );

    \I__1031\ : Odrv4
    port map (
            O => \N__5088\,
            I => \BANK1_c\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__5085\,
            I => \BANK1_c\
        );

    \I__1029\ : CascadeMux
    port map (
            O => \N__5080\,
            I => \N__5077\
        );

    \I__1028\ : InMux
    port map (
            O => \N__5077\,
            I => \N__5074\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__5074\,
            I => \N__5071\
        );

    \I__1026\ : Span4Mux_v
    port map (
            O => \N__5071\,
            I => \N__5068\
        );

    \I__1025\ : Sp12to4
    port map (
            O => \N__5068\,
            I => \N__5065\
        );

    \I__1024\ : Odrv12
    port map (
            O => \N__5065\,
            I => \A_c_21\
        );

    \I__1023\ : InMux
    port map (
            O => \N__5062\,
            I => \N__5056\
        );

    \I__1022\ : InMux
    port map (
            O => \N__5061\,
            I => \N__5056\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__5056\,
            I => \U400_SDRAM_un1_SDRAM_COUNTER59_2_0\
        );

    \I__1020\ : IoInMux
    port map (
            O => \N__5053\,
            I => \N__5050\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__5050\,
            I => \N__5047\
        );

    \I__1018\ : Span4Mux_s2_h
    port map (
            O => \N__5047\,
            I => \N__5044\
        );

    \I__1017\ : Span4Mux_h
    port map (
            O => \N__5044\,
            I => \N__5041\
        );

    \I__1016\ : Span4Mux_v
    port map (
            O => \N__5041\,
            I => \N__5037\
        );

    \I__1015\ : InMux
    port map (
            O => \N__5040\,
            I => \N__5034\
        );

    \I__1014\ : Odrv4
    port map (
            O => \N__5037\,
            I => \BANK0_c\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__5034\,
            I => \BANK0_c\
        );

    \I__1012\ : InMux
    port map (
            O => \N__5029\,
            I => \N__5026\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__5026\,
            I => \N__5022\
        );

    \I__1010\ : InMux
    port map (
            O => \N__5025\,
            I => \N__5019\
        );

    \I__1009\ : Odrv4
    port map (
            O => \N__5022\,
            I => \U400_SDRAM_SDRAM_CMD_1_sqmuxa_1\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__5019\,
            I => \U400_SDRAM_SDRAM_CMD_1_sqmuxa_1\
        );

    \I__1007\ : InMux
    port map (
            O => \N__5014\,
            I => \N__5007\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5013\,
            I => \N__5004\
        );

    \I__1005\ : CascadeMux
    port map (
            O => \N__5012\,
            I => \N__4997\
        );

    \I__1004\ : CascadeMux
    port map (
            O => \N__5011\,
            I => \N__4993\
        );

    \I__1003\ : CascadeMux
    port map (
            O => \N__5010\,
            I => \N__4990\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__5007\,
            I => \N__4978\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__5004\,
            I => \N__4978\
        );

    \I__1000\ : InMux
    port map (
            O => \N__5003\,
            I => \N__4975\
        );

    \I__999\ : InMux
    port map (
            O => \N__5002\,
            I => \N__4972\
        );

    \I__998\ : InMux
    port map (
            O => \N__5001\,
            I => \N__4967\
        );

    \I__997\ : InMux
    port map (
            O => \N__5000\,
            I => \N__4967\
        );

    \I__996\ : InMux
    port map (
            O => \N__4997\,
            I => \N__4962\
        );

    \I__995\ : InMux
    port map (
            O => \N__4996\,
            I => \N__4962\
        );

    \I__994\ : InMux
    port map (
            O => \N__4993\,
            I => \N__4959\
        );

    \I__993\ : InMux
    port map (
            O => \N__4990\,
            I => \N__4954\
        );

    \I__992\ : InMux
    port map (
            O => \N__4989\,
            I => \N__4954\
        );

    \I__991\ : CascadeMux
    port map (
            O => \N__4988\,
            I => \N__4950\
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__4987\,
            I => \N__4944\
        );

    \I__989\ : InMux
    port map (
            O => \N__4986\,
            I => \N__4939\
        );

    \I__988\ : InMux
    port map (
            O => \N__4985\,
            I => \N__4939\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__4984\,
            I => \N__4936\
        );

    \I__986\ : InMux
    port map (
            O => \N__4983\,
            I => \N__4933\
        );

    \I__985\ : Span4Mux_h
    port map (
            O => \N__4978\,
            I => \N__4924\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__4975\,
            I => \N__4924\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__4972\,
            I => \N__4924\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__4967\,
            I => \N__4924\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__4962\,
            I => \N__4919\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__4959\,
            I => \N__4914\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__4954\,
            I => \N__4914\
        );

    \I__978\ : InMux
    port map (
            O => \N__4953\,
            I => \N__4909\
        );

    \I__977\ : InMux
    port map (
            O => \N__4950\,
            I => \N__4909\
        );

    \I__976\ : InMux
    port map (
            O => \N__4949\,
            I => \N__4904\
        );

    \I__975\ : InMux
    port map (
            O => \N__4948\,
            I => \N__4904\
        );

    \I__974\ : InMux
    port map (
            O => \N__4947\,
            I => \N__4899\
        );

    \I__973\ : InMux
    port map (
            O => \N__4944\,
            I => \N__4899\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__4939\,
            I => \N__4896\
        );

    \I__971\ : InMux
    port map (
            O => \N__4936\,
            I => \N__4893\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__4933\,
            I => \N__4888\
        );

    \I__969\ : Span4Mux_v
    port map (
            O => \N__4924\,
            I => \N__4888\
        );

    \I__968\ : InMux
    port map (
            O => \N__4923\,
            I => \N__4885\
        );

    \I__967\ : InMux
    port map (
            O => \N__4922\,
            I => \N__4882\
        );

    \I__966\ : Span4Mux_h
    port map (
            O => \N__4919\,
            I => \N__4871\
        );

    \I__965\ : Span4Mux_h
    port map (
            O => \N__4914\,
            I => \N__4871\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__4909\,
            I => \N__4871\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__4904\,
            I => \N__4871\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__4899\,
            I => \N__4871\
        );

    \I__961\ : Odrv12
    port map (
            O => \N__4896\,
            I => \U400_SDRAM_SDRAM_COUNTER_2\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4893\,
            I => \U400_SDRAM_SDRAM_COUNTER_2\
        );

    \I__959\ : Odrv4
    port map (
            O => \N__4888\,
            I => \U400_SDRAM_SDRAM_COUNTER_2\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__4885\,
            I => \U400_SDRAM_SDRAM_COUNTER_2\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__4882\,
            I => \U400_SDRAM_SDRAM_COUNTER_2\
        );

    \I__956\ : Odrv4
    port map (
            O => \N__4871\,
            I => \U400_SDRAM_SDRAM_COUNTER_2\
        );

    \I__955\ : InMux
    port map (
            O => \N__4858\,
            I => \N__4850\
        );

    \I__954\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4844\
        );

    \I__953\ : InMux
    port map (
            O => \N__4856\,
            I => \N__4837\
        );

    \I__952\ : InMux
    port map (
            O => \N__4855\,
            I => \N__4837\
        );

    \I__951\ : InMux
    port map (
            O => \N__4854\,
            I => \N__4837\
        );

    \I__950\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4834\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__4850\,
            I => \N__4828\
        );

    \I__948\ : InMux
    port map (
            O => \N__4849\,
            I => \N__4821\
        );

    \I__947\ : InMux
    port map (
            O => \N__4848\,
            I => \N__4821\
        );

    \I__946\ : InMux
    port map (
            O => \N__4847\,
            I => \N__4821\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4844\,
            I => \N__4815\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4837\,
            I => \N__4810\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__4834\,
            I => \N__4810\
        );

    \I__942\ : InMux
    port map (
            O => \N__4833\,
            I => \N__4807\
        );

    \I__941\ : InMux
    port map (
            O => \N__4832\,
            I => \N__4802\
        );

    \I__940\ : InMux
    port map (
            O => \N__4831\,
            I => \N__4802\
        );

    \I__939\ : Span4Mux_v
    port map (
            O => \N__4828\,
            I => \N__4792\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4821\,
            I => \N__4789\
        );

    \I__937\ : InMux
    port map (
            O => \N__4820\,
            I => \N__4786\
        );

    \I__936\ : InMux
    port map (
            O => \N__4819\,
            I => \N__4781\
        );

    \I__935\ : InMux
    port map (
            O => \N__4818\,
            I => \N__4781\
        );

    \I__934\ : Span4Mux_h
    port map (
            O => \N__4815\,
            I => \N__4772\
        );

    \I__933\ : Span4Mux_v
    port map (
            O => \N__4810\,
            I => \N__4772\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4807\,
            I => \N__4772\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4802\,
            I => \N__4772\
        );

    \I__930\ : InMux
    port map (
            O => \N__4801\,
            I => \N__4767\
        );

    \I__929\ : InMux
    port map (
            O => \N__4800\,
            I => \N__4767\
        );

    \I__928\ : InMux
    port map (
            O => \N__4799\,
            I => \N__4762\
        );

    \I__927\ : InMux
    port map (
            O => \N__4798\,
            I => \N__4762\
        );

    \I__926\ : InMux
    port map (
            O => \N__4797\,
            I => \N__4755\
        );

    \I__925\ : InMux
    port map (
            O => \N__4796\,
            I => \N__4755\
        );

    \I__924\ : InMux
    port map (
            O => \N__4795\,
            I => \N__4755\
        );

    \I__923\ : Odrv4
    port map (
            O => \N__4792\,
            I => \N_60\
        );

    \I__922\ : Odrv4
    port map (
            O => \N__4789\,
            I => \N_60\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4786\,
            I => \N_60\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4781\,
            I => \N_60\
        );

    \I__919\ : Odrv4
    port map (
            O => \N__4772\,
            I => \N_60\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__4767\,
            I => \N_60\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__4762\,
            I => \N_60\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4755\,
            I => \N_60\
        );

    \I__915\ : InMux
    port map (
            O => \N__4738\,
            I => \N__4735\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4735\,
            I => \U400_ADDRESS_DECODE.m145_nsZ0Z_1\
        );

    \I__913\ : InMux
    port map (
            O => \N__4732\,
            I => \N__4728\
        );

    \I__912\ : InMux
    port map (
            O => \N__4731\,
            I => \N__4725\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__4728\,
            I => \N__4716\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__4725\,
            I => \N__4713\
        );

    \I__909\ : InMux
    port map (
            O => \N__4724\,
            I => \N__4708\
        );

    \I__908\ : InMux
    port map (
            O => \N__4723\,
            I => \N__4708\
        );

    \I__907\ : InMux
    port map (
            O => \N__4722\,
            I => \N__4699\
        );

    \I__906\ : InMux
    port map (
            O => \N__4721\,
            I => \N__4699\
        );

    \I__905\ : InMux
    port map (
            O => \N__4720\,
            I => \N__4699\
        );

    \I__904\ : InMux
    port map (
            O => \N__4719\,
            I => \N__4699\
        );

    \I__903\ : Span4Mux_h
    port map (
            O => \N__4716\,
            I => \N__4696\
        );

    \I__902\ : Odrv4
    port map (
            O => \N__4713\,
            I => \N_100_0_i\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4708\,
            I => \N_100_0_i\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__4699\,
            I => \N_100_0_i\
        );

    \I__899\ : Odrv4
    port map (
            O => \N__4696\,
            I => \N_100_0_i\
        );

    \I__898\ : IoInMux
    port map (
            O => \N__4687\,
            I => \N__4684\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__4684\,
            I => \N__4681\
        );

    \I__896\ : IoSpan4Mux
    port map (
            O => \N__4681\,
            I => \N__4678\
        );

    \I__895\ : Span4Mux_s1_h
    port map (
            O => \N__4678\,
            I => \N__4674\
        );

    \I__894\ : CascadeMux
    port map (
            O => \N__4677\,
            I => \N__4671\
        );

    \I__893\ : Span4Mux_h
    port map (
            O => \N__4674\,
            I => \N__4668\
        );

    \I__892\ : InMux
    port map (
            O => \N__4671\,
            I => \N__4665\
        );

    \I__891\ : Odrv4
    port map (
            O => \N__4668\,
            I => \CONSTANT_ONE_NET\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__4665\,
            I => \CONSTANT_ONE_NET\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__4660\,
            I => \N__4649\
        );

    \I__888\ : CascadeMux
    port map (
            O => \N__4659\,
            I => \N__4641\
        );

    \I__887\ : InMux
    port map (
            O => \N__4658\,
            I => \N__4638\
        );

    \I__886\ : InMux
    port map (
            O => \N__4657\,
            I => \N__4635\
        );

    \I__885\ : CascadeMux
    port map (
            O => \N__4656\,
            I => \N__4632\
        );

    \I__884\ : InMux
    port map (
            O => \N__4655\,
            I => \N__4627\
        );

    \I__883\ : InMux
    port map (
            O => \N__4654\,
            I => \N__4624\
        );

    \I__882\ : InMux
    port map (
            O => \N__4653\,
            I => \N__4619\
        );

    \I__881\ : InMux
    port map (
            O => \N__4652\,
            I => \N__4619\
        );

    \I__880\ : InMux
    port map (
            O => \N__4649\,
            I => \N__4612\
        );

    \I__879\ : InMux
    port map (
            O => \N__4648\,
            I => \N__4612\
        );

    \I__878\ : InMux
    port map (
            O => \N__4647\,
            I => \N__4612\
        );

    \I__877\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4609\
        );

    \I__876\ : CascadeMux
    port map (
            O => \N__4645\,
            I => \N__4604\
        );

    \I__875\ : InMux
    port map (
            O => \N__4644\,
            I => \N__4593\
        );

    \I__874\ : InMux
    port map (
            O => \N__4641\,
            I => \N__4593\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__4638\,
            I => \N__4588\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4635\,
            I => \N__4588\
        );

    \I__871\ : InMux
    port map (
            O => \N__4632\,
            I => \N__4581\
        );

    \I__870\ : InMux
    port map (
            O => \N__4631\,
            I => \N__4581\
        );

    \I__869\ : InMux
    port map (
            O => \N__4630\,
            I => \N__4581\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4627\,
            I => \N__4576\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4624\,
            I => \N__4576\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__4619\,
            I => \N__4571\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__4612\,
            I => \N__4571\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4609\,
            I => \N__4568\
        );

    \I__863\ : InMux
    port map (
            O => \N__4608\,
            I => \N__4563\
        );

    \I__862\ : InMux
    port map (
            O => \N__4607\,
            I => \N__4563\
        );

    \I__861\ : InMux
    port map (
            O => \N__4604\,
            I => \N__4560\
        );

    \I__860\ : InMux
    port map (
            O => \N__4603\,
            I => \N__4553\
        );

    \I__859\ : InMux
    port map (
            O => \N__4602\,
            I => \N__4553\
        );

    \I__858\ : InMux
    port map (
            O => \N__4601\,
            I => \N__4553\
        );

    \I__857\ : InMux
    port map (
            O => \N__4600\,
            I => \N__4550\
        );

    \I__856\ : InMux
    port map (
            O => \N__4599\,
            I => \N__4547\
        );

    \I__855\ : InMux
    port map (
            O => \N__4598\,
            I => \N__4544\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__4593\,
            I => \N__4539\
        );

    \I__853\ : Span4Mux_v
    port map (
            O => \N__4588\,
            I => \N__4539\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__4581\,
            I => \N__4534\
        );

    \I__851\ : Span4Mux_h
    port map (
            O => \N__4576\,
            I => \N__4534\
        );

    \I__850\ : Span4Mux_h
    port map (
            O => \N__4571\,
            I => \N__4531\
        );

    \I__849\ : Span4Mux_h
    port map (
            O => \N__4568\,
            I => \N__4522\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__4563\,
            I => \N__4522\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4560\,
            I => \N__4522\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4553\,
            I => \N__4522\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__4550\,
            I => \U400_SDRAM_SDRAM_COUNTER_0\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__4547\,
            I => \U400_SDRAM_SDRAM_COUNTER_0\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__4544\,
            I => \U400_SDRAM_SDRAM_COUNTER_0\
        );

    \I__842\ : Odrv4
    port map (
            O => \N__4539\,
            I => \U400_SDRAM_SDRAM_COUNTER_0\
        );

    \I__841\ : Odrv4
    port map (
            O => \N__4534\,
            I => \U400_SDRAM_SDRAM_COUNTER_0\
        );

    \I__840\ : Odrv4
    port map (
            O => \N__4531\,
            I => \U400_SDRAM_SDRAM_COUNTER_0\
        );

    \I__839\ : Odrv4
    port map (
            O => \N__4522\,
            I => \U400_SDRAM_SDRAM_COUNTER_0\
        );

    \I__838\ : CEMux
    port map (
            O => \N__4507\,
            I => \N__4504\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4504\,
            I => \N__4499\
        );

    \I__836\ : CEMux
    port map (
            O => \N__4503\,
            I => \N__4496\
        );

    \I__835\ : CEMux
    port map (
            O => \N__4502\,
            I => \N__4493\
        );

    \I__834\ : Span4Mux_h
    port map (
            O => \N__4499\,
            I => \N__4490\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__4496\,
            I => \N__4487\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4493\,
            I => \N__4484\
        );

    \I__831\ : Odrv4
    port map (
            O => \N__4490\,
            I => \U400_SDRAM_SDRAM_COUNTERe_0_i\
        );

    \I__830\ : Odrv4
    port map (
            O => \N__4487\,
            I => \U400_SDRAM_SDRAM_COUNTERe_0_i\
        );

    \I__829\ : Odrv4
    port map (
            O => \N__4484\,
            I => \U400_SDRAM_SDRAM_COUNTERe_0_i\
        );

    \I__828\ : InMux
    port map (
            O => \N__4477\,
            I => \N__4472\
        );

    \I__827\ : InMux
    port map (
            O => \N__4476\,
            I => \N__4467\
        );

    \I__826\ : InMux
    port map (
            O => \N__4475\,
            I => \N__4467\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__4472\,
            I => \N__4464\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__4467\,
            I => \N__4461\
        );

    \I__823\ : Span4Mux_v
    port map (
            O => \N__4464\,
            I => \N__4458\
        );

    \I__822\ : Odrv12
    port map (
            O => \N__4461\,
            I => \U400_ADDRESS_DECODE.N_135_0\
        );

    \I__821\ : Odrv4
    port map (
            O => \N__4458\,
            I => \U400_ADDRESS_DECODE.N_135_0\
        );

    \I__820\ : CascadeMux
    port map (
            O => \N__4453\,
            I => \N__4449\
        );

    \I__819\ : InMux
    port map (
            O => \N__4452\,
            I => \N__4441\
        );

    \I__818\ : InMux
    port map (
            O => \N__4449\,
            I => \N__4441\
        );

    \I__817\ : InMux
    port map (
            O => \N__4448\,
            I => \N__4441\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__4441\,
            I => \U400_SDRAM_TA_COUNTER_4\
        );

    \I__815\ : InMux
    port map (
            O => \N__4438\,
            I => \N__4433\
        );

    \I__814\ : InMux
    port map (
            O => \N__4437\,
            I => \N__4428\
        );

    \I__813\ : InMux
    port map (
            O => \N__4436\,
            I => \N__4428\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__4433\,
            I => \U400_SDRAM_TA_COUNTER_1\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__4428\,
            I => \U400_SDRAM_TA_COUNTER_1\
        );

    \I__810\ : CascadeMux
    port map (
            O => \N__4423\,
            I => \U400_ADDRESS_DECODE.N_177_mux_cascade_\
        );

    \I__809\ : CascadeMux
    port map (
            O => \N__4420\,
            I => \N__4416\
        );

    \I__808\ : CascadeMux
    port map (
            O => \N__4419\,
            I => \N__4413\
        );

    \I__807\ : InMux
    port map (
            O => \N__4416\,
            I => \N__4405\
        );

    \I__806\ : InMux
    port map (
            O => \N__4413\,
            I => \N__4405\
        );

    \I__805\ : InMux
    port map (
            O => \N__4412\,
            I => \N__4405\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__4405\,
            I => \U400_SDRAM_TA_COUNTER_0\
        );

    \I__803\ : InMux
    port map (
            O => \N__4402\,
            I => \N__4389\
        );

    \I__802\ : InMux
    port map (
            O => \N__4401\,
            I => \N__4389\
        );

    \I__801\ : InMux
    port map (
            O => \N__4400\,
            I => \N__4389\
        );

    \I__800\ : InMux
    port map (
            O => \N__4399\,
            I => \N__4389\
        );

    \I__799\ : InMux
    port map (
            O => \N__4398\,
            I => \N__4386\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4389\,
            I => \N__4383\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__4386\,
            I => \U400_SDRAM_TACK\
        );

    \I__796\ : Odrv4
    port map (
            O => \N__4383\,
            I => \U400_SDRAM_TACK\
        );

    \I__795\ : InMux
    port map (
            O => \N__4378\,
            I => \N__4375\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__4375\,
            I => \N__4372\
        );

    \I__793\ : Span12Mux_v
    port map (
            O => \N__4372\,
            I => \N__4369\
        );

    \I__792\ : Odrv12
    port map (
            O => \N__4369\,
            I => \RnW_c\
        );

    \I__791\ : CascadeMux
    port map (
            O => \N__4366\,
            I => \N__4359\
        );

    \I__790\ : CascadeMux
    port map (
            O => \N__4365\,
            I => \N__4356\
        );

    \I__789\ : CascadeMux
    port map (
            O => \N__4364\,
            I => \N__4352\
        );

    \I__788\ : CascadeMux
    port map (
            O => \N__4363\,
            I => \N__4349\
        );

    \I__787\ : InMux
    port map (
            O => \N__4362\,
            I => \N__4344\
        );

    \I__786\ : InMux
    port map (
            O => \N__4359\,
            I => \N__4341\
        );

    \I__785\ : InMux
    port map (
            O => \N__4356\,
            I => \N__4338\
        );

    \I__784\ : InMux
    port map (
            O => \N__4355\,
            I => \N__4335\
        );

    \I__783\ : InMux
    port map (
            O => \N__4352\,
            I => \N__4330\
        );

    \I__782\ : InMux
    port map (
            O => \N__4349\,
            I => \N__4330\
        );

    \I__781\ : InMux
    port map (
            O => \N__4348\,
            I => \N__4326\
        );

    \I__780\ : CascadeMux
    port map (
            O => \N__4347\,
            I => \N__4322\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__4344\,
            I => \N__4317\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__4341\,
            I => \N__4317\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__4338\,
            I => \N__4310\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__4335\,
            I => \N__4310\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__4330\,
            I => \N__4310\
        );

    \I__774\ : InMux
    port map (
            O => \N__4329\,
            I => \N__4307\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__4326\,
            I => \N__4304\
        );

    \I__772\ : InMux
    port map (
            O => \N__4325\,
            I => \N__4299\
        );

    \I__771\ : InMux
    port map (
            O => \N__4322\,
            I => \N__4299\
        );

    \I__770\ : Span4Mux_h
    port map (
            O => \N__4317\,
            I => \N__4296\
        );

    \I__769\ : Span4Mux_v
    port map (
            O => \N__4310\,
            I => \N__4293\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__4307\,
            I => \U400_SDRAM_WRITE_CYCLE\
        );

    \I__767\ : Odrv4
    port map (
            O => \N__4304\,
            I => \U400_SDRAM_WRITE_CYCLE\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__4299\,
            I => \U400_SDRAM_WRITE_CYCLE\
        );

    \I__765\ : Odrv4
    port map (
            O => \N__4296\,
            I => \U400_SDRAM_WRITE_CYCLE\
        );

    \I__764\ : Odrv4
    port map (
            O => \N__4293\,
            I => \U400_SDRAM_WRITE_CYCLE\
        );

    \I__763\ : InMux
    port map (
            O => \N__4282\,
            I => \N__4279\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__4279\,
            I => \N_48\
        );

    \I__761\ : InMux
    port map (
            O => \N__4276\,
            I => \N__4273\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__4273\,
            I => \N_142_0\
        );

    \I__759\ : InMux
    port map (
            O => \N__4270\,
            I => \N__4267\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__4267\,
            I => \N__4263\
        );

    \I__757\ : InMux
    port map (
            O => \N__4266\,
            I => \N__4260\
        );

    \I__756\ : Odrv12
    port map (
            O => \N__4263\,
            I => \U400_ADDRESS_DECODE.N_12_0\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__4260\,
            I => \U400_ADDRESS_DECODE.N_12_0\
        );

    \I__754\ : InMux
    port map (
            O => \N__4255\,
            I => \N__4252\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__4252\,
            I => \N__4249\
        );

    \I__752\ : Odrv4
    port map (
            O => \N__4249\,
            I => \U400_ADDRESS_DECODE.N_21_0\
        );

    \I__751\ : CascadeMux
    port map (
            O => \N__4246\,
            I => \N__4242\
        );

    \I__750\ : CascadeMux
    port map (
            O => \N__4245\,
            I => \N__4239\
        );

    \I__749\ : InMux
    port map (
            O => \N__4242\,
            I => \N__4234\
        );

    \I__748\ : InMux
    port map (
            O => \N__4239\,
            I => \N__4234\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__4234\,
            I => \N__4231\
        );

    \I__746\ : Odrv12
    port map (
            O => \N__4231\,
            I => \A_c_23\
        );

    \I__745\ : InMux
    port map (
            O => \N__4228\,
            I => \N__4225\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__4225\,
            I => \N_137_0\
        );

    \I__743\ : InMux
    port map (
            O => \N__4222\,
            I => \N__4219\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__4219\,
            I => \N__4215\
        );

    \I__741\ : InMux
    port map (
            O => \N__4218\,
            I => \N__4212\
        );

    \I__740\ : Odrv4
    port map (
            O => \N__4215\,
            I => \N_190_mux\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__4212\,
            I => \N_190_mux\
        );

    \I__738\ : InMux
    port map (
            O => \N__4207\,
            I => \N__4204\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__4204\,
            I => \N_138_0\
        );

    \I__736\ : InMux
    port map (
            O => \N__4201\,
            I => \N__4197\
        );

    \I__735\ : InMux
    port map (
            O => \N__4200\,
            I => \N__4194\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__4197\,
            I => \N_23_0\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__4194\,
            I => \N_23_0\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__4189\,
            I => \N__4185\
        );

    \I__731\ : CascadeMux
    port map (
            O => \N__4188\,
            I => \N__4182\
        );

    \I__730\ : InMux
    port map (
            O => \N__4185\,
            I => \N__4177\
        );

    \I__729\ : InMux
    port map (
            O => \N__4182\,
            I => \N__4177\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__4177\,
            I => \U400_SDRAM.CS1_ENZ0\
        );

    \I__727\ : IoInMux
    port map (
            O => \N__4174\,
            I => \N__4171\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__4171\,
            I => \N__4168\
        );

    \I__725\ : Odrv12
    port map (
            O => \N__4168\,
            I => \CS1n_c\
        );

    \I__724\ : InMux
    port map (
            O => \N__4165\,
            I => \N__4162\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__4162\,
            I => \U400_ADDRESS_DECODE.m94_amZ0Z_1\
        );

    \I__722\ : CascadeMux
    port map (
            O => \N__4159\,
            I => \U400_ADDRESS_DECODE.m94_amZ0_cascade_\
        );

    \I__721\ : InMux
    port map (
            O => \N__4156\,
            I => \N__4153\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__4153\,
            I => \U400_ADDRESS_DECODE.N_95_0\
        );

    \I__719\ : InMux
    port map (
            O => \N__4150\,
            I => \N__4141\
        );

    \I__718\ : InMux
    port map (
            O => \N__4149\,
            I => \N__4136\
        );

    \I__717\ : InMux
    port map (
            O => \N__4148\,
            I => \N__4136\
        );

    \I__716\ : InMux
    port map (
            O => \N__4147\,
            I => \N__4131\
        );

    \I__715\ : InMux
    port map (
            O => \N__4146\,
            I => \N__4131\
        );

    \I__714\ : InMux
    port map (
            O => \N__4145\,
            I => \N__4126\
        );

    \I__713\ : InMux
    port map (
            O => \N__4144\,
            I => \N__4126\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__4141\,
            I => \U400_SDRAM_RAM_CYCLE_START\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__4136\,
            I => \U400_SDRAM_RAM_CYCLE_START\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__4131\,
            I => \U400_SDRAM_RAM_CYCLE_START\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__4126\,
            I => \U400_SDRAM_RAM_CYCLE_START\
        );

    \I__708\ : InMux
    port map (
            O => \N__4117\,
            I => \N__4112\
        );

    \I__707\ : InMux
    port map (
            O => \N__4116\,
            I => \N__4107\
        );

    \I__706\ : InMux
    port map (
            O => \N__4115\,
            I => \N__4107\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__4112\,
            I => \U400_ADDRESS_DECODE.N_15_0\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__4107\,
            I => \U400_ADDRESS_DECODE.N_15_0\
        );

    \I__703\ : CascadeMux
    port map (
            O => \N__4102\,
            I => \N__4097\
        );

    \I__702\ : CascadeMux
    port map (
            O => \N__4101\,
            I => \N__4094\
        );

    \I__701\ : InMux
    port map (
            O => \N__4100\,
            I => \N__4091\
        );

    \I__700\ : InMux
    port map (
            O => \N__4097\,
            I => \N__4088\
        );

    \I__699\ : InMux
    port map (
            O => \N__4094\,
            I => \N__4085\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__4091\,
            I => \N_13_0\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__4088\,
            I => \N_13_0\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__4085\,
            I => \N_13_0\
        );

    \I__695\ : CascadeMux
    port map (
            O => \N__4078\,
            I => \N__4072\
        );

    \I__694\ : InMux
    port map (
            O => \N__4077\,
            I => \N__4068\
        );

    \I__693\ : InMux
    port map (
            O => \N__4076\,
            I => \N__4065\
        );

    \I__692\ : InMux
    port map (
            O => \N__4075\,
            I => \N__4062\
        );

    \I__691\ : InMux
    port map (
            O => \N__4072\,
            I => \N__4056\
        );

    \I__690\ : InMux
    port map (
            O => \N__4071\,
            I => \N__4056\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__4068\,
            I => \N__4050\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__4065\,
            I => \N__4050\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__4062\,
            I => \N__4047\
        );

    \I__686\ : InMux
    port map (
            O => \N__4061\,
            I => \N__4044\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__4056\,
            I => \N__4041\
        );

    \I__684\ : InMux
    port map (
            O => \N__4055\,
            I => \N__4038\
        );

    \I__683\ : Span4Mux_h
    port map (
            O => \N__4050\,
            I => \N__4035\
        );

    \I__682\ : Span4Mux_v
    port map (
            O => \N__4047\,
            I => \N__4026\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__4044\,
            I => \N__4026\
        );

    \I__680\ : Span4Mux_h
    port map (
            O => \N__4041\,
            I => \N__4026\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__4038\,
            I => \N__4026\
        );

    \I__678\ : Odrv4
    port map (
            O => \N__4035\,
            I => \U400_SDRAM_SDRAM_CMD11\
        );

    \I__677\ : Odrv4
    port map (
            O => \N__4026\,
            I => \U400_SDRAM_SDRAM_CMD11\
        );

    \I__676\ : CascadeMux
    port map (
            O => \N__4021\,
            I => \U400_ADDRESS_DECODE.m20_amZ0_cascade_\
        );

    \I__675\ : CascadeMux
    port map (
            O => \N__4018\,
            I => \N__4011\
        );

    \I__674\ : InMux
    port map (
            O => \N__4017\,
            I => \N__3992\
        );

    \I__673\ : InMux
    port map (
            O => \N__4016\,
            I => \N__3992\
        );

    \I__672\ : InMux
    port map (
            O => \N__4015\,
            I => \N__3992\
        );

    \I__671\ : InMux
    port map (
            O => \N__4014\,
            I => \N__3983\
        );

    \I__670\ : InMux
    port map (
            O => \N__4011\,
            I => \N__3983\
        );

    \I__669\ : InMux
    port map (
            O => \N__4010\,
            I => \N__3983\
        );

    \I__668\ : InMux
    port map (
            O => \N__4009\,
            I => \N__3978\
        );

    \I__667\ : InMux
    port map (
            O => \N__4008\,
            I => \N__3978\
        );

    \I__666\ : InMux
    port map (
            O => \N__4007\,
            I => \N__3972\
        );

    \I__665\ : InMux
    port map (
            O => \N__4006\,
            I => \N__3972\
        );

    \I__664\ : InMux
    port map (
            O => \N__4005\,
            I => \N__3963\
        );

    \I__663\ : InMux
    port map (
            O => \N__4004\,
            I => \N__3963\
        );

    \I__662\ : InMux
    port map (
            O => \N__4003\,
            I => \N__3963\
        );

    \I__661\ : InMux
    port map (
            O => \N__4002\,
            I => \N__3956\
        );

    \I__660\ : InMux
    port map (
            O => \N__4001\,
            I => \N__3956\
        );

    \I__659\ : InMux
    port map (
            O => \N__4000\,
            I => \N__3956\
        );

    \I__658\ : InMux
    port map (
            O => \N__3999\,
            I => \N__3953\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3992\,
            I => \N__3950\
        );

    \I__656\ : InMux
    port map (
            O => \N__3991\,
            I => \N__3947\
        );

    \I__655\ : InMux
    port map (
            O => \N__3990\,
            I => \N__3944\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__3983\,
            I => \N__3941\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3978\,
            I => \N__3938\
        );

    \I__652\ : InMux
    port map (
            O => \N__3977\,
            I => \N__3935\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__3972\,
            I => \N__3931\
        );

    \I__650\ : InMux
    port map (
            O => \N__3971\,
            I => \N__3926\
        );

    \I__649\ : InMux
    port map (
            O => \N__3970\,
            I => \N__3926\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__3963\,
            I => \N__3921\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__3956\,
            I => \N__3921\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3953\,
            I => \N__3916\
        );

    \I__645\ : Span4Mux_v
    port map (
            O => \N__3950\,
            I => \N__3916\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3947\,
            I => \N__3913\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__3944\,
            I => \N__3904\
        );

    \I__642\ : Span4Mux_h
    port map (
            O => \N__3941\,
            I => \N__3904\
        );

    \I__641\ : Span4Mux_h
    port map (
            O => \N__3938\,
            I => \N__3904\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__3935\,
            I => \N__3904\
        );

    \I__639\ : InMux
    port map (
            O => \N__3934\,
            I => \N__3901\
        );

    \I__638\ : Span4Mux_h
    port map (
            O => \N__3931\,
            I => \N__3898\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__3926\,
            I => \N__3893\
        );

    \I__636\ : Span4Mux_h
    port map (
            O => \N__3921\,
            I => \N__3893\
        );

    \I__635\ : Odrv4
    port map (
            O => \N__3916\,
            I => \U400_SDRAM_SDRAM_COUNTER_3\
        );

    \I__634\ : Odrv12
    port map (
            O => \N__3913\,
            I => \U400_SDRAM_SDRAM_COUNTER_3\
        );

    \I__633\ : Odrv4
    port map (
            O => \N__3904\,
            I => \U400_SDRAM_SDRAM_COUNTER_3\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__3901\,
            I => \U400_SDRAM_SDRAM_COUNTER_3\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__3898\,
            I => \U400_SDRAM_SDRAM_COUNTER_3\
        );

    \I__630\ : Odrv4
    port map (
            O => \N__3893\,
            I => \U400_SDRAM_SDRAM_COUNTER_3\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__3880\,
            I => \N__3876\
        );

    \I__628\ : InMux
    port map (
            O => \N__3879\,
            I => \N__3872\
        );

    \I__627\ : InMux
    port map (
            O => \N__3876\,
            I => \N__3867\
        );

    \I__626\ : InMux
    port map (
            O => \N__3875\,
            I => \N__3867\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3872\,
            I => \U400_ADDRESS_DECODE.N_6_0\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3867\,
            I => \U400_ADDRESS_DECODE.N_6_0\
        );

    \I__623\ : InMux
    port map (
            O => \N__3862\,
            I => \N__3859\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__3859\,
            I => \U400_ADDRESS_DECODE.m94_bmZ0\
        );

    \I__621\ : CascadeMux
    port map (
            O => \N__3856\,
            I => \N__3852\
        );

    \I__620\ : InMux
    port map (
            O => \N__3855\,
            I => \N__3843\
        );

    \I__619\ : InMux
    port map (
            O => \N__3852\,
            I => \N__3840\
        );

    \I__618\ : InMux
    port map (
            O => \N__3851\,
            I => \N__3837\
        );

    \I__617\ : CascadeMux
    port map (
            O => \N__3850\,
            I => \N__3834\
        );

    \I__616\ : InMux
    port map (
            O => \N__3849\,
            I => \N__3831\
        );

    \I__615\ : CascadeMux
    port map (
            O => \N__3848\,
            I => \N__3827\
        );

    \I__614\ : InMux
    port map (
            O => \N__3847\,
            I => \N__3819\
        );

    \I__613\ : InMux
    port map (
            O => \N__3846\,
            I => \N__3816\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__3843\,
            I => \N__3810\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__3840\,
            I => \N__3805\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__3837\,
            I => \N__3805\
        );

    \I__609\ : InMux
    port map (
            O => \N__3834\,
            I => \N__3802\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__3831\,
            I => \N__3799\
        );

    \I__607\ : InMux
    port map (
            O => \N__3830\,
            I => \N__3792\
        );

    \I__606\ : InMux
    port map (
            O => \N__3827\,
            I => \N__3792\
        );

    \I__605\ : InMux
    port map (
            O => \N__3826\,
            I => \N__3792\
        );

    \I__604\ : InMux
    port map (
            O => \N__3825\,
            I => \N__3789\
        );

    \I__603\ : InMux
    port map (
            O => \N__3824\,
            I => \N__3784\
        );

    \I__602\ : InMux
    port map (
            O => \N__3823\,
            I => \N__3784\
        );

    \I__601\ : InMux
    port map (
            O => \N__3822\,
            I => \N__3781\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__3819\,
            I => \N__3776\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3816\,
            I => \N__3776\
        );

    \I__598\ : InMux
    port map (
            O => \N__3815\,
            I => \N__3769\
        );

    \I__597\ : InMux
    port map (
            O => \N__3814\,
            I => \N__3769\
        );

    \I__596\ : InMux
    port map (
            O => \N__3813\,
            I => \N__3769\
        );

    \I__595\ : Span4Mux_v
    port map (
            O => \N__3810\,
            I => \N__3764\
        );

    \I__594\ : Span4Mux_v
    port map (
            O => \N__3805\,
            I => \N__3764\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3802\,
            I => \N__3753\
        );

    \I__592\ : Span4Mux_h
    port map (
            O => \N__3799\,
            I => \N__3753\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__3792\,
            I => \N__3753\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3789\,
            I => \N__3753\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3784\,
            I => \N__3753\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3781\,
            I => \U400_SDRAM_SDRAM_COUNTER_1\
        );

    \I__587\ : Odrv12
    port map (
            O => \N__3776\,
            I => \U400_SDRAM_SDRAM_COUNTER_1\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__3769\,
            I => \U400_SDRAM_SDRAM_COUNTER_1\
        );

    \I__585\ : Odrv4
    port map (
            O => \N__3764\,
            I => \U400_SDRAM_SDRAM_COUNTER_1\
        );

    \I__584\ : Odrv4
    port map (
            O => \N__3753\,
            I => \U400_SDRAM_SDRAM_COUNTER_1\
        );

    \I__583\ : InMux
    port map (
            O => \N__3742\,
            I => \N__3739\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__3739\,
            I => \U400_ADDRESS_DECODE.m20_bmZ0\
        );

    \I__581\ : InMux
    port map (
            O => \N__3736\,
            I => \N__3733\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3733\,
            I => \N__3730\
        );

    \I__579\ : Span4Mux_v
    port map (
            O => \N__3730\,
            I => \N__3727\
        );

    \I__578\ : Span4Mux_h
    port map (
            O => \N__3727\,
            I => \N__3723\
        );

    \I__577\ : InMux
    port map (
            O => \N__3726\,
            I => \N__3720\
        );

    \I__576\ : Odrv4
    port map (
            O => \N__3723\,
            I => \U400_ADDRESS_DECODE.N_20_0\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__3720\,
            I => \U400_ADDRESS_DECODE.N_20_0\
        );

    \I__574\ : InMux
    port map (
            O => \N__3715\,
            I => \N__3711\
        );

    \I__573\ : InMux
    port map (
            O => \N__3714\,
            I => \N__3708\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3711\,
            I => \U400_ADDRESS_DECODE.N_179_mux\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3708\,
            I => \U400_ADDRESS_DECODE.N_179_mux\
        );

    \I__570\ : CascadeMux
    port map (
            O => \N__3703\,
            I => \U400_ADDRESS_DECODE.N_8_0_cascade_\
        );

    \I__569\ : SRMux
    port map (
            O => \N__3700\,
            I => \N__3696\
        );

    \I__568\ : SRMux
    port map (
            O => \N__3699\,
            I => \N__3692\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__3696\,
            I => \N__3689\
        );

    \I__566\ : SRMux
    port map (
            O => \N__3695\,
            I => \N__3686\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__3692\,
            I => \N__3683\
        );

    \I__564\ : Span4Mux_s3_v
    port map (
            O => \N__3689\,
            I => \N__3678\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__3686\,
            I => \N__3678\
        );

    \I__562\ : Span4Mux_s2_h
    port map (
            O => \N__3683\,
            I => \N__3673\
        );

    \I__561\ : Span4Mux_s2_h
    port map (
            O => \N__3678\,
            I => \N__3673\
        );

    \I__560\ : Odrv4
    port map (
            O => \N__3673\,
            I => \U400_SDRAM.SDRAM_CONFIGURED_RNIJKCAZ0Z2\
        );

    \I__559\ : CascadeMux
    port map (
            O => \N__3670\,
            I => \N__3667\
        );

    \I__558\ : InMux
    port map (
            O => \N__3667\,
            I => \N__3661\
        );

    \I__557\ : InMux
    port map (
            O => \N__3666\,
            I => \N__3661\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__3661\,
            I => \N__3658\
        );

    \I__555\ : Span4Mux_v
    port map (
            O => \N__3658\,
            I => \N__3655\
        );

    \I__554\ : Span4Mux_h
    port map (
            O => \N__3655\,
            I => \N__3652\
        );

    \I__553\ : Odrv4
    port map (
            O => \N__3652\,
            I => \TSn_c\
        );

    \I__552\ : InMux
    port map (
            O => \N__3649\,
            I => \N__3646\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3646\,
            I => \U400_ADDRESS_DECODE.m165_nsZ0Z_1\
        );

    \I__550\ : CascadeMux
    port map (
            O => \N__3643\,
            I => \N_13_0_cascade_\
        );

    \I__549\ : InMux
    port map (
            O => \N__3640\,
            I => \N__3632\
        );

    \I__548\ : InMux
    port map (
            O => \N__3639\,
            I => \N__3627\
        );

    \I__547\ : InMux
    port map (
            O => \N__3638\,
            I => \N__3627\
        );

    \I__546\ : InMux
    port map (
            O => \N__3637\,
            I => \N__3623\
        );

    \I__545\ : InMux
    port map (
            O => \N__3636\,
            I => \N__3620\
        );

    \I__544\ : InMux
    port map (
            O => \N__3635\,
            I => \N__3617\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__3632\,
            I => \N__3612\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__3627\,
            I => \N__3612\
        );

    \I__541\ : InMux
    port map (
            O => \N__3626\,
            I => \N__3609\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__3623\,
            I => \U400_ADDRESS_DECODE.N_10_0\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3620\,
            I => \U400_ADDRESS_DECODE.N_10_0\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3617\,
            I => \U400_ADDRESS_DECODE.N_10_0\
        );

    \I__537\ : Odrv4
    port map (
            O => \N__3612\,
            I => \U400_ADDRESS_DECODE.N_10_0\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3609\,
            I => \U400_ADDRESS_DECODE.N_10_0\
        );

    \I__535\ : InMux
    port map (
            O => \N__3598\,
            I => \N__3593\
        );

    \I__534\ : InMux
    port map (
            O => \N__3597\,
            I => \N__3590\
        );

    \I__533\ : InMux
    port map (
            O => \N__3596\,
            I => \N__3587\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3593\,
            I => \N__3584\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__3590\,
            I => \N__3581\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__3587\,
            I => \N__3577\
        );

    \I__529\ : Span4Mux_v
    port map (
            O => \N__3584\,
            I => \N__3572\
        );

    \I__528\ : Span4Mux_h
    port map (
            O => \N__3581\,
            I => \N__3572\
        );

    \I__527\ : InMux
    port map (
            O => \N__3580\,
            I => \N__3569\
        );

    \I__526\ : Odrv4
    port map (
            O => \N__3577\,
            I => \U400_ADDRESS_DECODE.N_8_0\
        );

    \I__525\ : Odrv4
    port map (
            O => \N__3572\,
            I => \U400_ADDRESS_DECODE.N_8_0\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__3569\,
            I => \U400_ADDRESS_DECODE.N_8_0\
        );

    \I__523\ : CascadeMux
    port map (
            O => \N__3562\,
            I => \U400_ADDRESS_DECODE.N_179_mux_cascade_\
        );

    \I__522\ : InMux
    port map (
            O => \N__3559\,
            I => \N__3554\
        );

    \I__521\ : InMux
    port map (
            O => \N__3558\,
            I => \N__3551\
        );

    \I__520\ : InMux
    port map (
            O => \N__3557\,
            I => \N__3548\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3554\,
            I => \U400_ADDRESS_DECODE.N_47_0\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__3551\,
            I => \U400_ADDRESS_DECODE.N_47_0\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3548\,
            I => \U400_ADDRESS_DECODE.N_47_0\
        );

    \I__516\ : InMux
    port map (
            O => \N__3541\,
            I => \N__3538\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__3538\,
            I => \U400_ADDRESS_DECODE.N_62_0\
        );

    \I__514\ : CascadeMux
    port map (
            O => \N__3535\,
            I => \U400_ADDRESS_DECODE.N_62_0_cascade_\
        );

    \I__513\ : CascadeMux
    port map (
            O => \N__3532\,
            I => \U400_ADDRESS_DECODE.m141_bmZ0_cascade_\
        );

    \I__512\ : InMux
    port map (
            O => \N__3529\,
            I => \N__3526\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3526\,
            I => \U400_ADDRESS_DECODE.m141_amZ0\
        );

    \I__510\ : CascadeMux
    port map (
            O => \N__3523\,
            I => \N__3519\
        );

    \I__509\ : CascadeMux
    port map (
            O => \N__3522\,
            I => \N__3516\
        );

    \I__508\ : InMux
    port map (
            O => \N__3519\,
            I => \N__3513\
        );

    \I__507\ : InMux
    port map (
            O => \N__3516\,
            I => \N__3510\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__3513\,
            I => \U400_SDRAM.CS0_ENZ0\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__3510\,
            I => \U400_SDRAM.CS0_ENZ0\
        );

    \I__504\ : IoInMux
    port map (
            O => \N__3505\,
            I => \N__3502\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__3502\,
            I => \N__3499\
        );

    \I__502\ : IoSpan4Mux
    port map (
            O => \N__3499\,
            I => \N__3496\
        );

    \I__501\ : Span4Mux_s2_h
    port map (
            O => \N__3496\,
            I => \N__3493\
        );

    \I__500\ : Odrv4
    port map (
            O => \N__3493\,
            I => \CS0n_c\
        );

    \I__499\ : CascadeMux
    port map (
            O => \N__3490\,
            I => \N__3487\
        );

    \I__498\ : InMux
    port map (
            O => \N__3487\,
            I => \N__3484\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3484\,
            I => \N__3481\
        );

    \I__496\ : Span4Mux_v
    port map (
            O => \N__3481\,
            I => \N__3478\
        );

    \I__495\ : Sp12to4
    port map (
            O => \N__3478\,
            I => \N__3475\
        );

    \I__494\ : Span12Mux_s9_h
    port map (
            O => \N__3475\,
            I => \N__3472\
        );

    \I__493\ : Odrv12
    port map (
            O => \N__3472\,
            I => \A_c_26\
        );

    \I__492\ : IoInMux
    port map (
            O => \N__3469\,
            I => \N__3466\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__3466\,
            I => \N__3463\
        );

    \I__490\ : Odrv4
    port map (
            O => \N__3463\,
            I => \MA_c_12\
        );

    \I__489\ : CascadeMux
    port map (
            O => \N__3460\,
            I => \N__3457\
        );

    \I__488\ : InMux
    port map (
            O => \N__3457\,
            I => \N__3454\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__3454\,
            I => \N__3451\
        );

    \I__486\ : Sp12to4
    port map (
            O => \N__3451\,
            I => \N__3448\
        );

    \I__485\ : Span12Mux_s10_v
    port map (
            O => \N__3448\,
            I => \N__3445\
        );

    \I__484\ : Odrv12
    port map (
            O => \N__3445\,
            I => \A_c_19\
        );

    \I__483\ : IoInMux
    port map (
            O => \N__3442\,
            I => \N__3439\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__3439\,
            I => \N__3436\
        );

    \I__481\ : Odrv4
    port map (
            O => \N__3436\,
            I => \MA_c_9\
        );

    \I__480\ : CascadeMux
    port map (
            O => \N__3433\,
            I => \N__3429\
        );

    \I__479\ : InMux
    port map (
            O => \N__3432\,
            I => \N__3426\
        );

    \I__478\ : InMux
    port map (
            O => \N__3429\,
            I => \N__3423\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__3426\,
            I => \N__3420\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__3423\,
            I => \U400_SDRAM_RAM_CYCLE\
        );

    \I__475\ : Odrv12
    port map (
            O => \N__3420\,
            I => \U400_SDRAM_RAM_CYCLE\
        );

    \I__474\ : InMux
    port map (
            O => \N__3415\,
            I => \N__3412\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__3412\,
            I => \U400_SDRAM_RAM_CYCLE_START_2_0\
        );

    \I__472\ : InMux
    port map (
            O => \N__3409\,
            I => \N__3406\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__3406\,
            I => \U400_ADDRESS_DECODE.N_33_0\
        );

    \I__470\ : InMux
    port map (
            O => \N__3403\,
            I => \N__3400\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3400\,
            I => \U400_ADDRESS_DECODE.m43_amZ0\
        );

    \I__468\ : InMux
    port map (
            O => \N__3397\,
            I => \N__3394\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__3394\,
            I => \U400_ADDRESS_DECODE.m87_nsZ0Z_1\
        );

    \I__466\ : CascadeMux
    port map (
            O => \N__3391\,
            I => \U400_ADDRESS_DECODE.N_88_0_cascade_\
        );

    \I__465\ : CascadeMux
    port map (
            O => \N__3388\,
            I => \N_96_0_cascade_\
        );

    \I__464\ : InMux
    port map (
            O => \N__3385\,
            I => \N__3381\
        );

    \I__463\ : InMux
    port map (
            O => \N__3384\,
            I => \N__3378\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__3381\,
            I => \N_73_0\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__3378\,
            I => \N_73_0\
        );

    \I__460\ : InMux
    port map (
            O => \N__3373\,
            I => \N__3370\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__3370\,
            I => \U400_ADDRESS_DECODE.m63_nsZ0Z_1\
        );

    \I__458\ : CascadeMux
    port map (
            O => \N__3367\,
            I => \U400_ADDRESS_DECODE.N_139_0_cascade_\
        );

    \I__457\ : CascadeMux
    port map (
            O => \N__3364\,
            I => \N__3360\
        );

    \I__456\ : CascadeMux
    port map (
            O => \N__3363\,
            I => \N__3357\
        );

    \I__455\ : InMux
    port map (
            O => \N__3360\,
            I => \N__3354\
        );

    \I__454\ : InMux
    port map (
            O => \N__3357\,
            I => \N__3351\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3354\,
            I => \N__3348\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__3351\,
            I => \U400_ADDRESS_DECODE.m133Z0Z_0\
        );

    \I__451\ : Odrv12
    port map (
            O => \N__3348\,
            I => \U400_ADDRESS_DECODE.m133Z0Z_0\
        );

    \I__450\ : CascadeMux
    port map (
            O => \N__3343\,
            I => \U400_ADDRESS_DECODE.m41_amZ0_cascade_\
        );

    \I__449\ : InMux
    port map (
            O => \N__3340\,
            I => \N__3337\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__3337\,
            I => \U400_ADDRESS_DECODE.m41_bmZ0\
        );

    \I__447\ : CascadeMux
    port map (
            O => \N__3334\,
            I => \U400_ADDRESS_DECODE.m54Z0Z_0_cascade_\
        );

    \I__446\ : InMux
    port map (
            O => \N__3331\,
            I => \N__3328\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__3328\,
            I => \U400_ADDRESS_DECODE.m56_bmZ0\
        );

    \I__444\ : InMux
    port map (
            O => \N__3325\,
            I => \N__3320\
        );

    \I__443\ : InMux
    port map (
            O => \N__3324\,
            I => \N__3317\
        );

    \I__442\ : InMux
    port map (
            O => \N__3323\,
            I => \N__3314\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__3320\,
            I => \U400_ADDRESS_DECODE.N_185\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__3317\,
            I => \U400_ADDRESS_DECODE.N_185\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__3314\,
            I => \U400_ADDRESS_DECODE.N_185\
        );

    \I__438\ : CascadeMux
    port map (
            O => \N__3307\,
            I => \U400_ADDRESS_DECODE.N_185_mux_cascade_\
        );

    \I__437\ : InMux
    port map (
            O => \N__3304\,
            I => \N__3301\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__3301\,
            I => \N__3298\
        );

    \I__435\ : Odrv4
    port map (
            O => \N__3298\,
            I => \U400_ADDRESS_DECODE.N_42_0\
        );

    \I__434\ : CascadeMux
    port map (
            O => \N__3295\,
            I => \U400_ADDRESS_DECODE.m43_bmZ0_cascade_\
        );

    \I__433\ : InMux
    port map (
            O => \N__3292\,
            I => \N__3289\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__3289\,
            I => \N_44_0\
        );

    \I__431\ : InMux
    port map (
            O => \N__3286\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_5\
        );

    \I__430\ : InMux
    port map (
            O => \N__3283\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_6\
        );

    \I__429\ : InMux
    port map (
            O => \N__3280\,
            I => \N__3276\
        );

    \I__428\ : InMux
    port map (
            O => \N__3279\,
            I => \N__3273\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__3276\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__3273\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__425\ : InMux
    port map (
            O => \N__3268\,
            I => \N__3264\
        );

    \I__424\ : InMux
    port map (
            O => \N__3267\,
            I => \N__3261\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__3264\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__3261\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__421\ : CascadeMux
    port map (
            O => \N__3256\,
            I => \N__3252\
        );

    \I__420\ : InMux
    port map (
            O => \N__3255\,
            I => \N__3249\
        );

    \I__419\ : InMux
    port map (
            O => \N__3252\,
            I => \N__3246\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__3249\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3246\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__416\ : InMux
    port map (
            O => \N__3241\,
            I => \N__3237\
        );

    \I__415\ : InMux
    port map (
            O => \N__3240\,
            I => \N__3234\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__3237\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__3234\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__412\ : CascadeMux
    port map (
            O => \N__3229\,
            I => \N_60_cascade_\
        );

    \I__411\ : CascadeMux
    port map (
            O => \N__3226\,
            I => \U400_ADDRESS_DECODE.N_98_0_cascade_\
        );

    \I__410\ : InMux
    port map (
            O => \N__3223\,
            I => \N__3216\
        );

    \I__409\ : InMux
    port map (
            O => \N__3222\,
            I => \N__3216\
        );

    \I__408\ : InMux
    port map (
            O => \N__3221\,
            I => \N__3213\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__3216\,
            I => \U400_SDRAM_SDRAM_CMD_5_sqmuxa\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__3213\,
            I => \U400_SDRAM_SDRAM_CMD_5_sqmuxa\
        );

    \I__405\ : CascadeMux
    port map (
            O => \N__3208\,
            I => \N__3205\
        );

    \I__404\ : InMux
    port map (
            O => \N__3205\,
            I => \N__3202\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__3202\,
            I => \N__3199\
        );

    \I__402\ : Span12Mux_s10_v
    port map (
            O => \N__3199\,
            I => \N__3196\
        );

    \I__401\ : Odrv12
    port map (
            O => \N__3196\,
            I => \A_c_18\
        );

    \I__400\ : InMux
    port map (
            O => \N__3193\,
            I => \N__3190\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__3190\,
            I => \N__3187\
        );

    \I__398\ : Span4Mux_h
    port map (
            O => \N__3187\,
            I => \N__3184\
        );

    \I__397\ : Sp12to4
    port map (
            O => \N__3184\,
            I => \N__3181\
        );

    \I__396\ : Span12Mux_v
    port map (
            O => \N__3181\,
            I => \N__3178\
        );

    \I__395\ : Odrv12
    port map (
            O => \N__3178\,
            I => \A_c_24\
        );

    \I__394\ : IoInMux
    port map (
            O => \N__3175\,
            I => \N__3172\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__3172\,
            I => \N__3169\
        );

    \I__392\ : Span4Mux_s1_v
    port map (
            O => \N__3169\,
            I => \N__3166\
        );

    \I__391\ : Odrv4
    port map (
            O => \N__3166\,
            I => \MA_c_8\
        );

    \I__390\ : InMux
    port map (
            O => \N__3163\,
            I => \N__3160\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__3160\,
            I => \N__3157\
        );

    \I__388\ : Odrv12
    port map (
            O => \N__3157\,
            I => \A_c_8\
        );

    \I__387\ : CascadeMux
    port map (
            O => \N__3154\,
            I => \N__3151\
        );

    \I__386\ : InMux
    port map (
            O => \N__3151\,
            I => \N__3148\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__3148\,
            I => \N__3145\
        );

    \I__384\ : Span4Mux_v
    port map (
            O => \N__3145\,
            I => \N__3142\
        );

    \I__383\ : Span4Mux_v
    port map (
            O => \N__3142\,
            I => \N__3139\
        );

    \I__382\ : Odrv4
    port map (
            O => \N__3139\,
            I => \A_c_16\
        );

    \I__381\ : IoInMux
    port map (
            O => \N__3136\,
            I => \N__3133\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__3133\,
            I => \N__3130\
        );

    \I__379\ : Odrv12
    port map (
            O => \N__3130\,
            I => \MA_c_6\
        );

    \I__378\ : InMux
    port map (
            O => \N__3127\,
            I => \N__3124\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__3124\,
            I => \U400_SDRAM.SDRAM_COUNTER_s_1\
        );

    \I__376\ : InMux
    port map (
            O => \N__3121\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_0\
        );

    \I__375\ : InMux
    port map (
            O => \N__3118\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_1\
        );

    \I__374\ : InMux
    port map (
            O => \N__3115\,
            I => \N__3112\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__3112\,
            I => \U400_SDRAM.SDRAM_COUNTER_s_3\
        );

    \I__372\ : InMux
    port map (
            O => \N__3109\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_2\
        );

    \I__371\ : InMux
    port map (
            O => \N__3106\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_3\
        );

    \I__370\ : InMux
    port map (
            O => \N__3103\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_4\
        );

    \I__369\ : CascadeMux
    port map (
            O => \N__3100\,
            I => \U400_ADDRESS_DECODE.m71_amZ0_cascade_\
        );

    \I__368\ : InMux
    port map (
            O => \N__3097\,
            I => \N__3094\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__3094\,
            I => \U400_ADDRESS_DECODE.m71_bmZ0\
        );

    \I__366\ : CascadeMux
    port map (
            O => \N__3091\,
            I => \U400_ADDRESS_DECODE.N_72_0_cascade_\
        );

    \I__365\ : CascadeMux
    port map (
            O => \N__3088\,
            I => \N_73_0_cascade_\
        );

    \I__364\ : InMux
    port map (
            O => \N__3085\,
            I => \N__3082\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__3082\,
            I => \U400_ADDRESS_DECODE.m56_amZ0\
        );

    \I__362\ : InMux
    port map (
            O => \N__3079\,
            I => \N__3076\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__3076\,
            I => \N_57_0\
        );

    \I__360\ : CascadeMux
    port map (
            O => \N__3073\,
            I => \U400_ADDRESS_DECODE.N_7_0_cascade_\
        );

    \I__359\ : IoInMux
    port map (
            O => \N__3070\,
            I => \N__3067\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__3067\,
            I => \N__3064\
        );

    \I__357\ : Odrv12
    port map (
            O => \N__3064\,
            I => \RESETn_c_i\
        );

    \I__356\ : InMux
    port map (
            O => \N__3061\,
            I => \N__3058\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__3058\,
            I => \N__3055\
        );

    \I__354\ : Odrv12
    port map (
            O => \N__3055\,
            I => \A_c_9\
        );

    \I__353\ : CascadeMux
    port map (
            O => \N__3052\,
            I => \N__3049\
        );

    \I__352\ : InMux
    port map (
            O => \N__3049\,
            I => \N__3046\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__3046\,
            I => \N__3043\
        );

    \I__350\ : Span4Mux_v
    port map (
            O => \N__3043\,
            I => \N__3040\
        );

    \I__349\ : Odrv4
    port map (
            O => \N__3040\,
            I => \A_c_17\
        );

    \I__348\ : IoInMux
    port map (
            O => \N__3037\,
            I => \N__3034\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__3034\,
            I => \N__3031\
        );

    \I__346\ : Span4Mux_s1_v
    port map (
            O => \N__3031\,
            I => \N__3028\
        );

    \I__345\ : Odrv4
    port map (
            O => \N__3028\,
            I => \MA_c_7\
        );

    \I__344\ : CascadeMux
    port map (
            O => \N__3025\,
            I => \U400_ADDRESS_DECODE.m84_amZ0_cascade_\
        );

    \I__343\ : InMux
    port map (
            O => \N__3022\,
            I => \N__3019\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__3019\,
            I => \U400_ADDRESS_DECODE.m84_bmZ0\
        );

    \I__341\ : InMux
    port map (
            O => \N__3016\,
            I => \N__3013\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__3013\,
            I => \N_85_0\
        );

    \I__339\ : InMux
    port map (
            O => \N__3010\,
            I => \N__3007\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__3007\,
            I => \U400_ADDRESS_DECODE.N_46_0\
        );

    \I__337\ : CascadeMux
    port map (
            O => \N__3004\,
            I => \U400_ADDRESS_DECODE.N_47_0_cascade_\
        );

    \I__336\ : InMux
    port map (
            O => \N__3001\,
            I => \N__2998\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__2998\,
            I => \U400_ADDRESS_DECODE.m71_amZ0Z_1\
        );

    \I__334\ : IoInMux
    port map (
            O => \N__2995\,
            I => \N__2992\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2992\,
            I => \N__2989\
        );

    \I__332\ : Odrv12
    port map (
            O => \N__2989\,
            I => \WEn_c\
        );

    \I__331\ : IoInMux
    port map (
            O => \N__2986\,
            I => \N__2983\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__2983\,
            I => \N__2980\
        );

    \I__329\ : Odrv12
    port map (
            O => \N__2980\,
            I => \RASn_c\
        );

    \I__328\ : InMux
    port map (
            O => \N__2977\,
            I => \N__2974\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__2974\,
            I => \N__2971\
        );

    \I__326\ : Span4Mux_h
    port map (
            O => \N__2971\,
            I => \N__2968\
        );

    \I__325\ : Odrv4
    port map (
            O => \N__2968\,
            I => \A_c_30\
        );

    \I__324\ : InMux
    port map (
            O => \N__2965\,
            I => \N__2962\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__2962\,
            I => \N__2959\
        );

    \I__322\ : Span4Mux_h
    port map (
            O => \N__2959\,
            I => \N__2956\
        );

    \I__321\ : Odrv4
    port map (
            O => \N__2956\,
            I => \A_c_29\
        );

    \I__320\ : CascadeMux
    port map (
            O => \N__2953\,
            I => \N__2950\
        );

    \I__319\ : InMux
    port map (
            O => \N__2950\,
            I => \N__2947\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__2947\,
            I => \A_c_28\
        );

    \I__317\ : InMux
    port map (
            O => \N__2944\,
            I => \N__2941\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__2941\,
            I => \N__2938\
        );

    \I__315\ : Odrv4
    port map (
            O => \N__2938\,
            I => \U400_ADDRESS_DECODE.m2Z0Z_1\
        );

    \I__314\ : CascadeMux
    port map (
            O => \N__2935\,
            I => \U400_ADDRESS_DECODE.N_185_cascade_\
        );

    \I__313\ : InMux
    port map (
            O => \N__2932\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_2\
        );

    \I__312\ : InMux
    port map (
            O => \N__2929\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_3\
        );

    \I__311\ : InMux
    port map (
            O => \N__2926\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_4\
        );

    \I__310\ : InMux
    port map (
            O => \N__2923\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_5\
        );

    \I__309\ : InMux
    port map (
            O => \N__2920\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_6\
        );

    \I__308\ : InMux
    port map (
            O => \N__2917\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_7\
        );

    \I__307\ : InMux
    port map (
            O => \N__2914\,
            I => \N__2910\
        );

    \I__306\ : InMux
    port map (
            O => \N__2913\,
            I => \N__2907\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__2910\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__2907\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__303\ : InMux
    port map (
            O => \N__2902\,
            I => \N__2898\
        );

    \I__302\ : InMux
    port map (
            O => \N__2901\,
            I => \N__2895\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2898\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__2895\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__299\ : InMux
    port map (
            O => \N__2890\,
            I => \N__2886\
        );

    \I__298\ : InMux
    port map (
            O => \N__2889\,
            I => \N__2883\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__2886\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__2883\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__295\ : InMux
    port map (
            O => \N__2878\,
            I => \N__2874\
        );

    \I__294\ : InMux
    port map (
            O => \N__2877\,
            I => \N__2871\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__2874\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_8\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2871\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_8\
        );

    \I__291\ : InMux
    port map (
            O => \N__2866\,
            I => \N__2862\
        );

    \I__290\ : InMux
    port map (
            O => \N__2865\,
            I => \N__2859\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2862\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2859\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__287\ : CascadeMux
    port map (
            O => \N__2854\,
            I => \U400_SDRAM.un1_REFRESH_COUNTERlt7_0_cascade_\
        );

    \I__286\ : InMux
    port map (
            O => \N__2851\,
            I => \N__2847\
        );

    \I__285\ : InMux
    port map (
            O => \N__2850\,
            I => \N__2844\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__2847\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__2844\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__282\ : IoInMux
    port map (
            O => \N__2839\,
            I => \N__2836\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2836\,
            I => \N__2833\
        );

    \I__280\ : Odrv12
    port map (
            O => \N__2833\,
            I => \CASn_c\
        );

    \I__279\ : InMux
    port map (
            O => \N__2830\,
            I => \N__2827\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2827\,
            I => \A_c_31\
        );

    \I__277\ : InMux
    port map (
            O => \N__2824\,
            I => \N__2821\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__2821\,
            I => \N__2818\
        );

    \I__275\ : Span4Mux_s1_v
    port map (
            O => \N__2818\,
            I => \N__2815\
        );

    \I__274\ : Odrv4
    port map (
            O => \N__2815\,
            I => \A_c_27\
        );

    \I__273\ : InMux
    port map (
            O => \N__2812\,
            I => \N__2808\
        );

    \I__272\ : InMux
    port map (
            O => \N__2811\,
            I => \N__2805\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__2808\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2805\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__269\ : CascadeMux
    port map (
            O => \N__2800\,
            I => \N__2795\
        );

    \I__268\ : InMux
    port map (
            O => \N__2799\,
            I => \N__2792\
        );

    \I__267\ : InMux
    port map (
            O => \N__2798\,
            I => \N__2789\
        );

    \I__266\ : InMux
    port map (
            O => \N__2795\,
            I => \N__2786\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__2792\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__2789\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__2786\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__262\ : InMux
    port map (
            O => \N__2779\,
            I => \N__2776\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__2776\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__260\ : InMux
    port map (
            O => \N__2773\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_1\
        );

    \I__259\ : IoInMux
    port map (
            O => \N__2770\,
            I => \N__2767\
        );

    \I__258\ : LocalMux
    port map (
            O => \N__2767\,
            I => \N__2764\
        );

    \I__257\ : IoSpan4Mux
    port map (
            O => \N__2764\,
            I => \N__2761\
        );

    \I__256\ : Span4Mux_s3_h
    port map (
            O => \N__2761\,
            I => \N__2758\
        );

    \I__255\ : Span4Mux_h
    port map (
            O => \N__2758\,
            I => \N__2755\
        );

    \I__254\ : Span4Mux_h
    port map (
            O => \N__2755\,
            I => \N__2752\
        );

    \I__253\ : Span4Mux_v
    port map (
            O => \N__2752\,
            I => \N__2749\
        );

    \I__252\ : Odrv4
    port map (
            O => \N__2749\,
            I => \CLK40_ibuf_gb_io_gb_input\
        );

    \INVU400_SDRAM.MA_nesr_2C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_2C_net\,
            I => \N__5248\
        );

    \INVU400_SDRAM.MA_nesr_1C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_1C_net\,
            I => \N__5247\
        );

    \INVU400_SDRAM.SDRAM_CONFIGUREDC\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_CONFIGUREDC_net\,
            I => \N__5241\
        );

    \INVU400_SDRAM.MA_nesr_10C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_10C_net\,
            I => \N__5244\
        );

    \INVU400_SDRAM.SDRAM_COUNTER_0C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_COUNTER_0C_net\,
            I => \N__5237\
        );

    \INVU400_SDRAM.BANK1C\ : INV
    port map (
            O => \INVU400_SDRAM.BANK1C_net\,
            I => \N__5240\
        );

    \INVU400_SDRAM.CS1_ENC\ : INV
    port map (
            O => \INVU400_SDRAM.CS1_ENC_net\,
            I => \N__5224\
        );

    \INVU400_SDRAM.WRITE_CYCLEC\ : INV
    port map (
            O => \INVU400_SDRAM.WRITE_CYCLEC_net\,
            I => \N__5233\
        );

    \INVU400_SDRAM.MA_nesr_12C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_12C_net\,
            I => \N__5239\
        );

    \INVU400_SDRAM.CS0_ENC\ : INV
    port map (
            O => \INVU400_SDRAM.CS0_ENC_net\,
            I => \N__5227\
        );

    \INVU400_SDRAM.SDRAM_CMD_1C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_CMD_1C_net\,
            I => \N__5232\
        );

    \INVU400_SDRAM.SDRAM_COUNTER_2C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            I => \N__5242\
        );

    \INVU400_SDRAM.MA_nesr_6C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_6C_net\,
            I => \N__5234\
        );

    \INVU400_SDRAM.MA_nesr_7C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_7C_net\,
            I => \N__5229\
        );

    \INVU400_SDRAM.SDRAM_CMD_0C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_CMD_0C_net\,
            I => \N__5226\
        );

    \INVU400_SDRAM.SDRAM_CMD_2C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_CMD_2C_net\,
            I => \N__5230\
        );

    \INVU400_SDRAM.RAM_CYCLEC\ : INV
    port map (
            O => \INVU400_SDRAM.RAM_CYCLEC_net\,
            I => \N__5235\
        );

    \INVU400_SDRAM.SDRAM_COUNTER_1C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_COUNTER_1C_net\,
            I => \N__5238\
        );

    \INVU400_SDRAM.RASnC\ : INV
    port map (
            O => \INVU400_SDRAM.RASnC_net\,
            I => \N__5223\
        );

    \INVU400_SDRAM.CASnC\ : INV
    port map (
            O => \INVU400_SDRAM.CASnC_net\,
            I => \N__5222\
        );

    \INVU400_SDRAM.REFRESH_COUNTER_2C\ : INV
    port map (
            O => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            I => \N__5228\
        );

    \INVU400_SDRAM.REFRESH_COUNTER_1C\ : INV
    port map (
            O => \INVU400_SDRAM.REFRESH_COUNTER_1C_net\,
            I => \N__5231\
        );

    \INVU400_SDRAM.REFRESH_COUNTER_0C\ : INV
    port map (
            O => \INVU400_SDRAM.REFRESH_COUNTER_0C_net\,
            I => \N__5225\
        );

    \IN_MUX_bfv_2_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_4_0_\
        );

    \IN_MUX_bfv_5_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_3_0_\
        );

    \CLK40_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2770\,
            GLOBALBUFFEROUTPUT => \CLK40_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3070\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_0_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2798\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__3699\
        );

    \U400_ADDRESS_DECODE.m2_1_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2830\,
            in2 => \_gnd_net_\,
            in3 => \N__2824\,
            lcout => \U400_ADDRESS_DECODE.m2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_1_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2799\,
            in2 => \_gnd_net_\,
            in3 => \N__2812\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__3700\
        );

    \U400_SDRAM.un3_REFRESH_COUNTER_cry_1_c_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2811\,
            in2 => \N__2800\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_4_0_\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_2_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2779\,
            in2 => \_gnd_net_\,
            in3 => \N__2773\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un3_REFRESH_COUNTER_cry_1\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_2\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3695\
        );

    \U400_SDRAM.REFRESH_COUNTER_3_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2890\,
            in2 => \_gnd_net_\,
            in3 => \N__2932\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un3_REFRESH_COUNTER_cry_2\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_3\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3695\
        );

    \U400_SDRAM.REFRESH_COUNTER_4_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2902\,
            in2 => \_gnd_net_\,
            in3 => \N__2929\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un3_REFRESH_COUNTER_cry_3\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_4\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3695\
        );

    \U400_SDRAM.REFRESH_COUNTER_5_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2914\,
            in2 => \_gnd_net_\,
            in3 => \N__2926\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un3_REFRESH_COUNTER_cry_4\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_5\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3695\
        );

    \U400_SDRAM.REFRESH_COUNTER_6_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2851\,
            in2 => \_gnd_net_\,
            in3 => \N__2923\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un3_REFRESH_COUNTER_cry_5\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_6\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3695\
        );

    \U400_SDRAM.REFRESH_COUNTER_7_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2866\,
            in2 => \_gnd_net_\,
            in3 => \N__2920\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un3_REFRESH_COUNTER_cry_6\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_7\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3695\
        );

    \U400_SDRAM.REFRESH_COUNTER_8_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2878\,
            in2 => \_gnd_net_\,
            in3 => \N__2917\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3695\
        );

    \U400_SDRAM.REFRESH_COUNTER_RNILA301_3_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__2913\,
            in1 => \N__2901\,
            in2 => \_gnd_net_\,
            in3 => \N__2889\,
            lcout => OPEN,
            ltout => \U400_SDRAM.un1_REFRESH_COUNTERlt7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_RNIJU602_8_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__2877\,
            in1 => \N__2865\,
            in2 => \N__2854\,
            in3 => \N__2850\,
            lcout => \U400_SDRAM_SDRAM_CMD11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.CASn_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6388\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CASnC_net\,
            ce => 'H',
            sr => \N__6730\
        );

    \U400_SDRAM.WEn_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6289\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CASnC_net\,
            ce => 'H',
            sr => \N__6730\
        );

    \U400_SDRAM.RASn_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5995\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.RASnC_net\,
            ce => 'H',
            sr => \N__6731\
        );

    \U400_ADDRESS_DECODE.m2_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__2977\,
            in1 => \N__2965\,
            in2 => \N__2953\,
            in3 => \N__2944\,
            lcout => \U400_ADDRESS_DECODE.N_170_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_1_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__3127\,
            in1 => \N__4723\,
            in2 => \N__5418\,
            in3 => \N__3222\,
            lcout => \U400_SDRAM_SDRAM_COUNTER_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_1C_net\,
            ce => \N__4502\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_3_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__3115\,
            in1 => \N__4724\,
            in2 => \N__5419\,
            in3 => \N__3223\,
            lcout => \U400_SDRAM_SDRAM_COUNTER_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_1C_net\,
            ce => \N__4502\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__5809\,
            in1 => \N__3221\,
            in2 => \N__3433\,
            in3 => \N__3016\,
            lcout => \U400_SDRAM_RAM_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.RAM_CYCLEC_net\,
            ce => 'H',
            sr => \N__6736\
        );

    \U400_ADDRESS_DECODE.SDRAM_COUNTERe_0_i_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__5806\,
            in1 => \N__3596\,
            in2 => \N__3363\,
            in3 => \N__3325\,
            lcout => \U400_SDRAM_SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m36_e_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4055\,
            in2 => \_gnd_net_\,
            in3 => \N__4144\,
            lcout => \U400_ADDRESS_DECODE.N_185\,
            ltout => \U400_ADDRESS_DECODE.N_185_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m71_am_1_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010111011111"
        )
    port map (
            in0 => \N__5000\,
            in1 => \N__3826\,
            in2 => \N__2935\,
            in3 => \N__3970\,
            lcout => \U400_ADDRESS_DECODE.m71_amZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m45_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011011"
        )
    port map (
            in0 => \N__3971\,
            in1 => \N__5001\,
            in2 => \N__3848\,
            in3 => \N__4818\,
            lcout => \U400_ADDRESS_DECODE.N_46_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m19_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__4819\,
            in1 => \N__5003\,
            in2 => \N__4366\,
            in3 => \N__3830\,
            lcout => \U400_ADDRESS_DECODE.N_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m84_bm_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3558\,
            in1 => \N__3990\,
            in2 => \_gnd_net_\,
            in3 => \N__3637\,
            lcout => \U400_ADDRESS_DECODE.m84_bmZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m84_am_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__4145\,
            in1 => \N__3597\,
            in2 => \_gnd_net_\,
            in3 => \N__4061\,
            lcout => OPEN,
            ltout => \U400_ADDRESS_DECODE.m84_amZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m84_ns_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__4655\,
            in1 => \_gnd_net_\,
            in2 => \N__3025\,
            in3 => \N__3022\,
            lcout => \N_85_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m71_bm_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010101"
        )
    port map (
            in0 => \N__4833\,
            in1 => \N__3847\,
            in2 => \N__5010\,
            in3 => \N__3977\,
            lcout => \U400_ADDRESS_DECODE.m71_bmZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m46_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3875\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4989\,
            lcout => \U400_ADDRESS_DECODE.N_47_0\,
            ltout => \U400_ADDRESS_DECODE.N_47_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m56_am_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010101010"
        )
    port map (
            in0 => \N__3010\,
            in1 => \_gnd_net_\,
            in2 => \N__3004\,
            in3 => \N__4652\,
            lcout => \U400_ADDRESS_DECODE.m56_amZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m71_am_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001010101"
        )
    port map (
            in0 => \N__4857\,
            in1 => \N__3324\,
            in2 => \N__3880\,
            in3 => \N__3001\,
            lcout => OPEN,
            ltout => \U400_ADDRESS_DECODE.m71_amZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m71_ns_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4653\,
            in2 => \N__3100\,
            in3 => \N__3097\,
            lcout => OPEN,
            ltout => \U400_ADDRESS_DECODE.N_72_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m72_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5807\,
            in2 => \N__3091\,
            in3 => \N__5856\,
            lcout => \N_73_0\,
            ltout => \N_73_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_2_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110111111101"
        )
    port map (
            in0 => \N__6555\,
            in1 => \N__5941\,
            in2 => \N__3088\,
            in3 => \N__3079\,
            lcout => \U400_SDRAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_CMD_2C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m56_ns_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3085\,
            in1 => \N__3331\,
            in2 => \_gnd_net_\,
            in3 => \N__5808\,
            lcout => \N_57_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m6_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4853\,
            in1 => \N__5002\,
            in2 => \_gnd_net_\,
            in3 => \N__3846\,
            lcout => OPEN,
            ltout => \U400_ADDRESS_DECODE.N_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m63_ns_1_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100101001100"
        )
    port map (
            in0 => \N__4348\,
            in1 => \N__3991\,
            in2 => \N__3073\,
            in3 => \N__3640\,
            lcout => \U400_ADDRESS_DECODE.m63_nsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_0_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111110101111"
        )
    port map (
            in0 => \N__6256\,
            in1 => \N__3292\,
            in2 => \N__6598\,
            in3 => \N__3385\,
            lcout => \U400_SDRAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_CMD_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6611\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_7_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__3061\,
            in1 => \N__5978\,
            in2 => \N__3052\,
            in3 => \N__6858\,
            lcout => \MA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_7C_net\,
            ce => \N__6802\,
            sr => \N__6735\
        );

    \U400_SDRAM.MA_nesr_8_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__6859\,
            in1 => \N__5994\,
            in2 => \N__3208\,
            in3 => \N__3193\,
            lcout => \MA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_7C_net\,
            ce => \N__6802\,
            sr => \N__6735\
        );

    \U400_SDRAM.MA_nesr_6_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__3163\,
            in1 => \N__6006\,
            in2 => \N__3154\,
            in3 => \N__6852\,
            lcout => \MA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_6C_net\,
            ce => \N__6801\,
            sr => \N__6739\
        );

    \U400_ADDRESS_DECODE.m133_0_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__6639\,
            in1 => \N__4646\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U400_ADDRESS_DECODE.m133Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_5_3_0_\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3822\,
            in2 => \_gnd_net_\,
            in3 => \N__3121\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_s_1\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_0\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_2_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4719\,
            in1 => \N__4983\,
            in2 => \_gnd_net_\,
            in3 => \N__3118\,
            lcout => \U400_SDRAM_SDRAM_COUNTER_2\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_1\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_2\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__4503\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3999\,
            in2 => \_gnd_net_\,
            in3 => \N__3109\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_s_3\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_2\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_4_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4720\,
            in1 => \N__3241\,
            in2 => \_gnd_net_\,
            in3 => \N__3106\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_3\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_4\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__4503\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_5_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4731\,
            in1 => \N__3268\,
            in2 => \_gnd_net_\,
            in3 => \N__3103\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_4\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_5\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__4503\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_6_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4721\,
            in1 => \N__3280\,
            in2 => \_gnd_net_\,
            in3 => \N__3286\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_5\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_6\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__4503\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_7_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__3255\,
            in1 => \N__4722\,
            in2 => \_gnd_net_\,
            in3 => \N__3283\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__4503\,
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m41_bm_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111101"
        )
    port map (
            in0 => \N__4923\,
            in1 => \N__3814\,
            in2 => \N__4364\,
            in3 => \N__4800\,
            lcout => \U400_ADDRESS_DECODE.m41_bmZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3279\,
            in1 => \N__3267\,
            in2 => \N__3256\,
            in3 => \N__3240\,
            lcout => \N_60\,
            ltout => \N_60_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m9_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4922\,
            in2 => \N__3229\,
            in3 => \N__3813\,
            lcout => \U400_ADDRESS_DECODE.N_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m97_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__3726\,
            in1 => \N__4117\,
            in2 => \_gnd_net_\,
            in3 => \N__4657\,
            lcout => OPEN,
            ltout => \U400_ADDRESS_DECODE.N_98_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.N_100_0_i_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110111011"
        )
    port map (
            in0 => \N__4266\,
            in1 => \N__6635\,
            in2 => \N__3226\,
            in3 => \N__5782\,
            lcout => \N_100_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m78_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__4658\,
            in1 => \N__5802\,
            in2 => \N__6640\,
            in3 => \N__3714\,
            lcout => \U400_SDRAM_SDRAM_CMD_5_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m41_am_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000111010"
        )
    port map (
            in0 => \N__5801\,
            in1 => \N__3815\,
            in2 => \N__4363\,
            in3 => \N__4801\,
            lcout => OPEN,
            ltout => \U400_ADDRESS_DECODE.m41_amZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m41_ns_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3934\,
            in2 => \N__3343\,
            in3 => \N__3340\,
            lcout => \U400_ADDRESS_DECODE.N_42_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m14_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4796\,
            in1 => \N__4948\,
            in2 => \_gnd_net_\,
            in3 => \N__4003\,
            lcout => \U400_ADDRESS_DECODE.N_15_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m5_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3823\,
            in2 => \_gnd_net_\,
            in3 => \N__4795\,
            lcout => \U400_ADDRESS_DECODE.N_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m87_ns_1_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100011011"
        )
    port map (
            in0 => \N__4004\,
            in1 => \N__3635\,
            in2 => \N__3850\,
            in3 => \N__4797\,
            lcout => \U400_ADDRESS_DECODE.m87_nsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m54_0_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__3824\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4949\,
            lcout => OPEN,
            ltout => \U400_ADDRESS_DECODE.m54Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m56_bm_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000110010001"
        )
    port map (
            in0 => \N__4005\,
            in1 => \N__4654\,
            in2 => \N__3334\,
            in3 => \N__4362\,
            lcout => \U400_ADDRESS_DECODE.m56_bmZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__6606\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3415\,
            lcout => \U400_SDRAM_RAM_CYCLE_START\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5236\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m36_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001101"
        )
    port map (
            in0 => \N__4010\,
            in1 => \N__3409\,
            in2 => \N__5011\,
            in3 => \N__3323\,
            lcout => OPEN,
            ltout => \U400_ADDRESS_DECODE.N_185_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m43_bm_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__4648\,
            in1 => \_gnd_net_\,
            in2 => \N__3307\,
            in3 => \N__3304\,
            lcout => OPEN,
            ltout => \U400_ADDRESS_DECODE.m43_bmZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m43_ns_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5783\,
            in2 => \N__3295\,
            in3 => \N__3403\,
            lcout => \N_44_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m32_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000010111011"
        )
    port map (
            in0 => \N__3825\,
            in1 => \N__4355\,
            in2 => \N__4988\,
            in3 => \N__4831\,
            lcout => \U400_ADDRESS_DECODE.N_33_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m43_am_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4832\,
            in1 => \N__4647\,
            in2 => \N__4018\,
            in3 => \N__4953\,
            lcout => \U400_ADDRESS_DECODE.m43_amZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m87_ns_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011011110110"
        )
    port map (
            in0 => \N__3397\,
            in1 => \N__4014\,
            in2 => \N__4660\,
            in3 => \N__3559\,
            lcout => OPEN,
            ltout => \U400_ADDRESS_DECODE.N_88_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m95_ns_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__4156\,
            in1 => \_gnd_net_\,
            in2 => \N__3391\,
            in3 => \N__5784\,
            lcout => OPEN,
            ltout => \N_96_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_1_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111011101"
        )
    port map (
            in0 => \N__6612\,
            in1 => \N__6357\,
            in2 => \N__3388\,
            in3 => \N__3384\,
            lcout => \U400_SDRAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_CMD_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m63_ns_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011000000110"
        )
    port map (
            in0 => \N__3373\,
            in1 => \N__4017\,
            in2 => \N__4659\,
            in3 => \N__3541\,
            lcout => \N_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m138_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__4985\,
            in1 => \N__3638\,
            in2 => \N__4347\,
            in3 => \N__4854\,
            lcout => OPEN,
            ltout => \U400_ADDRESS_DECODE.N_139_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m141_am_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__4855\,
            in1 => \N__4986\,
            in2 => \N__3367\,
            in3 => \N__4015\,
            lcout => \U400_ADDRESS_DECODE.m141_amZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m133_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000001000000"
        )
    port map (
            in0 => \N__5800\,
            in1 => \N__3598\,
            in2 => \N__3364\,
            in3 => \N__4075\,
            lcout => \N_190_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m61_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3639\,
            in1 => \N__4325\,
            in2 => \_gnd_net_\,
            in3 => \N__3557\,
            lcout => \U400_ADDRESS_DECODE.N_62_0\,
            ltout => \U400_ADDRESS_DECODE.N_62_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m141_bm_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__4016\,
            in1 => \N__5014\,
            in2 => \N__3535\,
            in3 => \N__4856\,
            lcout => OPEN,
            ltout => \U400_ADDRESS_DECODE.m141_bmZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m141_ns_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__4644\,
            in1 => \_gnd_net_\,
            in2 => \N__3532\,
            in3 => \N__3529\,
            lcout => \N_142_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.CS0_EN_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011101110"
        )
    port map (
            in0 => \N__4218\,
            in1 => \N__4228\,
            in2 => \N__3523\,
            in3 => \N__4200\,
            lcout => \U400_SDRAM.CS0_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS0_ENC_net\,
            ce => 'H',
            sr => \N__6732\
        );

    \U400_SDRAM.CS0n_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__5965\,
            in1 => \N__6367\,
            in2 => \N__3522\,
            in3 => \N__6249\,
            lcout => \CS0n_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS0_ENC_net\,
            ce => 'H',
            sr => \N__6732\
        );

    \U400_SDRAM.MA_nesr_12_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6023\,
            in1 => \N__6407\,
            in2 => \N__3490\,
            in3 => \N__6306\,
            lcout => \MA_c_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_12C_net\,
            ce => \N__6790\,
            sr => \N__6740\
        );

    \U400_SDRAM.MA_nesr_9_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6024\,
            in1 => \N__6408\,
            in2 => \N__3460\,
            in3 => \N__6307\,
            lcout => \MA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_12C_net\,
            ce => \N__6790\,
            sr => \N__6740\
        );

    \U400_ADDRESS_DECODE.m165_ns_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110100010"
        )
    port map (
            in0 => \N__3432\,
            in1 => \N__5496\,
            in2 => \N__3670\,
            in3 => \N__3649\,
            lcout => \U400_SDRAM_RAM_CYCLE_START_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m7_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3855\,
            in1 => \N__4820\,
            in2 => \N__4984\,
            in3 => \N__4006\,
            lcout => \U400_ADDRESS_DECODE.N_8_0\,
            ltout => \U400_ADDRESS_DECODE.N_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m11_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__4007\,
            in1 => \N__4607\,
            in2 => \N__3703\,
            in3 => \N__3636\,
            lcout => \U400_ADDRESS_DECODE.N_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNIJKCA2_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100110011"
        )
    port map (
            in0 => \N__4608\,
            in1 => \N__6626\,
            in2 => \N__5805\,
            in3 => \N__4100\,
            lcout => \U400_SDRAM.SDRAM_CONFIGURED_RNIJKCAZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m165_ns_1_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011111"
        )
    port map (
            in0 => \N__6625\,
            in1 => \N__3666\,
            in2 => \N__6687\,
            in3 => \N__4150\,
            lcout => \U400_ADDRESS_DECODE.m165_nsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m12_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__3851\,
            in1 => \N__4000\,
            in2 => \N__4987\,
            in3 => \N__4798\,
            lcout => \N_13_0\,
            ltout => \N_13_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m134_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__4799\,
            in1 => \N__4602\,
            in2 => \N__3643\,
            in3 => \N__4947\,
            lcout => \U400_ADDRESS_DECODE.N_135_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m64_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4601\,
            in1 => \N__4002\,
            in2 => \_gnd_net_\,
            in3 => \N__3626\,
            lcout => \N_65_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m75_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__4147\,
            in1 => \_gnd_net_\,
            in2 => \N__4078\,
            in3 => \N__3580\,
            lcout => \U400_ADDRESS_DECODE.N_179_mux\,
            ltout => \U400_ADDRESS_DECODE.N_179_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m77_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4603\,
            in2 => \N__3562\,
            in3 => \N__5803\,
            lcout => \U400_SDRAM_SDRAM_CMD_1_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m94_am_1_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001010"
        )
    port map (
            in0 => \N__4001\,
            in1 => \N__4071\,
            in2 => \N__3856\,
            in3 => \N__4146\,
            lcout => \U400_ADDRESS_DECODE.m94_amZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m94_am_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000100110010"
        )
    port map (
            in0 => \N__4009\,
            in1 => \N__4848\,
            in2 => \N__5012\,
            in3 => \N__4165\,
            lcout => OPEN,
            ltout => \U400_ADDRESS_DECODE.m94_amZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m94_ns_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__4631\,
            in1 => \_gnd_net_\,
            in2 => \N__4159\,
            in3 => \N__3862\,
            lcout => \U400_ADDRESS_DECODE.N_95_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m145_ns_1_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100001111"
        )
    port map (
            in0 => \N__4115\,
            in1 => \N__4076\,
            in2 => \N__4101\,
            in3 => \N__4148\,
            lcout => \U400_ADDRESS_DECODE.m145_nsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m20_am_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__4149\,
            in1 => \N__4116\,
            in2 => \N__4102\,
            in3 => \N__4077\,
            lcout => OPEN,
            ltout => \U400_ADDRESS_DECODE.m20_amZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m20_ns_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4630\,
            in2 => \N__4021\,
            in3 => \N__3742\,
            lcout => \U400_ADDRESS_DECODE.N_21_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m94_bm_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__4849\,
            in1 => \N__4008\,
            in2 => \_gnd_net_\,
            in3 => \N__3879\,
            lcout => \U400_ADDRESS_DECODE.m94_bmZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m20_bm_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__4996\,
            in1 => \N__3849\,
            in2 => \N__4365\,
            in3 => \N__4847\,
            lcout => \U400_ADDRESS_DECODE.m20_bmZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m153_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__5804\,
            in1 => \N__3736\,
            in2 => \N__4656\,
            in3 => \N__3715\,
            lcout => \U400_SDRAM_un1_SDRAM_COUNTER59_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.WRITE_CYCLE_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__4378\,
            in1 => \N__4329\,
            in2 => \_gnd_net_\,
            in3 => \N__5029\,
            lcout => \U400_SDRAM_WRITE_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.WRITE_CYCLEC_net\,
            ce => 'H',
            sr => \N__6733\
        );

    \U400_SDRAM.TACK_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__4398\,
            in1 => \N__4282\,
            in2 => \N__5788\,
            in3 => \N__4276\,
            lcout => \U400_SDRAM_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.WRITE_CYCLEC_net\,
            ce => 'H',
            sr => \N__6733\
        );

    \U400_ADDRESS_DECODE.m22_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000010110000"
        )
    port map (
            in0 => \N__5787\,
            in1 => \N__4270\,
            in2 => \N__6610\,
            in3 => \N__4255\,
            lcout => \N_23_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m137_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000111"
        )
    port map (
            in0 => \N__5786\,
            in1 => \N__4476\,
            in2 => \N__4246\,
            in3 => \N__5852\,
            lcout => \N_138_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m136_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001110000"
        )
    port map (
            in0 => \N__5785\,
            in1 => \N__4475\,
            in2 => \N__4245\,
            in3 => \N__5851\,
            lcout => \N_137_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.CS1_EN_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011101110"
        )
    port map (
            in0 => \N__4222\,
            in1 => \N__4207\,
            in2 => \N__4189\,
            in3 => \N__4201\,
            lcout => \U400_SDRAM.CS1_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS1_ENC_net\,
            ce => 'H',
            sr => \N__6734\
        );

    \U400_SDRAM.CS1n_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__6371\,
            in1 => \N__5979\,
            in2 => \N__4188\,
            in3 => \N__6288\,
            lcout => \CS1n_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS1_ENC_net\,
            ce => 'H',
            sr => \N__6734\
        );

    \U400_SDRAM.TA_COUNTER_4_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6608\,
            in2 => \_gnd_net_\,
            in3 => \N__5134\,
            lcout => \U400_SDRAM_TA_COUNTER_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5245\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_5_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6609\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4452\,
            lcout => \U400_SDRAM_TA_COUNTER_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5245\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m111_e_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4448\,
            in2 => \_gnd_net_\,
            in3 => \N__4436\,
            lcout => \N_174\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m102_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000101"
        )
    port map (
            in0 => \N__4437\,
            in1 => \_gnd_net_\,
            in2 => \N__4453\,
            in3 => \N__5893\,
            lcout => \U400_SDRAM_TA_OUT_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_1_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__4402\,
            in1 => \_gnd_net_\,
            in2 => \N__4420\,
            in3 => \N__6603\,
            lcout => \U400_SDRAM_TA_COUNTER_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5243\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_2_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6604\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4438\,
            lcout => \U400_SDRAM_TA_COUNTER_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5243\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m112_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100001111"
        )
    port map (
            in0 => \N__4401\,
            in1 => \N__5133\,
            in2 => \N__6624\,
            in3 => \N__5292\,
            lcout => OPEN,
            ltout => \U400_ADDRESS_DECODE.N_177_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_0_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110011111110"
        )
    port map (
            in0 => \N__5148\,
            in1 => \N__5161\,
            in2 => \N__4423\,
            in3 => \N__5863\,
            lcout => \U400_SDRAM_TA_COUNTER_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5243\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m26_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__4400\,
            in1 => \_gnd_net_\,
            in2 => \N__4419\,
            in3 => \_gnd_net_\,
            lcout => \U400_SDRAM_N_252_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_RNIF6C61_0_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6605\,
            in1 => \N__4412\,
            in2 => \_gnd_net_\,
            in3 => \N__4399\,
            lcout => \U400_SDRAM.N_252_0_0\,
            ltout => \U400_SDRAM.N_252_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_EN_i_RNO_0_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__5160\,
            in1 => \N__5144\,
            in2 => \N__5152\,
            in3 => \N__5887\,
            lcout => \U400_SDRAM.N_252_0_0_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_3_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__5888\,
            in1 => \_gnd_net_\,
            in2 => \N__5149\,
            in3 => \N__6602\,
            lcout => \U400_SDRAM_TA_COUNTER_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5243\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.BANK1_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__5062\,
            in1 => \N__5091\,
            in2 => \N__5122\,
            in3 => \N__4600\,
            lcout => \BANK1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.BANK1C_net\,
            ce => 'H',
            sr => \N__6737\
        );

    \U400_SDRAM.BANK0_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__5040\,
            in1 => \N__4599\,
            in2 => \N__5080\,
            in3 => \N__5061\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.BANK1C_net\,
            ce => 'H',
            sr => \N__6737\
        );

    \U400_SDRAM.BURST_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__5473\,
            in1 => \N__5892\,
            in2 => \N__5581\,
            in3 => \N__5025\,
            lcout => \U400_SDRAM_BURST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.BANK1C_net\,
            ce => 'H',
            sr => \N__6737\
        );

    \U400_ADDRESS_DECODE.m145_ns_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000101111"
        )
    port map (
            in0 => \N__5013\,
            in1 => \N__4858\,
            in2 => \N__4645\,
            in3 => \N__4738\,
            lcout => \U400_ADDRESS_DECODE.N_146_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_0_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001011011110"
        )
    port map (
            in0 => \N__4598\,
            in1 => \N__4732\,
            in2 => \N__4677\,
            in3 => \N__5380\,
            lcout => \U400_SDRAM_SDRAM_COUNTER_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_0C_net\,
            ce => \N__4507\,
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m149_e_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5564\,
            in2 => \_gnd_net_\,
            in3 => \N__5469\,
            lcout => \N_14_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m135_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__5725\,
            in1 => \N__5846\,
            in2 => \_gnd_net_\,
            in3 => \N__4477\,
            lcout => \U400_ADDRESS_DECODE.N_136_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m146_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__5847\,
            in1 => \N__5726\,
            in2 => \_gnd_net_\,
            in3 => \N__5425\,
            lcout => OPEN,
            ltout => \U400_ADDRESS_DECODE.N_147_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m149_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111010101"
        )
    port map (
            in0 => \N__6580\,
            in1 => \N__5400\,
            in2 => \N__5389\,
            in3 => \N__5386\,
            lcout => \N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_10_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001010"
        )
    port map (
            in0 => \N__6401\,
            in1 => \N__5374\,
            in2 => \N__6037\,
            in3 => \N__6297\,
            lcout => \MA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_10C_net\,
            ce => \N__6776\,
            sr => \N__6742\
        );

    \U400_SDRAM.MA_nesr_11_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6298\,
            in1 => \N__6027\,
            in2 => \N__5344\,
            in3 => \N__6402\,
            lcout => \MA_c_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_10C_net\,
            ce => \N__6776\,
            sr => \N__6742\
        );

    \U400_ADDRESS_DECODE.m3_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6685\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6607\,
            lcout => \U400_ADDRESS_DECODE.N_4_0\,
            ltout => \U400_ADDRESS_DECODE.N_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m123_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000111"
        )
    port map (
            in0 => \N__5603\,
            in1 => \N__5634\,
            in2 => \N__5320\,
            in3 => \N__5541\,
            lcout => \N_124_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_EN_i_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__6438\,
            in1 => \N__5305\,
            in2 => \_gnd_net_\,
            in3 => \N__5299\,
            lcout => \TA_EN_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5246\,
            ce => 'H',
            sr => \N__6741\
        );

    \U400_SDRAM.TA_OUT_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001110110001"
        )
    port map (
            in0 => \N__5293\,
            in1 => \N__5281\,
            in2 => \N__5265\,
            in3 => \N__5275\,
            lcout => \TA_OUT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5246\,
            ce => 'H',
            sr => \N__6741\
        );

    \U400_ADDRESS_DECODE.m113_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6581\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5886\,
            lcout => \U400_ADDRESS_DECODE.N_114_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5727\,
            in2 => \_gnd_net_\,
            in3 => \N__5857\,
            lcout => \U400_SDRAM_SDRAM_CONFIGURED\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_CONFIGUREDC_net\,
            ce => 'H',
            sr => \N__6738\
        );

    \U400_SDRAM.SDRAM_CMD_RNIMFKP_0_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011011110111"
        )
    port map (
            in0 => \N__6026\,
            in1 => \N__6390\,
            in2 => \N__6754\,
            in3 => \N__6291\,
            lcout => \U400_SDRAM.un1_MA20_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6025\,
            in1 => \N__6389\,
            in2 => \_gnd_net_\,
            in3 => \N__6290\,
            lcout => \U400_SDRAM.MA19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m128_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100001111"
        )
    port map (
            in0 => \N__5434\,
            in1 => \_gnd_net_\,
            in2 => \N__5605\,
            in3 => \N__5650\,
            lcout => \N_129_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m126_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__5648\,
            in1 => \N__5433\,
            in2 => \_gnd_net_\,
            in3 => \N__5596\,
            lcout => \N_127_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m127_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101001111"
        )
    port map (
            in0 => \N__5534\,
            in1 => \N__5649\,
            in2 => \N__5604\,
            in3 => \N__5489\,
            lcout => \N_128_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m121_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001000000"
        )
    port map (
            in0 => \N__5461\,
            in1 => \N__6556\,
            in2 => \N__6691\,
            in3 => \N__5576\,
            lcout => \U400_ADDRESS_DECODE.N_122_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.m125_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__5577\,
            in1 => \N__5542\,
            in2 => \N__5497\,
            in3 => \N__5462\,
            lcout => \U400_ADDRESS_DECODE.N_186_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_RNO_0_5_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111010"
        )
    port map (
            in0 => \N__6305\,
            in1 => \N__6418\,
            in2 => \N__6409\,
            in3 => \N__6032\,
            lcout => \U400_SDRAM.MA_5_iv_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_RNO_0_1_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101001110"
        )
    port map (
            in0 => \N__6031\,
            in1 => \N__6403\,
            in2 => \N__6322\,
            in3 => \N__6304\,
            lcout => \U400_SDRAM.MA_5_iv_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_1_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__6223\,
            in1 => \N__6214\,
            in2 => \_gnd_net_\,
            in3 => \N__6833\,
            lcout => \MA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_1C_net\,
            ce => \N__6777\,
            sr => \N__6746\
        );

    \U400_SDRAM.MA_nesr_5_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011111111"
        )
    port map (
            in0 => \N__6834\,
            in1 => \N__6199\,
            in2 => \_gnd_net_\,
            in3 => \N__6190\,
            lcout => \MA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_1C_net\,
            ce => \N__6777\,
            sr => \N__6746\
        );

    \U400_SDRAM.MA_nesr_3_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__6835\,
            in1 => \N__6166\,
            in2 => \N__6154\,
            in3 => \N__6035\,
            lcout => \MA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_1C_net\,
            ce => \N__6777\,
            sr => \N__6746\
        );

    \U400_SDRAM.MA_nesr_2_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__6121\,
            in1 => \N__6034\,
            in2 => \N__6106\,
            in3 => \N__6850\,
            lcout => \MA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_2C_net\,
            ce => \N__6800\,
            sr => \N__6747\
        );

    \U400_SDRAM.MA_nesr_4_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__6851\,
            in1 => \N__6091\,
            in2 => \N__6079\,
            in3 => \N__6036\,
            lcout => \MA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_2C_net\,
            ce => \N__6800\,
            sr => \N__6747\
        );

    \U400_SDRAM.MA_nesr_0_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__6049\,
            in1 => \N__6033\,
            in2 => \N__6874\,
            in3 => \N__6849\,
            lcout => \MA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_2C_net\,
            ce => \N__6800\,
            sr => \N__6747\
        );

    \U400_ADDRESS_DECODE.N_4_0_i_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__6686\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6519\,
            lcout => \N_4_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TAn_obuft_RNO_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6445\,
            lcout => \N_304_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 30 2025 12:31:54

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    CMA : out std_logic_vector(10 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    A : in std_logic_vector(20 downto 0);
    RAMENn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    DBRn : in std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__12169\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7827\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \N_861_i\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A20C_net\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \A_c_14\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_\ : std_logic;
signal \LATCH_CLK_c\ : std_logic;
signal \U712_CHIP_RAM.LATCH_CLK_RNOZ0Z_0\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DBENn_8_0\ : std_logic;
signal \U712_CHIP_RAM.N_341\ : std_logic;
signal \U712_CHIP_RAM.N_341_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0\ : std_logic;
signal \A_c_20\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.N_387_cascade_\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_186_cascade_\ : std_logic;
signal \U712_CHIP_RAM.BANK0_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_387\ : std_logic;
signal \U712_CHIP_RAM.N_385_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_223\ : std_logic;
signal \U712_CHIP_RAM.N_335_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_342_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_6_0_a2_2\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_6_0_a2_1\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_6_0_cascade_\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0\ : std_logic;
signal \U712_CHIP_RAM.N_385\ : std_logic;
signal \U712_CHIP_RAM.N_338_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_305_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_239_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_208\ : std_logic;
signal \U712_CYCLE_TERM.N_217_i_0_en_0\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.START_RSTZ0\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \U712_REG_SM.N_270_cascade_\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_289\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.BANK0_RNOZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z20\ : std_logic;
signal \U712_CHIP_RAM.N_305\ : std_logic;
signal \U712_CHIP_RAM.BANK0_RNOZ0Z_1_cascade_\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \U712_CHIP_RAM.BANK0_RNOZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.N_186\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_0_a2_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_306\ : std_logic;
signal \U712_CHIP_RAM.N_333_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_0_0_a2_1_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER18_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_239\ : std_logic;
signal \U712_CHIP_RAM.N_269\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_0_0_a2_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \bfn_10_12_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.N_46\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CYCLE_TERM.N_217_i_0_en\ : std_logic;
signal \U712_REG_SM.START_RST_0_sqmuxa\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_0\ : std_logic;
signal \U712_REG_SM.N_285_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER18\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_srsts_i_0_a2_0_0_0\ : std_logic;
signal \U712_REG_SM.N_222\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ1Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_284_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.N_134\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\ : std_logic;
signal \N_116_i\ : std_logic;
signal \U712_CHIP_RAM.N_207_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_333\ : std_logic;
signal \U712_CHIP_RAM.N_310_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \U712_CHIP_RAM.N_334\ : std_logic;
signal \U712_CHIP_RAM.N_297\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_202\ : std_logic;
signal \U712_CHIP_RAM.N_184_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_304\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERlde_0_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.N_392_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_0\ : std_logic;
signal \U712_REG_SM.N_196\ : std_logic;
signal \U712_REG_SM.N_383\ : std_logic;
signal \U712_REG_SM.N_383_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.N_321_cascade_\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \N_156_i\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1Z0Z_0\ : std_logic;
signal \N_126_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_315\ : std_logic;
signal \U712_BYTE_ENABLE.N_319\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_1\ : std_logic;
signal \U712_REG_SM.un1_STATE_COUNT_4_i_i_0\ : std_logic;
signal \U712_REG_SM.N_26\ : std_logic;
signal \U712_REG_SM.N_274\ : std_logic;
signal \DMA_LATCH_EN_c\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_8\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.N_207\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_262\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_237\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.N_335\ : std_logic;
signal \U712_CHIP_RAM.N_261\ : std_logic;
signal \U712_CHIP_RAM.N_180\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_386\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_338\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_1_2\ : std_logic;
signal \U712_CHIP_RAM.N_342\ : std_logic;
signal \U712_CHIP_RAM.N_293_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_294\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_1_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.N_235_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_REG_SM.N_281\ : std_logic;
signal \U712_REG_SM.N_235\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_212\ : std_logic;
signal \U712_REG_SM.REG_TACK_RNOZ0Z_0\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0Z0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_220_cascade_\ : std_logic;
signal \N_151_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_314\ : std_logic;
signal \U712_BYTE_ENABLE.UUBE\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \WEn_c\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_2\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_236_cascade_\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_273\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \A_c_19\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \UMBEn_c\ : std_logic;
signal \U712_BYTE_ENABLE_UUBE_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \U712_BYTE_ENABLE_un1_UDSn_i\ : std_logic;
signal \LLBEn_c\ : std_logic;
signal \DS_ENm\ : std_logic;
signal \N_119\ : std_logic;
signal \A_c_1\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \N_220_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \CASn_c\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_0\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \RnW_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \WRITE_CYCLEm\ : std_logic;
signal \N_238\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__4113\,
            RESETB => \N__5976\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12169\,
            DIN => \N__12168\,
            DOUT => \N__12167\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12169\,
            PADOUT => \N__12168\,
            PADIN => \N__12167\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5586\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12160\,
            DIN => \N__12159\,
            DOUT => \N__12158\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12160\,
            PADOUT => \N__12159\,
            PADIN => \N__12158\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12151\,
            DIN => \N__12150\,
            DOUT => \N__12149\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12151\,
            PADOUT => \N__12150\,
            PADIN => \N__12149\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9246\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12142\,
            DIN => \N__12141\,
            DOUT => \N__12140\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12142\,
            PADOUT => \N__12141\,
            PADIN => \N__12140\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11064\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12133\,
            DIN => \N__12132\,
            DOUT => \N__12131\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12133\,
            PADOUT => \N__12132\,
            PADIN => \N__12131\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12124\,
            DIN => \N__12123\,
            DOUT => \N__12122\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12124\,
            PADOUT => \N__12123\,
            PADIN => \N__12122\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12115\,
            DIN => \N__12114\,
            DOUT => \N__12113\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12115\,
            PADOUT => \N__12114\,
            PADIN => \N__12113\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12106\,
            DIN => \N__12105\,
            DOUT => \N__12104\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12106\,
            PADOUT => \N__12105\,
            PADIN => \N__12104\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12097\,
            DIN => \N__12096\,
            DOUT => \N__12095\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12097\,
            PADOUT => \N__12096\,
            PADIN => \N__12095\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12088\,
            DIN => \N__12087\,
            DOUT => \N__12086\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12088\,
            PADOUT => \N__12087\,
            PADIN => \N__12086\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12079\,
            DIN => \N__12078\,
            DOUT => \N__12077\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12079\,
            PADOUT => \N__12078\,
            PADIN => \N__12077\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8979\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12070\,
            DIN => \N__12069\,
            DOUT => \N__12068\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12070\,
            PADOUT => \N__12069\,
            PADIN => \N__12068\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9063\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12061\,
            DIN => \N__12060\,
            DOUT => \N__12059\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12061\,
            PADOUT => \N__12060\,
            PADIN => \N__12059\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12052\,
            DIN => \N__12051\,
            DOUT => \N__12050\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12052\,
            PADOUT => \N__12051\,
            PADIN => \N__12050\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4674\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12043\,
            DIN => \N__12042\,
            DOUT => \N__12041\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12043\,
            PADOUT => \N__12042\,
            PADIN => \N__12041\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12034\,
            DIN => \N__12033\,
            DOUT => \N__12032\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12034\,
            PADOUT => \N__12033\,
            PADIN => \N__12032\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12025\,
            DIN => \N__12024\,
            DOUT => \N__12023\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12025\,
            PADOUT => \N__12024\,
            PADIN => \N__12023\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4296\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12016\,
            DIN => \N__12015\,
            DOUT => \N__12014\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12016\,
            PADOUT => \N__12015\,
            PADIN => \N__12014\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12007\,
            DIN => \N__12006\,
            DOUT => \N__12005\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12007\,
            PADOUT => \N__12006\,
            PADIN => \N__12005\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11998\,
            DIN => \N__11997\,
            DOUT => \N__11996\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11998\,
            PADOUT => \N__11997\,
            PADIN => \N__11996\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11049\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11989\,
            DIN => \N__11988\,
            DOUT => \N__11987\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11989\,
            PADOUT => \N__11988\,
            PADIN => \N__11987\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11980\,
            DIN => \N__11979\,
            DOUT => \N__11978\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11980\,
            PADOUT => \N__11979\,
            PADIN => \N__11978\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9003\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11971\,
            DIN => \N__11970\,
            DOUT => \N__11969\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11971\,
            PADOUT => \N__11970\,
            PADIN => \N__11969\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11962\,
            DIN => \N__11961\,
            DOUT => \N__11960\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11962\,
            PADOUT => \N__11961\,
            PADIN => \N__11960\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9774\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11953\,
            DIN => \N__11952\,
            DOUT => \N__11951\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11953\,
            PADOUT => \N__11952\,
            PADIN => \N__11951\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11944\,
            DIN => \N__11943\,
            DOUT => \N__11942\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11944\,
            PADOUT => \N__11943\,
            PADIN => \N__11942\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11935\,
            DIN => \N__11934\,
            DOUT => \N__11933\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11935\,
            PADOUT => \N__11934\,
            PADIN => \N__11933\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11926\,
            DIN => \N__11925\,
            DOUT => \N__11924\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11926\,
            PADOUT => \N__11925\,
            PADIN => \N__11924\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11917\,
            DIN => \N__11916\,
            DOUT => \N__11915\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11917\,
            PADOUT => \N__11916\,
            PADIN => \N__11915\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11908\,
            DIN => \N__11907\,
            DOUT => \N__11906\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11908\,
            PADOUT => \N__11907\,
            PADIN => \N__11906\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5997\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11899\,
            DIN => \N__11898\,
            DOUT => \N__11897\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11899\,
            PADOUT => \N__11898\,
            PADIN => \N__11897\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11890\,
            DIN => \N__11889\,
            DOUT => \N__11888\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11890\,
            PADOUT => \N__11889\,
            PADIN => \N__11888\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11881\,
            DIN => \N__11880\,
            DOUT => \N__11879\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11881\,
            PADOUT => \N__11880\,
            PADIN => \N__11879\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11872\,
            DIN => \N__11871\,
            DOUT => \N__11870\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11872\,
            PADOUT => \N__11871\,
            PADIN => \N__11870\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11863\,
            DIN => \N__11862\,
            DOUT => \N__11861\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11863\,
            PADOUT => \N__11862\,
            PADIN => \N__11861\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11854\,
            DIN => \N__11853\,
            DOUT => \N__11852\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11854\,
            PADOUT => \N__11853\,
            PADIN => \N__11852\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7698\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11845\,
            DIN => \N__11844\,
            DOUT => \N__11843\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11845\,
            PADOUT => \N__11844\,
            PADIN => \N__11843\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4986\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11836\,
            DIN => \N__11835\,
            DOUT => \N__11834\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11836\,
            PADOUT => \N__11835\,
            PADIN => \N__11834\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11827\,
            DIN => \N__11826\,
            DOUT => \N__11825\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11827\,
            PADOUT => \N__11826\,
            PADIN => \N__11825\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4722\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11818\,
            DIN => \N__11817\,
            DOUT => \N__11816\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11818\,
            PADOUT => \N__11817\,
            PADIN => \N__11816\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10728\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11809\,
            DIN => \N__11808\,
            DOUT => \N__11807\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11809\,
            PADOUT => \N__11808\,
            PADIN => \N__11807\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11800\,
            DIN => \N__11799\,
            DOUT => \N__11798\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11800\,
            PADOUT => \N__11799\,
            PADIN => \N__11798\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11791\,
            DIN => \N__11790\,
            DOUT => \N__11789\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11791\,
            PADOUT => \N__11790\,
            PADIN => \N__11789\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11782\,
            DIN => \N__11781\,
            DOUT => \N__11780\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11782\,
            PADOUT => \N__11781\,
            PADIN => \N__11780\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11773\,
            DIN => \N__11772\,
            DOUT => \N__11771\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11773\,
            PADOUT => \N__11772\,
            PADIN => \N__11771\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7566\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11764\,
            DIN => \N__11763\,
            DOUT => \N__11762\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11764\,
            PADOUT => \N__11763\,
            PADIN => \N__11762\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11755\,
            DIN => \N__11754\,
            DOUT => \N__11753\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11755\,
            PADOUT => \N__11754\,
            PADIN => \N__11753\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8569\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11746\,
            DIN => \N__11745\,
            DOUT => \N__11744\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11746\,
            PADOUT => \N__11745\,
            PADIN => \N__11744\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8952\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11737\,
            DIN => \N__11736\,
            DOUT => \N__11735\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11737\,
            PADOUT => \N__11736\,
            PADIN => \N__11735\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9804\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11728\,
            DIN => \N__11727\,
            DOUT => \N__11726\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11728\,
            PADOUT => \N__11727\,
            PADIN => \N__11726\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5805\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11719\,
            DIN => \N__11718\,
            DOUT => \N__11717\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11719\,
            PADOUT => \N__11718\,
            PADIN => \N__11717\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7935\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11710\,
            DIN => \N__11709\,
            DOUT => \N__11708\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11710\,
            PADOUT => \N__11709\,
            PADIN => \N__11708\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4718\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11701\,
            DIN => \N__11700\,
            DOUT => \N__11699\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11701\,
            PADOUT => \N__11700\,
            PADIN => \N__11699\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11692\,
            DIN => \N__11691\,
            DOUT => \N__11690\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11692\,
            PADOUT => \N__11691\,
            PADIN => \N__11690\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11683\,
            DIN => \N__11682\,
            DOUT => \N__11681\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11683\,
            PADOUT => \N__11682\,
            PADIN => \N__11681\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7239\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11674\,
            DIN => \N__11673\,
            DOUT => \N__11672\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11674\,
            PADOUT => \N__11673\,
            PADIN => \N__11672\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7713\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11665\,
            DIN => \N__11664\,
            DOUT => \N__11663\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11665\,
            PADOUT => \N__11664\,
            PADIN => \N__11663\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4209\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11656\,
            DIN => \N__11655\,
            DOUT => \N__11654\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11656\,
            PADOUT => \N__11655\,
            PADIN => \N__11654\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5769\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11647\,
            DIN => \N__11646\,
            DOUT => \N__11645\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11647\,
            PADOUT => \N__11646\,
            PADIN => \N__11645\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11638\,
            DIN => \N__11637\,
            DOUT => \N__11636\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11638\,
            PADOUT => \N__11637\,
            PADIN => \N__11636\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11629\,
            DIN => \N__11628\,
            DOUT => \N__11627\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11629\,
            PADOUT => \N__11628\,
            PADIN => \N__11627\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11620\,
            DIN => \N__11619\,
            DOUT => \N__11618\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11620\,
            PADOUT => \N__11619\,
            PADIN => \N__11618\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11611\,
            DIN => \N__11610\,
            DOUT => \N__11609\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11611\,
            PADOUT => \N__11610\,
            PADIN => \N__11609\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4821\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11602\,
            DIN => \N__11601\,
            DOUT => \N__11600\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11602\,
            PADOUT => \N__11601\,
            PADIN => \N__11600\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9414\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11593\,
            DIN => \N__11592\,
            DOUT => \N__11591\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11593\,
            PADOUT => \N__11592\,
            PADIN => \N__11591\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11584\,
            DIN => \N__11583\,
            DOUT => \N__11582\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11584\,
            PADOUT => \N__11583\,
            PADIN => \N__11582\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5427\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11575\,
            DIN => \N__11574\,
            DOUT => \N__11573\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11575\,
            PADOUT => \N__11574\,
            PADIN => \N__11573\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4158\,
            DIN0 => OPEN,
            DOUT0 => \N__4488\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11566\,
            DIN => \N__11565\,
            DOUT => \N__11564\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11566\,
            PADOUT => \N__11565\,
            PADIN => \N__11564\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7794\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11557\,
            DIN => \N__11556\,
            DOUT => \N__11555\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11557\,
            PADOUT => \N__11556\,
            PADIN => \N__11555\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11548\,
            DIN => \N__11547\,
            DOUT => \N__11546\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11548\,
            PADOUT => \N__11547\,
            PADIN => \N__11546\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11539\,
            DIN => \N__11538\,
            DOUT => \N__11537\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11539\,
            PADOUT => \N__11538\,
            PADIN => \N__11537\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7524\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11530\,
            DIN => \N__11529\,
            DOUT => \N__11528\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11530\,
            PADOUT => \N__11529\,
            PADIN => \N__11528\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11521\,
            DIN => \N__11520\,
            DOUT => \N__11519\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11521\,
            PADOUT => \N__11520\,
            PADIN => \N__11519\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11512\,
            DIN => \N__11511\,
            DOUT => \N__11510\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11512\,
            PADOUT => \N__11511\,
            PADIN => \N__11510\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11503\,
            DIN => \N__11502\,
            DOUT => \N__11501\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11503\,
            PADOUT => \N__11502\,
            PADIN => \N__11501\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11494\,
            DIN => \N__11493\,
            DOUT => \N__11492\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11494\,
            PADOUT => \N__11493\,
            PADIN => \N__11492\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4449\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11485\,
            DIN => \N__11484\,
            DOUT => \N__11483\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11485\,
            PADOUT => \N__11484\,
            PADIN => \N__11483\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9792\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11476\,
            DIN => \N__11475\,
            DOUT => \N__11474\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11476\,
            PADOUT => \N__11475\,
            PADIN => \N__11474\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8517\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11467\,
            DIN => \N__11466\,
            DOUT => \N__11465\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11467\,
            PADOUT => \N__11466\,
            PADIN => \N__11465\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4608\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11458\,
            DIN => \N__11457\,
            DOUT => \N__11456\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11458\,
            PADOUT => \N__11457\,
            PADIN => \N__11456\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11449\,
            DIN => \N__11448\,
            DOUT => \N__11447\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11449\,
            PADOUT => \N__11448\,
            PADIN => \N__11447\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11440\,
            DIN => \N__11439\,
            DOUT => \N__11438\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11440\,
            PADOUT => \N__11439\,
            PADIN => \N__11438\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9087\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11431\,
            DIN => \N__11430\,
            DOUT => \N__11429\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11431\,
            PADOUT => \N__11430\,
            PADIN => \N__11429\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11422\,
            DIN => \N__11421\,
            DOUT => \N__11420\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11422\,
            PADOUT => \N__11421\,
            PADIN => \N__11420\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11413\,
            DIN => \N__11412\,
            DOUT => \N__11411\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11413\,
            PADOUT => \N__11412\,
            PADIN => \N__11411\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4242\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11404\,
            DIN => \N__11403\,
            DOUT => \N__11402\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11404\,
            PADOUT => \N__11403\,
            PADIN => \N__11402\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9732\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11395\,
            DIN => \N__11394\,
            DOUT => \N__11393\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11395\,
            PADOUT => \N__11394\,
            PADIN => \N__11393\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8571\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11386\,
            DIN => \N__11385\,
            DOUT => \N__11384\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11386\,
            PADOUT => \N__11385\,
            PADIN => \N__11384\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11377\,
            DIN => \N__11376\,
            DOUT => \N__11375\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11377\,
            PADOUT => \N__11376\,
            PADIN => \N__11375\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8570\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11368\,
            DIN => \N__11367\,
            DOUT => \N__11366\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11368\,
            PADOUT => \N__11367\,
            PADIN => \N__11366\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4173\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2773\ : InMux
    port map (
            O => \N__11349\,
            I => \N__11346\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__11346\,
            I => \N__11342\
        );

    \I__2771\ : InMux
    port map (
            O => \N__11345\,
            I => \N__11338\
        );

    \I__2770\ : Span4Mux_v
    port map (
            O => \N__11342\,
            I => \N__11335\
        );

    \I__2769\ : InMux
    port map (
            O => \N__11341\,
            I => \N__11331\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__11338\,
            I => \N__11328\
        );

    \I__2767\ : Span4Mux_v
    port map (
            O => \N__11335\,
            I => \N__11325\
        );

    \I__2766\ : InMux
    port map (
            O => \N__11334\,
            I => \N__11322\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__11331\,
            I => \N__11319\
        );

    \I__2764\ : Span12Mux_h
    port map (
            O => \N__11328\,
            I => \N__11316\
        );

    \I__2763\ : Sp12to4
    port map (
            O => \N__11325\,
            I => \N__11313\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__11322\,
            I => \N__11310\
        );

    \I__2761\ : Span12Mux_h
    port map (
            O => \N__11319\,
            I => \N__11307\
        );

    \I__2760\ : Span12Mux_h
    port map (
            O => \N__11316\,
            I => \N__11304\
        );

    \I__2759\ : Span12Mux_h
    port map (
            O => \N__11313\,
            I => \N__11299\
        );

    \I__2758\ : Span12Mux_v
    port map (
            O => \N__11310\,
            I => \N__11299\
        );

    \I__2757\ : Span12Mux_v
    port map (
            O => \N__11307\,
            I => \N__11296\
        );

    \I__2756\ : Span12Mux_v
    port map (
            O => \N__11304\,
            I => \N__11291\
        );

    \I__2755\ : Span12Mux_h
    port map (
            O => \N__11299\,
            I => \N__11291\
        );

    \I__2754\ : Odrv12
    port map (
            O => \N__11296\,
            I => \RnW_c\
        );

    \I__2753\ : Odrv12
    port map (
            O => \N__11291\,
            I => \RnW_c\
        );

    \I__2752\ : InMux
    port map (
            O => \N__11286\,
            I => \N__11283\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__11283\,
            I => \N__11280\
        );

    \I__2750\ : Span4Mux_v
    port map (
            O => \N__11280\,
            I => \N__11276\
        );

    \I__2749\ : InMux
    port map (
            O => \N__11279\,
            I => \N__11273\
        );

    \I__2748\ : Span4Mux_v
    port map (
            O => \N__11276\,
            I => \N__11267\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__11273\,
            I => \N__11267\
        );

    \I__2746\ : InMux
    port map (
            O => \N__11272\,
            I => \N__11263\
        );

    \I__2745\ : Span4Mux_h
    port map (
            O => \N__11267\,
            I => \N__11260\
        );

    \I__2744\ : InMux
    port map (
            O => \N__11266\,
            I => \N__11257\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__11263\,
            I => \N__11254\
        );

    \I__2742\ : Span4Mux_v
    port map (
            O => \N__11260\,
            I => \N__11249\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__11257\,
            I => \N__11249\
        );

    \I__2740\ : Sp12to4
    port map (
            O => \N__11254\,
            I => \N__11244\
        );

    \I__2739\ : Span4Mux_v
    port map (
            O => \N__11249\,
            I => \N__11241\
        );

    \I__2738\ : InMux
    port map (
            O => \N__11248\,
            I => \N__11236\
        );

    \I__2737\ : InMux
    port map (
            O => \N__11247\,
            I => \N__11236\
        );

    \I__2736\ : Span12Mux_v
    port map (
            O => \N__11244\,
            I => \N__11233\
        );

    \I__2735\ : Sp12to4
    port map (
            O => \N__11241\,
            I => \N__11230\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__11236\,
            I => \N__11227\
        );

    \I__2733\ : Span12Mux_h
    port map (
            O => \N__11233\,
            I => \N__11224\
        );

    \I__2732\ : Span12Mux_h
    port map (
            O => \N__11230\,
            I => \N__11221\
        );

    \I__2731\ : Span4Mux_v
    port map (
            O => \N__11227\,
            I => \N__11218\
        );

    \I__2730\ : Odrv12
    port map (
            O => \N__11224\,
            I => \CASUn_c\
        );

    \I__2729\ : Odrv12
    port map (
            O => \N__11221\,
            I => \CASUn_c\
        );

    \I__2728\ : Odrv4
    port map (
            O => \N__11218\,
            I => \CASUn_c\
        );

    \I__2727\ : CascadeMux
    port map (
            O => \N__11211\,
            I => \N__11206\
        );

    \I__2726\ : InMux
    port map (
            O => \N__11210\,
            I => \N__11202\
        );

    \I__2725\ : InMux
    port map (
            O => \N__11209\,
            I => \N__11197\
        );

    \I__2724\ : InMux
    port map (
            O => \N__11206\,
            I => \N__11197\
        );

    \I__2723\ : InMux
    port map (
            O => \N__11205\,
            I => \N__11194\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__11202\,
            I => \N__11191\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__11197\,
            I => \N__11187\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__11194\,
            I => \N__11184\
        );

    \I__2719\ : Span4Mux_v
    port map (
            O => \N__11191\,
            I => \N__11181\
        );

    \I__2718\ : CascadeMux
    port map (
            O => \N__11190\,
            I => \N__11177\
        );

    \I__2717\ : Sp12to4
    port map (
            O => \N__11187\,
            I => \N__11172\
        );

    \I__2716\ : Sp12to4
    port map (
            O => \N__11184\,
            I => \N__11172\
        );

    \I__2715\ : Sp12to4
    port map (
            O => \N__11181\,
            I => \N__11169\
        );

    \I__2714\ : InMux
    port map (
            O => \N__11180\,
            I => \N__11164\
        );

    \I__2713\ : InMux
    port map (
            O => \N__11177\,
            I => \N__11164\
        );

    \I__2712\ : Span12Mux_v
    port map (
            O => \N__11172\,
            I => \N__11161\
        );

    \I__2711\ : Span12Mux_h
    port map (
            O => \N__11169\,
            I => \N__11156\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__11164\,
            I => \N__11156\
        );

    \I__2709\ : Span12Mux_h
    port map (
            O => \N__11161\,
            I => \N__11151\
        );

    \I__2708\ : Span12Mux_v
    port map (
            O => \N__11156\,
            I => \N__11151\
        );

    \I__2707\ : Odrv12
    port map (
            O => \N__11151\,
            I => \CASLn_c\
        );

    \I__2706\ : InMux
    port map (
            O => \N__11148\,
            I => \N__11144\
        );

    \I__2705\ : InMux
    port map (
            O => \N__11147\,
            I => \N__11141\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__11144\,
            I => \N__11138\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__11141\,
            I => \N__11133\
        );

    \I__2702\ : Span4Mux_v
    port map (
            O => \N__11138\,
            I => \N__11129\
        );

    \I__2701\ : InMux
    port map (
            O => \N__11137\,
            I => \N__11124\
        );

    \I__2700\ : InMux
    port map (
            O => \N__11136\,
            I => \N__11124\
        );

    \I__2699\ : Span4Mux_h
    port map (
            O => \N__11133\,
            I => \N__11120\
        );

    \I__2698\ : InMux
    port map (
            O => \N__11132\,
            I => \N__11117\
        );

    \I__2697\ : Span4Mux_v
    port map (
            O => \N__11129\,
            I => \N__11112\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__11124\,
            I => \N__11112\
        );

    \I__2695\ : InMux
    port map (
            O => \N__11123\,
            I => \N__11109\
        );

    \I__2694\ : Sp12to4
    port map (
            O => \N__11120\,
            I => \N__11106\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__11117\,
            I => \N__11101\
        );

    \I__2692\ : Span4Mux_v
    port map (
            O => \N__11112\,
            I => \N__11101\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__11109\,
            I => \N__11097\
        );

    \I__2690\ : Span12Mux_v
    port map (
            O => \N__11106\,
            I => \N__11089\
        );

    \I__2689\ : Sp12to4
    port map (
            O => \N__11101\,
            I => \N__11089\
        );

    \I__2688\ : InMux
    port map (
            O => \N__11100\,
            I => \N__11086\
        );

    \I__2687\ : Span4Mux_v
    port map (
            O => \N__11097\,
            I => \N__11083\
        );

    \I__2686\ : InMux
    port map (
            O => \N__11096\,
            I => \N__11080\
        );

    \I__2685\ : InMux
    port map (
            O => \N__11095\,
            I => \N__11075\
        );

    \I__2684\ : InMux
    port map (
            O => \N__11094\,
            I => \N__11075\
        );

    \I__2683\ : Odrv12
    port map (
            O => \N__11089\,
            I => \WRITE_CYCLEm\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__11086\,
            I => \WRITE_CYCLEm\
        );

    \I__2681\ : Odrv4
    port map (
            O => \N__11083\,
            I => \WRITE_CYCLEm\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__11080\,
            I => \WRITE_CYCLEm\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__11075\,
            I => \WRITE_CYCLEm\
        );

    \I__2678\ : IoInMux
    port map (
            O => \N__11064\,
            I => \N__11061\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__11061\,
            I => \N__11058\
        );

    \I__2676\ : Span4Mux_s3_h
    port map (
            O => \N__11058\,
            I => \N__11055\
        );

    \I__2675\ : Span4Mux_v
    port map (
            O => \N__11055\,
            I => \N__11052\
        );

    \I__2674\ : Odrv4
    port map (
            O => \N__11052\,
            I => \N_238\
        );

    \I__2673\ : IoInMux
    port map (
            O => \N__11049\,
            I => \N__11046\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__11046\,
            I => \N__11043\
        );

    \I__2671\ : IoSpan4Mux
    port map (
            O => \N__11043\,
            I => \N__11040\
        );

    \I__2670\ : Span4Mux_s3_v
    port map (
            O => \N__11040\,
            I => \N__11037\
        );

    \I__2669\ : Sp12to4
    port map (
            O => \N__11037\,
            I => \N__11034\
        );

    \I__2668\ : Span12Mux_v
    port map (
            O => \N__11034\,
            I => \N__11031\
        );

    \I__2667\ : Odrv12
    port map (
            O => \N__11031\,
            I => \CMA_c_0\
        );

    \I__2666\ : InMux
    port map (
            O => \N__11028\,
            I => \N__11024\
        );

    \I__2665\ : InMux
    port map (
            O => \N__11027\,
            I => \N__11019\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__11024\,
            I => \N__11016\
        );

    \I__2663\ : InMux
    port map (
            O => \N__11023\,
            I => \N__11013\
        );

    \I__2662\ : InMux
    port map (
            O => \N__11022\,
            I => \N__11010\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__11019\,
            I => \N__11007\
        );

    \I__2660\ : Span4Mux_v
    port map (
            O => \N__11016\,
            I => \N__11000\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__11013\,
            I => \N__11000\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__11010\,
            I => \N__11000\
        );

    \I__2657\ : Span4Mux_h
    port map (
            O => \N__11007\,
            I => \N__10995\
        );

    \I__2656\ : Span4Mux_h
    port map (
            O => \N__11000\,
            I => \N__10995\
        );

    \I__2655\ : Sp12to4
    port map (
            O => \N__10995\,
            I => \N__10992\
        );

    \I__2654\ : Span12Mux_v
    port map (
            O => \N__10992\,
            I => \N__10989\
        );

    \I__2653\ : Odrv12
    port map (
            O => \N__10989\,
            I => \DRA_c_1\
        );

    \I__2652\ : InMux
    port map (
            O => \N__10986\,
            I => \N__10983\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__10983\,
            I => \N__10979\
        );

    \I__2650\ : InMux
    port map (
            O => \N__10982\,
            I => \N__10976\
        );

    \I__2649\ : Sp12to4
    port map (
            O => \N__10979\,
            I => \N__10971\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__10976\,
            I => \N__10971\
        );

    \I__2647\ : Span12Mux_v
    port map (
            O => \N__10971\,
            I => \N__10968\
        );

    \I__2646\ : Span12Mux_h
    port map (
            O => \N__10968\,
            I => \N__10965\
        );

    \I__2645\ : Odrv12
    port map (
            O => \N__10965\,
            I => \DRA_c_0\
        );

    \I__2644\ : InMux
    port map (
            O => \N__10962\,
            I => \N__10959\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__10959\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2642\ : InMux
    port map (
            O => \N__10956\,
            I => \N__10953\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__10953\,
            I => \N__10949\
        );

    \I__2640\ : InMux
    port map (
            O => \N__10952\,
            I => \N__10946\
        );

    \I__2639\ : Span4Mux_h
    port map (
            O => \N__10949\,
            I => \N__10943\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__10946\,
            I => \N__10940\
        );

    \I__2637\ : Span4Mux_h
    port map (
            O => \N__10943\,
            I => \N__10937\
        );

    \I__2636\ : Span12Mux_v
    port map (
            O => \N__10940\,
            I => \N__10934\
        );

    \I__2635\ : Odrv4
    port map (
            O => \N__10937\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2634\ : Odrv12
    port map (
            O => \N__10934\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2633\ : InMux
    port map (
            O => \N__10929\,
            I => \N__10926\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__10926\,
            I => \N__10920\
        );

    \I__2631\ : InMux
    port map (
            O => \N__10925\,
            I => \N__10915\
        );

    \I__2630\ : InMux
    port map (
            O => \N__10924\,
            I => \N__10915\
        );

    \I__2629\ : InMux
    port map (
            O => \N__10923\,
            I => \N__10912\
        );

    \I__2628\ : Span4Mux_h
    port map (
            O => \N__10920\,
            I => \N__10907\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__10915\,
            I => \N__10907\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__10912\,
            I => \N__10904\
        );

    \I__2625\ : Span4Mux_v
    port map (
            O => \N__10907\,
            I => \N__10901\
        );

    \I__2624\ : Span12Mux_v
    port map (
            O => \N__10904\,
            I => \N__10898\
        );

    \I__2623\ : Sp12to4
    port map (
            O => \N__10901\,
            I => \N__10895\
        );

    \I__2622\ : Span12Mux_h
    port map (
            O => \N__10898\,
            I => \N__10892\
        );

    \I__2621\ : Odrv12
    port map (
            O => \N__10895\,
            I => \DRA_c_5\
        );

    \I__2620\ : Odrv12
    port map (
            O => \N__10892\,
            I => \DRA_c_5\
        );

    \I__2619\ : InMux
    port map (
            O => \N__10887\,
            I => \N__10884\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__10884\,
            I => \N__10881\
        );

    \I__2617\ : Odrv4
    port map (
            O => \N__10881\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2616\ : InMux
    port map (
            O => \N__10878\,
            I => \N__10873\
        );

    \I__2615\ : InMux
    port map (
            O => \N__10877\,
            I => \N__10870\
        );

    \I__2614\ : InMux
    port map (
            O => \N__10876\,
            I => \N__10867\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__10873\,
            I => \N__10862\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__10870\,
            I => \N__10859\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__10867\,
            I => \N__10856\
        );

    \I__2610\ : InMux
    port map (
            O => \N__10866\,
            I => \N__10851\
        );

    \I__2609\ : InMux
    port map (
            O => \N__10865\,
            I => \N__10851\
        );

    \I__2608\ : Span4Mux_h
    port map (
            O => \N__10862\,
            I => \N__10845\
        );

    \I__2607\ : Span4Mux_h
    port map (
            O => \N__10859\,
            I => \N__10845\
        );

    \I__2606\ : Span4Mux_h
    port map (
            O => \N__10856\,
            I => \N__10842\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__10851\,
            I => \N__10839\
        );

    \I__2604\ : InMux
    port map (
            O => \N__10850\,
            I => \N__10836\
        );

    \I__2603\ : Odrv4
    port map (
            O => \N__10845\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\
        );

    \I__2602\ : Odrv4
    port map (
            O => \N__10842\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\
        );

    \I__2601\ : Odrv12
    port map (
            O => \N__10839\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__10836\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\
        );

    \I__2599\ : CascadeMux
    port map (
            O => \N__10827\,
            I => \N__10822\
        );

    \I__2598\ : CascadeMux
    port map (
            O => \N__10826\,
            I => \N__10816\
        );

    \I__2597\ : CascadeMux
    port map (
            O => \N__10825\,
            I => \N__10813\
        );

    \I__2596\ : InMux
    port map (
            O => \N__10822\,
            I => \N__10810\
        );

    \I__2595\ : CascadeMux
    port map (
            O => \N__10821\,
            I => \N__10807\
        );

    \I__2594\ : CascadeMux
    port map (
            O => \N__10820\,
            I => \N__10804\
        );

    \I__2593\ : CascadeMux
    port map (
            O => \N__10819\,
            I => \N__10799\
        );

    \I__2592\ : InMux
    port map (
            O => \N__10816\,
            I => \N__10795\
        );

    \I__2591\ : InMux
    port map (
            O => \N__10813\,
            I => \N__10792\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__10810\,
            I => \N__10789\
        );

    \I__2589\ : InMux
    port map (
            O => \N__10807\,
            I => \N__10784\
        );

    \I__2588\ : InMux
    port map (
            O => \N__10804\,
            I => \N__10784\
        );

    \I__2587\ : InMux
    port map (
            O => \N__10803\,
            I => \N__10781\
        );

    \I__2586\ : InMux
    port map (
            O => \N__10802\,
            I => \N__10778\
        );

    \I__2585\ : InMux
    port map (
            O => \N__10799\,
            I => \N__10775\
        );

    \I__2584\ : CascadeMux
    port map (
            O => \N__10798\,
            I => \N__10772\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__10795\,
            I => \N__10769\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__10792\,
            I => \N__10762\
        );

    \I__2581\ : Span4Mux_h
    port map (
            O => \N__10789\,
            I => \N__10762\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__10784\,
            I => \N__10762\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__10781\,
            I => \N__10755\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__10778\,
            I => \N__10755\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__10775\,
            I => \N__10755\
        );

    \I__2576\ : InMux
    port map (
            O => \N__10772\,
            I => \N__10752\
        );

    \I__2575\ : Span4Mux_v
    port map (
            O => \N__10769\,
            I => \N__10747\
        );

    \I__2574\ : Span4Mux_v
    port map (
            O => \N__10762\,
            I => \N__10747\
        );

    \I__2573\ : Span4Mux_h
    port map (
            O => \N__10755\,
            I => \N__10744\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__10752\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2571\ : Odrv4
    port map (
            O => \N__10747\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__10744\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2569\ : InMux
    port map (
            O => \N__10737\,
            I => \N__10734\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__10734\,
            I => \N__10731\
        );

    \I__2567\ : Odrv4
    port map (
            O => \N__10731\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__2566\ : IoInMux
    port map (
            O => \N__10728\,
            I => \N__10725\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__10725\,
            I => \N__10722\
        );

    \I__2564\ : Span4Mux_s0_h
    port map (
            O => \N__10722\,
            I => \N__10719\
        );

    \I__2563\ : Sp12to4
    port map (
            O => \N__10719\,
            I => \N__10716\
        );

    \I__2562\ : Span12Mux_s6_v
    port map (
            O => \N__10716\,
            I => \N__10713\
        );

    \I__2561\ : Span12Mux_h
    port map (
            O => \N__10713\,
            I => \N__10710\
        );

    \I__2560\ : Odrv12
    port map (
            O => \N__10710\,
            I => \CMA_c_3\
        );

    \I__2559\ : InMux
    port map (
            O => \N__10707\,
            I => \N__10704\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__10704\,
            I => \N__10663\
        );

    \I__2557\ : ClkMux
    port map (
            O => \N__10703\,
            I => \N__10569\
        );

    \I__2556\ : ClkMux
    port map (
            O => \N__10702\,
            I => \N__10569\
        );

    \I__2555\ : ClkMux
    port map (
            O => \N__10701\,
            I => \N__10569\
        );

    \I__2554\ : ClkMux
    port map (
            O => \N__10700\,
            I => \N__10569\
        );

    \I__2553\ : ClkMux
    port map (
            O => \N__10699\,
            I => \N__10569\
        );

    \I__2552\ : ClkMux
    port map (
            O => \N__10698\,
            I => \N__10569\
        );

    \I__2551\ : ClkMux
    port map (
            O => \N__10697\,
            I => \N__10569\
        );

    \I__2550\ : ClkMux
    port map (
            O => \N__10696\,
            I => \N__10569\
        );

    \I__2549\ : ClkMux
    port map (
            O => \N__10695\,
            I => \N__10569\
        );

    \I__2548\ : ClkMux
    port map (
            O => \N__10694\,
            I => \N__10569\
        );

    \I__2547\ : ClkMux
    port map (
            O => \N__10693\,
            I => \N__10569\
        );

    \I__2546\ : ClkMux
    port map (
            O => \N__10692\,
            I => \N__10569\
        );

    \I__2545\ : ClkMux
    port map (
            O => \N__10691\,
            I => \N__10569\
        );

    \I__2544\ : ClkMux
    port map (
            O => \N__10690\,
            I => \N__10569\
        );

    \I__2543\ : ClkMux
    port map (
            O => \N__10689\,
            I => \N__10569\
        );

    \I__2542\ : ClkMux
    port map (
            O => \N__10688\,
            I => \N__10569\
        );

    \I__2541\ : ClkMux
    port map (
            O => \N__10687\,
            I => \N__10569\
        );

    \I__2540\ : ClkMux
    port map (
            O => \N__10686\,
            I => \N__10569\
        );

    \I__2539\ : ClkMux
    port map (
            O => \N__10685\,
            I => \N__10569\
        );

    \I__2538\ : ClkMux
    port map (
            O => \N__10684\,
            I => \N__10569\
        );

    \I__2537\ : ClkMux
    port map (
            O => \N__10683\,
            I => \N__10569\
        );

    \I__2536\ : ClkMux
    port map (
            O => \N__10682\,
            I => \N__10569\
        );

    \I__2535\ : ClkMux
    port map (
            O => \N__10681\,
            I => \N__10569\
        );

    \I__2534\ : ClkMux
    port map (
            O => \N__10680\,
            I => \N__10569\
        );

    \I__2533\ : ClkMux
    port map (
            O => \N__10679\,
            I => \N__10569\
        );

    \I__2532\ : ClkMux
    port map (
            O => \N__10678\,
            I => \N__10569\
        );

    \I__2531\ : ClkMux
    port map (
            O => \N__10677\,
            I => \N__10569\
        );

    \I__2530\ : ClkMux
    port map (
            O => \N__10676\,
            I => \N__10569\
        );

    \I__2529\ : ClkMux
    port map (
            O => \N__10675\,
            I => \N__10569\
        );

    \I__2528\ : ClkMux
    port map (
            O => \N__10674\,
            I => \N__10569\
        );

    \I__2527\ : ClkMux
    port map (
            O => \N__10673\,
            I => \N__10569\
        );

    \I__2526\ : ClkMux
    port map (
            O => \N__10672\,
            I => \N__10569\
        );

    \I__2525\ : ClkMux
    port map (
            O => \N__10671\,
            I => \N__10569\
        );

    \I__2524\ : ClkMux
    port map (
            O => \N__10670\,
            I => \N__10569\
        );

    \I__2523\ : ClkMux
    port map (
            O => \N__10669\,
            I => \N__10569\
        );

    \I__2522\ : ClkMux
    port map (
            O => \N__10668\,
            I => \N__10569\
        );

    \I__2521\ : ClkMux
    port map (
            O => \N__10667\,
            I => \N__10569\
        );

    \I__2520\ : ClkMux
    port map (
            O => \N__10666\,
            I => \N__10569\
        );

    \I__2519\ : Glb2LocalMux
    port map (
            O => \N__10663\,
            I => \N__10569\
        );

    \I__2518\ : ClkMux
    port map (
            O => \N__10662\,
            I => \N__10569\
        );

    \I__2517\ : ClkMux
    port map (
            O => \N__10661\,
            I => \N__10569\
        );

    \I__2516\ : ClkMux
    port map (
            O => \N__10660\,
            I => \N__10569\
        );

    \I__2515\ : ClkMux
    port map (
            O => \N__10659\,
            I => \N__10569\
        );

    \I__2514\ : ClkMux
    port map (
            O => \N__10658\,
            I => \N__10569\
        );

    \I__2513\ : GlobalMux
    port map (
            O => \N__10569\,
            I => \CLK80_PLL\
        );

    \I__2512\ : CEMux
    port map (
            O => \N__10566\,
            I => \N__10562\
        );

    \I__2511\ : CEMux
    port map (
            O => \N__10565\,
            I => \N__10557\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__10562\,
            I => \N__10551\
        );

    \I__2509\ : CEMux
    port map (
            O => \N__10561\,
            I => \N__10548\
        );

    \I__2508\ : CEMux
    port map (
            O => \N__10560\,
            I => \N__10544\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__10557\,
            I => \N__10540\
        );

    \I__2506\ : CEMux
    port map (
            O => \N__10556\,
            I => \N__10537\
        );

    \I__2505\ : CEMux
    port map (
            O => \N__10555\,
            I => \N__10534\
        );

    \I__2504\ : CEMux
    port map (
            O => \N__10554\,
            I => \N__10531\
        );

    \I__2503\ : Span4Mux_v
    port map (
            O => \N__10551\,
            I => \N__10526\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__10548\,
            I => \N__10526\
        );

    \I__2501\ : CEMux
    port map (
            O => \N__10547\,
            I => \N__10523\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__10544\,
            I => \N__10520\
        );

    \I__2499\ : CEMux
    port map (
            O => \N__10543\,
            I => \N__10517\
        );

    \I__2498\ : Span4Mux_h
    port map (
            O => \N__10540\,
            I => \N__10512\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__10537\,
            I => \N__10512\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__10534\,
            I => \N__10509\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__10531\,
            I => \N__10506\
        );

    \I__2494\ : Span4Mux_v
    port map (
            O => \N__10526\,
            I => \N__10503\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__10523\,
            I => \N__10500\
        );

    \I__2492\ : Span4Mux_h
    port map (
            O => \N__10520\,
            I => \N__10495\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__10517\,
            I => \N__10495\
        );

    \I__2490\ : Span4Mux_h
    port map (
            O => \N__10512\,
            I => \N__10492\
        );

    \I__2489\ : Span4Mux_v
    port map (
            O => \N__10509\,
            I => \N__10489\
        );

    \I__2488\ : Span4Mux_h
    port map (
            O => \N__10506\,
            I => \N__10486\
        );

    \I__2487\ : Span4Mux_h
    port map (
            O => \N__10503\,
            I => \N__10483\
        );

    \I__2486\ : Span4Mux_h
    port map (
            O => \N__10500\,
            I => \N__10480\
        );

    \I__2485\ : Span4Mux_v
    port map (
            O => \N__10495\,
            I => \N__10477\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__10492\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2483\ : Odrv4
    port map (
            O => \N__10489\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2482\ : Odrv4
    port map (
            O => \N__10486\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2481\ : Odrv4
    port map (
            O => \N__10483\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__10480\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2479\ : Odrv4
    port map (
            O => \N__10477\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2478\ : InMux
    port map (
            O => \N__10464\,
            I => \N__10460\
        );

    \I__2477\ : InMux
    port map (
            O => \N__10463\,
            I => \N__10457\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__10460\,
            I => \N__10450\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__10457\,
            I => \N__10450\
        );

    \I__2474\ : InMux
    port map (
            O => \N__10456\,
            I => \N__10447\
        );

    \I__2473\ : InMux
    port map (
            O => \N__10455\,
            I => \N__10444\
        );

    \I__2472\ : Span4Mux_v
    port map (
            O => \N__10450\,
            I => \N__10441\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__10447\,
            I => \N__10436\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__10444\,
            I => \N__10436\
        );

    \I__2469\ : Sp12to4
    port map (
            O => \N__10441\,
            I => \N__10433\
        );

    \I__2468\ : Span4Mux_v
    port map (
            O => \N__10436\,
            I => \N__10430\
        );

    \I__2467\ : Span12Mux_h
    port map (
            O => \N__10433\,
            I => \N__10427\
        );

    \I__2466\ : Sp12to4
    port map (
            O => \N__10430\,
            I => \N__10424\
        );

    \I__2465\ : Odrv12
    port map (
            O => \N__10427\,
            I => \DRA_c_6\
        );

    \I__2464\ : Odrv12
    port map (
            O => \N__10424\,
            I => \DRA_c_6\
        );

    \I__2463\ : InMux
    port map (
            O => \N__10419\,
            I => \N__10414\
        );

    \I__2462\ : InMux
    port map (
            O => \N__10418\,
            I => \N__10410\
        );

    \I__2461\ : InMux
    port map (
            O => \N__10417\,
            I => \N__10407\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__10414\,
            I => \N__10404\
        );

    \I__2459\ : InMux
    port map (
            O => \N__10413\,
            I => \N__10401\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__10410\,
            I => \N__10396\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__10407\,
            I => \N__10396\
        );

    \I__2456\ : Span12Mux_v
    port map (
            O => \N__10404\,
            I => \N__10391\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__10401\,
            I => \N__10391\
        );

    \I__2454\ : Span12Mux_h
    port map (
            O => \N__10396\,
            I => \N__10388\
        );

    \I__2453\ : Span12Mux_h
    port map (
            O => \N__10391\,
            I => \N__10385\
        );

    \I__2452\ : Odrv12
    port map (
            O => \N__10388\,
            I => \DRA_c_7\
        );

    \I__2451\ : Odrv12
    port map (
            O => \N__10385\,
            I => \DRA_c_7\
        );

    \I__2450\ : InMux
    port map (
            O => \N__10380\,
            I => \N__10377\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__10377\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2448\ : InMux
    port map (
            O => \N__10374\,
            I => \N__10369\
        );

    \I__2447\ : InMux
    port map (
            O => \N__10373\,
            I => \N__10366\
        );

    \I__2446\ : InMux
    port map (
            O => \N__10372\,
            I => \N__10363\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__10369\,
            I => \N__10357\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__10366\,
            I => \N__10357\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__10363\,
            I => \N__10354\
        );

    \I__2442\ : InMux
    port map (
            O => \N__10362\,
            I => \N__10351\
        );

    \I__2441\ : Span4Mux_v
    port map (
            O => \N__10357\,
            I => \N__10348\
        );

    \I__2440\ : Span4Mux_h
    port map (
            O => \N__10354\,
            I => \N__10343\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__10351\,
            I => \N__10343\
        );

    \I__2438\ : Sp12to4
    port map (
            O => \N__10348\,
            I => \N__10340\
        );

    \I__2437\ : Span4Mux_v
    port map (
            O => \N__10343\,
            I => \N__10337\
        );

    \I__2436\ : Span12Mux_h
    port map (
            O => \N__10340\,
            I => \N__10334\
        );

    \I__2435\ : Sp12to4
    port map (
            O => \N__10337\,
            I => \N__10331\
        );

    \I__2434\ : Odrv12
    port map (
            O => \N__10334\,
            I => \DRA_c_3\
        );

    \I__2433\ : Odrv12
    port map (
            O => \N__10331\,
            I => \DRA_c_3\
        );

    \I__2432\ : InMux
    port map (
            O => \N__10326\,
            I => \N__10322\
        );

    \I__2431\ : InMux
    port map (
            O => \N__10325\,
            I => \N__10319\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__10322\,
            I => \N__10316\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__10319\,
            I => \N__10312\
        );

    \I__2428\ : Span4Mux_v
    port map (
            O => \N__10316\,
            I => \N__10304\
        );

    \I__2427\ : InMux
    port map (
            O => \N__10315\,
            I => \N__10301\
        );

    \I__2426\ : Span4Mux_v
    port map (
            O => \N__10312\,
            I => \N__10293\
        );

    \I__2425\ : InMux
    port map (
            O => \N__10311\,
            I => \N__10290\
        );

    \I__2424\ : InMux
    port map (
            O => \N__10310\,
            I => \N__10284\
        );

    \I__2423\ : InMux
    port map (
            O => \N__10309\,
            I => \N__10281\
        );

    \I__2422\ : InMux
    port map (
            O => \N__10308\,
            I => \N__10278\
        );

    \I__2421\ : InMux
    port map (
            O => \N__10307\,
            I => \N__10275\
        );

    \I__2420\ : Span4Mux_h
    port map (
            O => \N__10304\,
            I => \N__10270\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__10301\,
            I => \N__10270\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10300\,
            I => \N__10267\
        );

    \I__2417\ : InMux
    port map (
            O => \N__10299\,
            I => \N__10264\
        );

    \I__2416\ : InMux
    port map (
            O => \N__10298\,
            I => \N__10261\
        );

    \I__2415\ : InMux
    port map (
            O => \N__10297\,
            I => \N__10258\
        );

    \I__2414\ : InMux
    port map (
            O => \N__10296\,
            I => \N__10255\
        );

    \I__2413\ : Span4Mux_h
    port map (
            O => \N__10293\,
            I => \N__10247\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__10290\,
            I => \N__10244\
        );

    \I__2411\ : InMux
    port map (
            O => \N__10289\,
            I => \N__10241\
        );

    \I__2410\ : InMux
    port map (
            O => \N__10288\,
            I => \N__10236\
        );

    \I__2409\ : InMux
    port map (
            O => \N__10287\,
            I => \N__10236\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__10284\,
            I => \N__10227\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__10281\,
            I => \N__10227\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__10278\,
            I => \N__10227\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__10275\,
            I => \N__10227\
        );

    \I__2404\ : Span4Mux_v
    port map (
            O => \N__10270\,
            I => \N__10222\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__10267\,
            I => \N__10222\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__10264\,
            I => \N__10215\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__10261\,
            I => \N__10215\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__10258\,
            I => \N__10215\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__10255\,
            I => \N__10212\
        );

    \I__2398\ : InMux
    port map (
            O => \N__10254\,
            I => \N__10209\
        );

    \I__2397\ : InMux
    port map (
            O => \N__10253\,
            I => \N__10204\
        );

    \I__2396\ : InMux
    port map (
            O => \N__10252\,
            I => \N__10204\
        );

    \I__2395\ : InMux
    port map (
            O => \N__10251\,
            I => \N__10201\
        );

    \I__2394\ : InMux
    port map (
            O => \N__10250\,
            I => \N__10198\
        );

    \I__2393\ : Span4Mux_h
    port map (
            O => \N__10247\,
            I => \N__10187\
        );

    \I__2392\ : Span4Mux_v
    port map (
            O => \N__10244\,
            I => \N__10187\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__10241\,
            I => \N__10187\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__10236\,
            I => \N__10187\
        );

    \I__2389\ : Span4Mux_v
    port map (
            O => \N__10227\,
            I => \N__10187\
        );

    \I__2388\ : Span4Mux_h
    port map (
            O => \N__10222\,
            I => \N__10180\
        );

    \I__2387\ : Span4Mux_v
    port map (
            O => \N__10215\,
            I => \N__10180\
        );

    \I__2386\ : Span4Mux_v
    port map (
            O => \N__10212\,
            I => \N__10180\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__10209\,
            I => \N__10175\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__10204\,
            I => \N__10175\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__10201\,
            I => \N__10166\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__10198\,
            I => \N__10166\
        );

    \I__2381\ : Sp12to4
    port map (
            O => \N__10187\,
            I => \N__10166\
        );

    \I__2380\ : Sp12to4
    port map (
            O => \N__10180\,
            I => \N__10166\
        );

    \I__2379\ : Span12Mux_v
    port map (
            O => \N__10175\,
            I => \N__10163\
        );

    \I__2378\ : Span12Mux_h
    port map (
            O => \N__10166\,
            I => \N__10160\
        );

    \I__2377\ : Span12Mux_h
    port map (
            O => \N__10163\,
            I => \N__10157\
        );

    \I__2376\ : Span12Mux_v
    port map (
            O => \N__10160\,
            I => \N__10154\
        );

    \I__2375\ : Odrv12
    port map (
            O => \N__10157\,
            I => \AGNUS_REV_c\
        );

    \I__2374\ : Odrv12
    port map (
            O => \N__10154\,
            I => \AGNUS_REV_c\
        );

    \I__2373\ : InMux
    port map (
            O => \N__10149\,
            I => \N__10143\
        );

    \I__2372\ : InMux
    port map (
            O => \N__10148\,
            I => \N__10140\
        );

    \I__2371\ : InMux
    port map (
            O => \N__10147\,
            I => \N__10137\
        );

    \I__2370\ : InMux
    port map (
            O => \N__10146\,
            I => \N__10134\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__10143\,
            I => \N__10129\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__10140\,
            I => \N__10129\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__10137\,
            I => \N__10126\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__10134\,
            I => \N__10123\
        );

    \I__2365\ : Span4Mux_v
    port map (
            O => \N__10129\,
            I => \N__10120\
        );

    \I__2364\ : Span4Mux_v
    port map (
            O => \N__10126\,
            I => \N__10117\
        );

    \I__2363\ : Span12Mux_v
    port map (
            O => \N__10123\,
            I => \N__10110\
        );

    \I__2362\ : Sp12to4
    port map (
            O => \N__10120\,
            I => \N__10110\
        );

    \I__2361\ : Sp12to4
    port map (
            O => \N__10117\,
            I => \N__10110\
        );

    \I__2360\ : Span12Mux_h
    port map (
            O => \N__10110\,
            I => \N__10107\
        );

    \I__2359\ : Odrv12
    port map (
            O => \N__10107\,
            I => \DRA_c_4\
        );

    \I__2358\ : InMux
    port map (
            O => \N__10104\,
            I => \N__10101\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__10101\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2356\ : ClkMux
    port map (
            O => \N__10098\,
            I => \N__10074\
        );

    \I__2355\ : ClkMux
    port map (
            O => \N__10097\,
            I => \N__10074\
        );

    \I__2354\ : ClkMux
    port map (
            O => \N__10096\,
            I => \N__10074\
        );

    \I__2353\ : ClkMux
    port map (
            O => \N__10095\,
            I => \N__10074\
        );

    \I__2352\ : ClkMux
    port map (
            O => \N__10094\,
            I => \N__10074\
        );

    \I__2351\ : ClkMux
    port map (
            O => \N__10093\,
            I => \N__10074\
        );

    \I__2350\ : ClkMux
    port map (
            O => \N__10092\,
            I => \N__10074\
        );

    \I__2349\ : ClkMux
    port map (
            O => \N__10091\,
            I => \N__10074\
        );

    \I__2348\ : GlobalMux
    port map (
            O => \N__10074\,
            I => \N__10071\
        );

    \I__2347\ : gio2CtrlBuf
    port map (
            O => \N__10071\,
            I => \C3_c_g\
        );

    \I__2346\ : CEMux
    port map (
            O => \N__10068\,
            I => \N__10023\
        );

    \I__2345\ : CEMux
    port map (
            O => \N__10067\,
            I => \N__10023\
        );

    \I__2344\ : CEMux
    port map (
            O => \N__10066\,
            I => \N__10023\
        );

    \I__2343\ : CEMux
    port map (
            O => \N__10065\,
            I => \N__10023\
        );

    \I__2342\ : CEMux
    port map (
            O => \N__10064\,
            I => \N__10023\
        );

    \I__2341\ : CEMux
    port map (
            O => \N__10063\,
            I => \N__10023\
        );

    \I__2340\ : CEMux
    port map (
            O => \N__10062\,
            I => \N__10023\
        );

    \I__2339\ : CEMux
    port map (
            O => \N__10061\,
            I => \N__10023\
        );

    \I__2338\ : CEMux
    port map (
            O => \N__10060\,
            I => \N__10023\
        );

    \I__2337\ : CEMux
    port map (
            O => \N__10059\,
            I => \N__10023\
        );

    \I__2336\ : CEMux
    port map (
            O => \N__10058\,
            I => \N__10023\
        );

    \I__2335\ : CEMux
    port map (
            O => \N__10057\,
            I => \N__10023\
        );

    \I__2334\ : CEMux
    port map (
            O => \N__10056\,
            I => \N__10023\
        );

    \I__2333\ : CEMux
    port map (
            O => \N__10055\,
            I => \N__10023\
        );

    \I__2332\ : CEMux
    port map (
            O => \N__10054\,
            I => \N__10023\
        );

    \I__2331\ : GlobalMux
    port map (
            O => \N__10023\,
            I => \N__10020\
        );

    \I__2330\ : gio2CtrlBuf
    port map (
            O => \N__10020\,
            I => \DBRn_c_i_0_g\
        );

    \I__2329\ : InMux
    port map (
            O => \N__10017\,
            I => \N__10010\
        );

    \I__2328\ : InMux
    port map (
            O => \N__10016\,
            I => \N__10007\
        );

    \I__2327\ : InMux
    port map (
            O => \N__10015\,
            I => \N__10004\
        );

    \I__2326\ : InMux
    port map (
            O => \N__10014\,
            I => \N__10001\
        );

    \I__2325\ : InMux
    port map (
            O => \N__10013\,
            I => \N__9998\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__10010\,
            I => \N__9995\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__10007\,
            I => \N__9975\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__10004\,
            I => \N__9962\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__10001\,
            I => \N__9955\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__9998\,
            I => \N__9947\
        );

    \I__2319\ : Glb2LocalMux
    port map (
            O => \N__9995\,
            I => \N__9849\
        );

    \I__2318\ : SRMux
    port map (
            O => \N__9994\,
            I => \N__9849\
        );

    \I__2317\ : SRMux
    port map (
            O => \N__9993\,
            I => \N__9849\
        );

    \I__2316\ : SRMux
    port map (
            O => \N__9992\,
            I => \N__9849\
        );

    \I__2315\ : SRMux
    port map (
            O => \N__9991\,
            I => \N__9849\
        );

    \I__2314\ : SRMux
    port map (
            O => \N__9990\,
            I => \N__9849\
        );

    \I__2313\ : SRMux
    port map (
            O => \N__9989\,
            I => \N__9849\
        );

    \I__2312\ : SRMux
    port map (
            O => \N__9988\,
            I => \N__9849\
        );

    \I__2311\ : SRMux
    port map (
            O => \N__9987\,
            I => \N__9849\
        );

    \I__2310\ : SRMux
    port map (
            O => \N__9986\,
            I => \N__9849\
        );

    \I__2309\ : SRMux
    port map (
            O => \N__9985\,
            I => \N__9849\
        );

    \I__2308\ : SRMux
    port map (
            O => \N__9984\,
            I => \N__9849\
        );

    \I__2307\ : SRMux
    port map (
            O => \N__9983\,
            I => \N__9849\
        );

    \I__2306\ : SRMux
    port map (
            O => \N__9982\,
            I => \N__9849\
        );

    \I__2305\ : SRMux
    port map (
            O => \N__9981\,
            I => \N__9849\
        );

    \I__2304\ : SRMux
    port map (
            O => \N__9980\,
            I => \N__9849\
        );

    \I__2303\ : SRMux
    port map (
            O => \N__9979\,
            I => \N__9849\
        );

    \I__2302\ : SRMux
    port map (
            O => \N__9978\,
            I => \N__9849\
        );

    \I__2301\ : Glb2LocalMux
    port map (
            O => \N__9975\,
            I => \N__9849\
        );

    \I__2300\ : SRMux
    port map (
            O => \N__9974\,
            I => \N__9849\
        );

    \I__2299\ : SRMux
    port map (
            O => \N__9973\,
            I => \N__9849\
        );

    \I__2298\ : SRMux
    port map (
            O => \N__9972\,
            I => \N__9849\
        );

    \I__2297\ : SRMux
    port map (
            O => \N__9971\,
            I => \N__9849\
        );

    \I__2296\ : SRMux
    port map (
            O => \N__9970\,
            I => \N__9849\
        );

    \I__2295\ : SRMux
    port map (
            O => \N__9969\,
            I => \N__9849\
        );

    \I__2294\ : SRMux
    port map (
            O => \N__9968\,
            I => \N__9849\
        );

    \I__2293\ : SRMux
    port map (
            O => \N__9967\,
            I => \N__9849\
        );

    \I__2292\ : SRMux
    port map (
            O => \N__9966\,
            I => \N__9849\
        );

    \I__2291\ : SRMux
    port map (
            O => \N__9965\,
            I => \N__9849\
        );

    \I__2290\ : Glb2LocalMux
    port map (
            O => \N__9962\,
            I => \N__9849\
        );

    \I__2289\ : SRMux
    port map (
            O => \N__9961\,
            I => \N__9849\
        );

    \I__2288\ : SRMux
    port map (
            O => \N__9960\,
            I => \N__9849\
        );

    \I__2287\ : SRMux
    port map (
            O => \N__9959\,
            I => \N__9849\
        );

    \I__2286\ : SRMux
    port map (
            O => \N__9958\,
            I => \N__9849\
        );

    \I__2285\ : Glb2LocalMux
    port map (
            O => \N__9955\,
            I => \N__9849\
        );

    \I__2284\ : SRMux
    port map (
            O => \N__9954\,
            I => \N__9849\
        );

    \I__2283\ : SRMux
    port map (
            O => \N__9953\,
            I => \N__9849\
        );

    \I__2282\ : SRMux
    port map (
            O => \N__9952\,
            I => \N__9849\
        );

    \I__2281\ : SRMux
    port map (
            O => \N__9951\,
            I => \N__9849\
        );

    \I__2280\ : SRMux
    port map (
            O => \N__9950\,
            I => \N__9849\
        );

    \I__2279\ : Glb2LocalMux
    port map (
            O => \N__9947\,
            I => \N__9849\
        );

    \I__2278\ : SRMux
    port map (
            O => \N__9946\,
            I => \N__9849\
        );

    \I__2277\ : SRMux
    port map (
            O => \N__9945\,
            I => \N__9849\
        );

    \I__2276\ : SRMux
    port map (
            O => \N__9944\,
            I => \N__9849\
        );

    \I__2275\ : SRMux
    port map (
            O => \N__9943\,
            I => \N__9849\
        );

    \I__2274\ : SRMux
    port map (
            O => \N__9942\,
            I => \N__9849\
        );

    \I__2273\ : GlobalMux
    port map (
            O => \N__9849\,
            I => \N__9846\
        );

    \I__2272\ : gio2CtrlBuf
    port map (
            O => \N__9846\,
            I => \RESETn_c_i_g\
        );

    \I__2271\ : InMux
    port map (
            O => \N__9843\,
            I => \N__9839\
        );

    \I__2270\ : InMux
    port map (
            O => \N__9842\,
            I => \N__9836\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__9839\,
            I => \N__9833\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__9836\,
            I => \N__9830\
        );

    \I__2267\ : Span12Mux_v
    port map (
            O => \N__9833\,
            I => \N__9826\
        );

    \I__2266\ : Span4Mux_h
    port map (
            O => \N__9830\,
            I => \N__9823\
        );

    \I__2265\ : CascadeMux
    port map (
            O => \N__9829\,
            I => \N__9820\
        );

    \I__2264\ : Span12Mux_h
    port map (
            O => \N__9826\,
            I => \N__9817\
        );

    \I__2263\ : Span4Mux_v
    port map (
            O => \N__9823\,
            I => \N__9814\
        );

    \I__2262\ : InMux
    port map (
            O => \N__9820\,
            I => \N__9811\
        );

    \I__2261\ : Odrv12
    port map (
            O => \N__9817\,
            I => \REG_CYCLEm\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__9814\,
            I => \REG_CYCLEm\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__9811\,
            I => \REG_CYCLEm\
        );

    \I__2258\ : IoInMux
    port map (
            O => \N__9804\,
            I => \N__9801\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__9801\,
            I => \N__9798\
        );

    \I__2256\ : Span12Mux_s6_v
    port map (
            O => \N__9798\,
            I => \N__9795\
        );

    \I__2255\ : Odrv12
    port map (
            O => \N__9795\,
            I => \DRDENn_c\
        );

    \I__2254\ : IoInMux
    port map (
            O => \N__9792\,
            I => \N__9789\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__9789\,
            I => \N__9786\
        );

    \I__2252\ : Span4Mux_s3_v
    port map (
            O => \N__9786\,
            I => \N__9783\
        );

    \I__2251\ : Span4Mux_h
    port map (
            O => \N__9783\,
            I => \N__9780\
        );

    \I__2250\ : Span4Mux_v
    port map (
            O => \N__9780\,
            I => \N__9777\
        );

    \I__2249\ : Odrv4
    port map (
            O => \N__9777\,
            I => \U712_BYTE_ENABLE_un1_UDSn_i\
        );

    \I__2248\ : IoInMux
    port map (
            O => \N__9774\,
            I => \N__9771\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__9771\,
            I => \N__9768\
        );

    \I__2246\ : Span4Mux_s0_v
    port map (
            O => \N__9768\,
            I => \N__9765\
        );

    \I__2245\ : Span4Mux_v
    port map (
            O => \N__9765\,
            I => \N__9762\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__9762\,
            I => \LLBEn_c\
        );

    \I__2243\ : CascadeMux
    port map (
            O => \N__9759\,
            I => \N__9756\
        );

    \I__2242\ : InMux
    port map (
            O => \N__9756\,
            I => \N__9752\
        );

    \I__2241\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9749\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__9752\,
            I => \N__9744\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__9749\,
            I => \N__9744\
        );

    \I__2238\ : Span4Mux_v
    port map (
            O => \N__9744\,
            I => \N__9740\
        );

    \I__2237\ : InMux
    port map (
            O => \N__9743\,
            I => \N__9737\
        );

    \I__2236\ : Odrv4
    port map (
            O => \N__9740\,
            I => \DS_ENm\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__9737\,
            I => \DS_ENm\
        );

    \I__2234\ : IoInMux
    port map (
            O => \N__9732\,
            I => \N__9729\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__9729\,
            I => \N__9726\
        );

    \I__2232\ : Span4Mux_s3_v
    port map (
            O => \N__9726\,
            I => \N__9723\
        );

    \I__2231\ : Span4Mux_h
    port map (
            O => \N__9723\,
            I => \N__9720\
        );

    \I__2230\ : Span4Mux_h
    port map (
            O => \N__9720\,
            I => \N__9717\
        );

    \I__2229\ : Odrv4
    port map (
            O => \N__9717\,
            I => \N_119\
        );

    \I__2228\ : InMux
    port map (
            O => \N__9714\,
            I => \N__9709\
        );

    \I__2227\ : InMux
    port map (
            O => \N__9713\,
            I => \N__9706\
        );

    \I__2226\ : InMux
    port map (
            O => \N__9712\,
            I => \N__9703\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__9709\,
            I => \N__9691\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__9706\,
            I => \N__9691\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__9703\,
            I => \N__9691\
        );

    \I__2222\ : InMux
    port map (
            O => \N__9702\,
            I => \N__9688\
        );

    \I__2221\ : InMux
    port map (
            O => \N__9701\,
            I => \N__9683\
        );

    \I__2220\ : InMux
    port map (
            O => \N__9700\,
            I => \N__9683\
        );

    \I__2219\ : InMux
    port map (
            O => \N__9699\,
            I => \N__9678\
        );

    \I__2218\ : InMux
    port map (
            O => \N__9698\,
            I => \N__9678\
        );

    \I__2217\ : Span4Mux_h
    port map (
            O => \N__9691\,
            I => \N__9673\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__9688\,
            I => \N__9673\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__9683\,
            I => \N__9668\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__9678\,
            I => \N__9668\
        );

    \I__2213\ : Span4Mux_v
    port map (
            O => \N__9673\,
            I => \N__9665\
        );

    \I__2212\ : Span4Mux_v
    port map (
            O => \N__9668\,
            I => \N__9662\
        );

    \I__2211\ : Sp12to4
    port map (
            O => \N__9665\,
            I => \N__9657\
        );

    \I__2210\ : Sp12to4
    port map (
            O => \N__9662\,
            I => \N__9657\
        );

    \I__2209\ : Span12Mux_h
    port map (
            O => \N__9657\,
            I => \N__9654\
        );

    \I__2208\ : Odrv12
    port map (
            O => \N__9654\,
            I => \A_c_1\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__9651\,
            I => \N__9643\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__9650\,
            I => \N__9638\
        );

    \I__2205\ : InMux
    port map (
            O => \N__9649\,
            I => \N__9633\
        );

    \I__2204\ : InMux
    port map (
            O => \N__9648\,
            I => \N__9633\
        );

    \I__2203\ : InMux
    port map (
            O => \N__9647\,
            I => \N__9629\
        );

    \I__2202\ : InMux
    port map (
            O => \N__9646\,
            I => \N__9624\
        );

    \I__2201\ : InMux
    port map (
            O => \N__9643\,
            I => \N__9624\
        );

    \I__2200\ : InMux
    port map (
            O => \N__9642\,
            I => \N__9621\
        );

    \I__2199\ : InMux
    port map (
            O => \N__9641\,
            I => \N__9616\
        );

    \I__2198\ : InMux
    port map (
            O => \N__9638\,
            I => \N__9616\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__9633\,
            I => \N__9613\
        );

    \I__2196\ : InMux
    port map (
            O => \N__9632\,
            I => \N__9610\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__9629\,
            I => \N__9603\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__9624\,
            I => \N__9603\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__9621\,
            I => \N__9603\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__9616\,
            I => \N__9600\
        );

    \I__2191\ : Span4Mux_h
    port map (
            O => \N__9613\,
            I => \N__9597\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__9610\,
            I => \N__9594\
        );

    \I__2189\ : Span4Mux_v
    port map (
            O => \N__9603\,
            I => \N__9590\
        );

    \I__2188\ : Span4Mux_v
    port map (
            O => \N__9600\,
            I => \N__9587\
        );

    \I__2187\ : Span4Mux_v
    port map (
            O => \N__9597\,
            I => \N__9582\
        );

    \I__2186\ : Span4Mux_v
    port map (
            O => \N__9594\,
            I => \N__9582\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9593\,
            I => \N__9579\
        );

    \I__2184\ : Sp12to4
    port map (
            O => \N__9590\,
            I => \N__9570\
        );

    \I__2183\ : Sp12to4
    port map (
            O => \N__9587\,
            I => \N__9570\
        );

    \I__2182\ : Sp12to4
    port map (
            O => \N__9582\,
            I => \N__9570\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__9579\,
            I => \N__9570\
        );

    \I__2180\ : Span12Mux_h
    port map (
            O => \N__9570\,
            I => \N__9567\
        );

    \I__2179\ : Odrv12
    port map (
            O => \N__9567\,
            I => \A_c_0\
        );

    \I__2178\ : CascadeMux
    port map (
            O => \N__9564\,
            I => \N__9560\
        );

    \I__2177\ : InMux
    port map (
            O => \N__9563\,
            I => \N__9552\
        );

    \I__2176\ : InMux
    port map (
            O => \N__9560\,
            I => \N__9552\
        );

    \I__2175\ : InMux
    port map (
            O => \N__9559\,
            I => \N__9547\
        );

    \I__2174\ : InMux
    port map (
            O => \N__9558\,
            I => \N__9547\
        );

    \I__2173\ : CascadeMux
    port map (
            O => \N__9557\,
            I => \N__9543\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__9552\,
            I => \N__9539\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__9547\,
            I => \N__9536\
        );

    \I__2170\ : InMux
    port map (
            O => \N__9546\,
            I => \N__9529\
        );

    \I__2169\ : InMux
    port map (
            O => \N__9543\,
            I => \N__9529\
        );

    \I__2168\ : InMux
    port map (
            O => \N__9542\,
            I => \N__9529\
        );

    \I__2167\ : Span4Mux_v
    port map (
            O => \N__9539\,
            I => \N__9525\
        );

    \I__2166\ : Span4Mux_v
    port map (
            O => \N__9536\,
            I => \N__9522\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__9529\,
            I => \N__9519\
        );

    \I__2164\ : CascadeMux
    port map (
            O => \N__9528\,
            I => \N__9516\
        );

    \I__2163\ : Span4Mux_v
    port map (
            O => \N__9525\,
            I => \N__9513\
        );

    \I__2162\ : Span4Mux_v
    port map (
            O => \N__9522\,
            I => \N__9508\
        );

    \I__2161\ : Span4Mux_h
    port map (
            O => \N__9519\,
            I => \N__9508\
        );

    \I__2160\ : InMux
    port map (
            O => \N__9516\,
            I => \N__9505\
        );

    \I__2159\ : Span4Mux_v
    port map (
            O => \N__9513\,
            I => \N__9502\
        );

    \I__2158\ : Span4Mux_v
    port map (
            O => \N__9508\,
            I => \N__9499\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__9505\,
            I => \N__9496\
        );

    \I__2156\ : Sp12to4
    port map (
            O => \N__9502\,
            I => \N__9489\
        );

    \I__2155\ : Sp12to4
    port map (
            O => \N__9499\,
            I => \N__9489\
        );

    \I__2154\ : Span12Mux_v
    port map (
            O => \N__9496\,
            I => \N__9489\
        );

    \I__2153\ : Span12Mux_h
    port map (
            O => \N__9489\,
            I => \N__9486\
        );

    \I__2152\ : Odrv12
    port map (
            O => \N__9486\,
            I => \SIZ_c_1\
        );

    \I__2151\ : InMux
    port map (
            O => \N__9483\,
            I => \N__9476\
        );

    \I__2150\ : InMux
    port map (
            O => \N__9482\,
            I => \N__9473\
        );

    \I__2149\ : InMux
    port map (
            O => \N__9481\,
            I => \N__9466\
        );

    \I__2148\ : InMux
    port map (
            O => \N__9480\,
            I => \N__9466\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9479\,
            I => \N__9466\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__9476\,
            I => \N__9462\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__9473\,
            I => \N__9459\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__9466\,
            I => \N__9456\
        );

    \I__2143\ : InMux
    port map (
            O => \N__9465\,
            I => \N__9453\
        );

    \I__2142\ : Span4Mux_v
    port map (
            O => \N__9462\,
            I => \N__9450\
        );

    \I__2141\ : Span4Mux_v
    port map (
            O => \N__9459\,
            I => \N__9447\
        );

    \I__2140\ : Span4Mux_h
    port map (
            O => \N__9456\,
            I => \N__9442\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__9453\,
            I => \N__9442\
        );

    \I__2138\ : Span4Mux_v
    port map (
            O => \N__9450\,
            I => \N__9439\
        );

    \I__2137\ : Span4Mux_v
    port map (
            O => \N__9447\,
            I => \N__9434\
        );

    \I__2136\ : Span4Mux_h
    port map (
            O => \N__9442\,
            I => \N__9434\
        );

    \I__2135\ : Span4Mux_v
    port map (
            O => \N__9439\,
            I => \N__9431\
        );

    \I__2134\ : Span4Mux_v
    port map (
            O => \N__9434\,
            I => \N__9428\
        );

    \I__2133\ : Span4Mux_h
    port map (
            O => \N__9431\,
            I => \N__9425\
        );

    \I__2132\ : Span4Mux_h
    port map (
            O => \N__9428\,
            I => \N__9422\
        );

    \I__2131\ : Sp12to4
    port map (
            O => \N__9425\,
            I => \N__9417\
        );

    \I__2130\ : Sp12to4
    port map (
            O => \N__9422\,
            I => \N__9417\
        );

    \I__2129\ : Odrv12
    port map (
            O => \N__9417\,
            I => \SIZ_c_0\
        );

    \I__2128\ : IoInMux
    port map (
            O => \N__9414\,
            I => \N__9411\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__9411\,
            I => \N__9408\
        );

    \I__2126\ : Span4Mux_s3_v
    port map (
            O => \N__9408\,
            I => \N__9405\
        );

    \I__2125\ : Odrv4
    port map (
            O => \N__9405\,
            I => \N_220_i\
        );

    \I__2124\ : CascadeMux
    port map (
            O => \N__9402\,
            I => \N__9393\
        );

    \I__2123\ : InMux
    port map (
            O => \N__9401\,
            I => \N__9389\
        );

    \I__2122\ : InMux
    port map (
            O => \N__9400\,
            I => \N__9384\
        );

    \I__2121\ : InMux
    port map (
            O => \N__9399\,
            I => \N__9384\
        );

    \I__2120\ : InMux
    port map (
            O => \N__9398\,
            I => \N__9381\
        );

    \I__2119\ : InMux
    port map (
            O => \N__9397\,
            I => \N__9374\
        );

    \I__2118\ : InMux
    port map (
            O => \N__9396\,
            I => \N__9374\
        );

    \I__2117\ : InMux
    port map (
            O => \N__9393\,
            I => \N__9371\
        );

    \I__2116\ : InMux
    port map (
            O => \N__9392\,
            I => \N__9367\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__9389\,
            I => \N__9364\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__9384\,
            I => \N__9353\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__9381\,
            I => \N__9350\
        );

    \I__2112\ : CascadeMux
    port map (
            O => \N__9380\,
            I => \N__9347\
        );

    \I__2111\ : CascadeMux
    port map (
            O => \N__9379\,
            I => \N__9344\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__9374\,
            I => \N__9337\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__9371\,
            I => \N__9337\
        );

    \I__2108\ : InMux
    port map (
            O => \N__9370\,
            I => \N__9334\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__9367\,
            I => \N__9327\
        );

    \I__2106\ : Span4Mux_v
    port map (
            O => \N__9364\,
            I => \N__9327\
        );

    \I__2105\ : InMux
    port map (
            O => \N__9363\,
            I => \N__9324\
        );

    \I__2104\ : InMux
    port map (
            O => \N__9362\,
            I => \N__9321\
        );

    \I__2103\ : InMux
    port map (
            O => \N__9361\,
            I => \N__9317\
        );

    \I__2102\ : InMux
    port map (
            O => \N__9360\,
            I => \N__9310\
        );

    \I__2101\ : InMux
    port map (
            O => \N__9359\,
            I => \N__9310\
        );

    \I__2100\ : InMux
    port map (
            O => \N__9358\,
            I => \N__9310\
        );

    \I__2099\ : InMux
    port map (
            O => \N__9357\,
            I => \N__9305\
        );

    \I__2098\ : InMux
    port map (
            O => \N__9356\,
            I => \N__9305\
        );

    \I__2097\ : Span4Mux_v
    port map (
            O => \N__9353\,
            I => \N__9300\
        );

    \I__2096\ : Span4Mux_v
    port map (
            O => \N__9350\,
            I => \N__9300\
        );

    \I__2095\ : InMux
    port map (
            O => \N__9347\,
            I => \N__9291\
        );

    \I__2094\ : InMux
    port map (
            O => \N__9344\,
            I => \N__9291\
        );

    \I__2093\ : InMux
    port map (
            O => \N__9343\,
            I => \N__9291\
        );

    \I__2092\ : InMux
    port map (
            O => \N__9342\,
            I => \N__9291\
        );

    \I__2091\ : Span4Mux_v
    port map (
            O => \N__9337\,
            I => \N__9288\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__9334\,
            I => \N__9285\
        );

    \I__2089\ : InMux
    port map (
            O => \N__9333\,
            I => \N__9280\
        );

    \I__2088\ : InMux
    port map (
            O => \N__9332\,
            I => \N__9280\
        );

    \I__2087\ : Span4Mux_h
    port map (
            O => \N__9327\,
            I => \N__9273\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__9324\,
            I => \N__9273\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__9321\,
            I => \N__9273\
        );

    \I__2084\ : InMux
    port map (
            O => \N__9320\,
            I => \N__9270\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__9317\,
            I => \N__9267\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__9310\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__9305\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2080\ : Odrv4
    port map (
            O => \N__9300\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__9291\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__9288\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2077\ : Odrv4
    port map (
            O => \N__9285\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__9280\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2075\ : Odrv4
    port map (
            O => \N__9273\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__9270\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2073\ : Odrv4
    port map (
            O => \N__9267\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2072\ : IoInMux
    port map (
            O => \N__9246\,
            I => \N__9243\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__9243\,
            I => \N__9240\
        );

    \I__2070\ : Span4Mux_s2_v
    port map (
            O => \N__9240\,
            I => \N__9237\
        );

    \I__2069\ : Span4Mux_v
    port map (
            O => \N__9237\,
            I => \N__9234\
        );

    \I__2068\ : Span4Mux_v
    port map (
            O => \N__9234\,
            I => \N__9231\
        );

    \I__2067\ : Span4Mux_h
    port map (
            O => \N__9231\,
            I => \N__9228\
        );

    \I__2066\ : Odrv4
    port map (
            O => \N__9228\,
            I => \CASn_c\
        );

    \I__2065\ : InMux
    port map (
            O => \N__9225\,
            I => \N__9222\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__9222\,
            I => \N__9219\
        );

    \I__2063\ : Span12Mux_h
    port map (
            O => \N__9219\,
            I => \N__9216\
        );

    \I__2062\ : Odrv12
    port map (
            O => \N__9216\,
            I => \RAS0n_c\
        );

    \I__2061\ : InMux
    port map (
            O => \N__9213\,
            I => \N__9209\
        );

    \I__2060\ : InMux
    port map (
            O => \N__9212\,
            I => \N__9204\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__9209\,
            I => \N__9201\
        );

    \I__2058\ : InMux
    port map (
            O => \N__9208\,
            I => \N__9198\
        );

    \I__2057\ : InMux
    port map (
            O => \N__9207\,
            I => \N__9195\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__9204\,
            I => \N__9192\
        );

    \I__2055\ : Span4Mux_h
    port map (
            O => \N__9201\,
            I => \N__9185\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__9198\,
            I => \N__9185\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__9195\,
            I => \N__9185\
        );

    \I__2052\ : Span4Mux_h
    port map (
            O => \N__9192\,
            I => \N__9182\
        );

    \I__2051\ : Span4Mux_h
    port map (
            O => \N__9185\,
            I => \N__9179\
        );

    \I__2050\ : Sp12to4
    port map (
            O => \N__9182\,
            I => \N__9176\
        );

    \I__2049\ : Span4Mux_v
    port map (
            O => \N__9179\,
            I => \N__9173\
        );

    \I__2048\ : Span12Mux_v
    port map (
            O => \N__9176\,
            I => \N__9170\
        );

    \I__2047\ : Sp12to4
    port map (
            O => \N__9173\,
            I => \N__9167\
        );

    \I__2046\ : Span12Mux_h
    port map (
            O => \N__9170\,
            I => \N__9164\
        );

    \I__2045\ : Span12Mux_v
    port map (
            O => \N__9167\,
            I => \N__9161\
        );

    \I__2044\ : Odrv12
    port map (
            O => \N__9164\,
            I => \DRA_c_9\
        );

    \I__2043\ : Odrv12
    port map (
            O => \N__9161\,
            I => \DRA_c_9\
        );

    \I__2042\ : InMux
    port map (
            O => \N__9156\,
            I => \N__9153\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__9153\,
            I => \N__9150\
        );

    \I__2040\ : Span4Mux_v
    port map (
            O => \N__9150\,
            I => \N__9147\
        );

    \I__2039\ : Odrv4
    port map (
            O => \N__9147\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2038\ : InMux
    port map (
            O => \N__9144\,
            I => \N__9141\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__9141\,
            I => \N__9136\
        );

    \I__2036\ : InMux
    port map (
            O => \N__9140\,
            I => \N__9133\
        );

    \I__2035\ : InMux
    port map (
            O => \N__9139\,
            I => \N__9130\
        );

    \I__2034\ : Span4Mux_v
    port map (
            O => \N__9136\,
            I => \N__9126\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__9133\,
            I => \N__9123\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__9130\,
            I => \N__9120\
        );

    \I__2031\ : InMux
    port map (
            O => \N__9129\,
            I => \N__9117\
        );

    \I__2030\ : Sp12to4
    port map (
            O => \N__9126\,
            I => \N__9108\
        );

    \I__2029\ : Span12Mux_v
    port map (
            O => \N__9123\,
            I => \N__9108\
        );

    \I__2028\ : Span12Mux_v
    port map (
            O => \N__9120\,
            I => \N__9108\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__9117\,
            I => \N__9108\
        );

    \I__2026\ : Span12Mux_h
    port map (
            O => \N__9108\,
            I => \N__9105\
        );

    \I__2025\ : Odrv12
    port map (
            O => \N__9105\,
            I => \DRA_c_8\
        );

    \I__2024\ : InMux
    port map (
            O => \N__9102\,
            I => \N__9099\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__9099\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2022\ : InMux
    port map (
            O => \N__9096\,
            I => \N__9093\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__9093\,
            I => \N__9090\
        );

    \I__2020\ : Odrv4
    port map (
            O => \N__9090\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__2019\ : IoInMux
    port map (
            O => \N__9087\,
            I => \N__9084\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__9084\,
            I => \N__9081\
        );

    \I__2017\ : Span12Mux_s5_h
    port map (
            O => \N__9081\,
            I => \N__9078\
        );

    \I__2016\ : Span12Mux_v
    port map (
            O => \N__9078\,
            I => \N__9075\
        );

    \I__2015\ : Odrv12
    port map (
            O => \N__9075\,
            I => \CMA_c_6\
        );

    \I__2014\ : InMux
    port map (
            O => \N__9072\,
            I => \N__9069\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__9069\,
            I => \N__9066\
        );

    \I__2012\ : Odrv12
    port map (
            O => \N__9066\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__2011\ : IoInMux
    port map (
            O => \N__9063\,
            I => \N__9060\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__9060\,
            I => \N__9057\
        );

    \I__2009\ : Span4Mux_s3_v
    port map (
            O => \N__9057\,
            I => \N__9054\
        );

    \I__2008\ : Odrv4
    port map (
            O => \N__9054\,
            I => \U712_BYTE_ENABLE_UUBE_i\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__9051\,
            I => \N__9047\
        );

    \I__2006\ : InMux
    port map (
            O => \N__9050\,
            I => \N__9044\
        );

    \I__2005\ : InMux
    port map (
            O => \N__9047\,
            I => \N__9041\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__9044\,
            I => \N__9038\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__9041\,
            I => \N__9034\
        );

    \I__2002\ : Span4Mux_h
    port map (
            O => \N__9038\,
            I => \N__9031\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__9037\,
            I => \N__9026\
        );

    \I__2000\ : Span4Mux_v
    port map (
            O => \N__9034\,
            I => \N__9023\
        );

    \I__1999\ : Span4Mux_v
    port map (
            O => \N__9031\,
            I => \N__9020\
        );

    \I__1998\ : InMux
    port map (
            O => \N__9030\,
            I => \N__9015\
        );

    \I__1997\ : InMux
    port map (
            O => \N__9029\,
            I => \N__9015\
        );

    \I__1996\ : InMux
    port map (
            O => \N__9026\,
            I => \N__9012\
        );

    \I__1995\ : Odrv4
    port map (
            O => \N__9023\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1994\ : Odrv4
    port map (
            O => \N__9020\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__9015\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__9012\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1991\ : IoInMux
    port map (
            O => \N__9003\,
            I => \N__9000\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__9000\,
            I => \N__8997\
        );

    \I__1989\ : Span4Mux_s3_v
    port map (
            O => \N__8997\,
            I => \N__8994\
        );

    \I__1988\ : Span4Mux_v
    port map (
            O => \N__8994\,
            I => \N__8991\
        );

    \I__1987\ : Span4Mux_h
    port map (
            O => \N__8991\,
            I => \N__8988\
        );

    \I__1986\ : Odrv4
    port map (
            O => \N__8988\,
            I => \CRCSn_c\
        );

    \I__1985\ : InMux
    port map (
            O => \N__8985\,
            I => \N__8982\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__8982\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__1983\ : IoInMux
    port map (
            O => \N__8979\,
            I => \N__8976\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__8976\,
            I => \N__8973\
        );

    \I__1981\ : IoSpan4Mux
    port map (
            O => \N__8973\,
            I => \N__8970\
        );

    \I__1980\ : Span4Mux_s0_h
    port map (
            O => \N__8970\,
            I => \N__8967\
        );

    \I__1979\ : Sp12to4
    port map (
            O => \N__8967\,
            I => \N__8964\
        );

    \I__1978\ : Span12Mux_h
    port map (
            O => \N__8964\,
            I => \N__8961\
        );

    \I__1977\ : Odrv12
    port map (
            O => \N__8961\,
            I => \CMA_c_7\
        );

    \I__1976\ : InMux
    port map (
            O => \N__8958\,
            I => \N__8955\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__8955\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__1974\ : IoInMux
    port map (
            O => \N__8952\,
            I => \N__8949\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__8949\,
            I => \N__8946\
        );

    \I__1972\ : Span12Mux_s5_h
    port map (
            O => \N__8946\,
            I => \N__8943\
        );

    \I__1971\ : Span12Mux_v
    port map (
            O => \N__8943\,
            I => \N__8940\
        );

    \I__1970\ : Odrv12
    port map (
            O => \N__8940\,
            I => \CMA_c_4\
        );

    \I__1969\ : InMux
    port map (
            O => \N__8937\,
            I => \N__8934\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__8934\,
            I => \N__8931\
        );

    \I__1967\ : Span4Mux_h
    port map (
            O => \N__8931\,
            I => \N__8928\
        );

    \I__1966\ : Span4Mux_h
    port map (
            O => \N__8928\,
            I => \N__8925\
        );

    \I__1965\ : Odrv4
    port map (
            O => \N__8925\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__1964\ : InMux
    port map (
            O => \N__8922\,
            I => \N__8919\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__8919\,
            I => \N__8916\
        );

    \I__1962\ : Odrv12
    port map (
            O => \N__8916\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__1961\ : InMux
    port map (
            O => \N__8913\,
            I => \N__8910\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__8910\,
            I => \N__8907\
        );

    \I__1959\ : Span4Mux_h
    port map (
            O => \N__8907\,
            I => \N__8904\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__8904\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__1957\ : InMux
    port map (
            O => \N__8901\,
            I => \N__8894\
        );

    \I__1956\ : InMux
    port map (
            O => \N__8900\,
            I => \N__8894\
        );

    \I__1955\ : InMux
    port map (
            O => \N__8899\,
            I => \N__8891\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__8894\,
            I => \N__8885\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__8891\,
            I => \N__8885\
        );

    \I__1952\ : InMux
    port map (
            O => \N__8890\,
            I => \N__8882\
        );

    \I__1951\ : Span4Mux_v
    port map (
            O => \N__8885\,
            I => \N__8877\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__8882\,
            I => \N__8877\
        );

    \I__1949\ : Span4Mux_h
    port map (
            O => \N__8877\,
            I => \N__8874\
        );

    \I__1948\ : Span4Mux_v
    port map (
            O => \N__8874\,
            I => \N__8871\
        );

    \I__1947\ : Sp12to4
    port map (
            O => \N__8871\,
            I => \N__8868\
        );

    \I__1946\ : Odrv12
    port map (
            O => \N__8868\,
            I => \DRA_c_2\
        );

    \I__1945\ : InMux
    port map (
            O => \N__8865\,
            I => \N__8862\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__8862\,
            I => \N__8859\
        );

    \I__1943\ : Span4Mux_h
    port map (
            O => \N__8859\,
            I => \N__8856\
        );

    \I__1942\ : Odrv4
    port map (
            O => \N__8856\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__8853\,
            I => \N__8850\
        );

    \I__1940\ : InMux
    port map (
            O => \N__8850\,
            I => \N__8842\
        );

    \I__1939\ : InMux
    port map (
            O => \N__8849\,
            I => \N__8842\
        );

    \I__1938\ : InMux
    port map (
            O => \N__8848\,
            I => \N__8837\
        );

    \I__1937\ : InMux
    port map (
            O => \N__8847\,
            I => \N__8837\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__8842\,
            I => \N__8831\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__8837\,
            I => \N__8831\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__8836\,
            I => \N__8827\
        );

    \I__1933\ : Span4Mux_h
    port map (
            O => \N__8831\,
            I => \N__8817\
        );

    \I__1932\ : InMux
    port map (
            O => \N__8830\,
            I => \N__8814\
        );

    \I__1931\ : InMux
    port map (
            O => \N__8827\,
            I => \N__8811\
        );

    \I__1930\ : InMux
    port map (
            O => \N__8826\,
            I => \N__8806\
        );

    \I__1929\ : InMux
    port map (
            O => \N__8825\,
            I => \N__8803\
        );

    \I__1928\ : InMux
    port map (
            O => \N__8824\,
            I => \N__8800\
        );

    \I__1927\ : InMux
    port map (
            O => \N__8823\,
            I => \N__8795\
        );

    \I__1926\ : InMux
    port map (
            O => \N__8822\,
            I => \N__8795\
        );

    \I__1925\ : InMux
    port map (
            O => \N__8821\,
            I => \N__8789\
        );

    \I__1924\ : InMux
    port map (
            O => \N__8820\,
            I => \N__8784\
        );

    \I__1923\ : Span4Mux_v
    port map (
            O => \N__8817\,
            I => \N__8779\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__8814\,
            I => \N__8779\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__8811\,
            I => \N__8770\
        );

    \I__1920\ : InMux
    port map (
            O => \N__8810\,
            I => \N__8765\
        );

    \I__1919\ : InMux
    port map (
            O => \N__8809\,
            I => \N__8765\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__8806\,
            I => \N__8762\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__8803\,
            I => \N__8759\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__8800\,
            I => \N__8754\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__8795\,
            I => \N__8754\
        );

    \I__1914\ : InMux
    port map (
            O => \N__8794\,
            I => \N__8747\
        );

    \I__1913\ : InMux
    port map (
            O => \N__8793\,
            I => \N__8747\
        );

    \I__1912\ : InMux
    port map (
            O => \N__8792\,
            I => \N__8747\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__8789\,
            I => \N__8744\
        );

    \I__1910\ : InMux
    port map (
            O => \N__8788\,
            I => \N__8741\
        );

    \I__1909\ : InMux
    port map (
            O => \N__8787\,
            I => \N__8738\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8784\,
            I => \N__8735\
        );

    \I__1907\ : Span4Mux_h
    port map (
            O => \N__8779\,
            I => \N__8732\
        );

    \I__1906\ : InMux
    port map (
            O => \N__8778\,
            I => \N__8727\
        );

    \I__1905\ : InMux
    port map (
            O => \N__8777\,
            I => \N__8727\
        );

    \I__1904\ : InMux
    port map (
            O => \N__8776\,
            I => \N__8718\
        );

    \I__1903\ : InMux
    port map (
            O => \N__8775\,
            I => \N__8718\
        );

    \I__1902\ : InMux
    port map (
            O => \N__8774\,
            I => \N__8718\
        );

    \I__1901\ : InMux
    port map (
            O => \N__8773\,
            I => \N__8718\
        );

    \I__1900\ : Span4Mux_v
    port map (
            O => \N__8770\,
            I => \N__8709\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__8765\,
            I => \N__8709\
        );

    \I__1898\ : Span4Mux_v
    port map (
            O => \N__8762\,
            I => \N__8709\
        );

    \I__1897\ : Span4Mux_v
    port map (
            O => \N__8759\,
            I => \N__8709\
        );

    \I__1896\ : Span12Mux_v
    port map (
            O => \N__8754\,
            I => \N__8704\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__8747\,
            I => \N__8704\
        );

    \I__1894\ : Odrv4
    port map (
            O => \N__8744\,
            I => \CPU_CYCLEm\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__8741\,
            I => \CPU_CYCLEm\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__8738\,
            I => \CPU_CYCLEm\
        );

    \I__1891\ : Odrv4
    port map (
            O => \N__8735\,
            I => \CPU_CYCLEm\
        );

    \I__1890\ : Odrv4
    port map (
            O => \N__8732\,
            I => \CPU_CYCLEm\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__8727\,
            I => \CPU_CYCLEm\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__8718\,
            I => \CPU_CYCLEm\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__8709\,
            I => \CPU_CYCLEm\
        );

    \I__1886\ : Odrv12
    port map (
            O => \N__8704\,
            I => \CPU_CYCLEm\
        );

    \I__1885\ : CascadeMux
    port map (
            O => \N__8685\,
            I => \N__8682\
        );

    \I__1884\ : InMux
    port map (
            O => \N__8682\,
            I => \N__8679\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__8679\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__1882\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8673\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__8673\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__1880\ : InMux
    port map (
            O => \N__8670\,
            I => \N__8667\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__8667\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1878\ : InMux
    port map (
            O => \N__8664\,
            I => \N__8661\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8661\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__1876\ : InMux
    port map (
            O => \N__8658\,
            I => \N__8655\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__8655\,
            I => \N__8652\
        );

    \I__1874\ : Span4Mux_v
    port map (
            O => \N__8652\,
            I => \N__8649\
        );

    \I__1873\ : Odrv4
    port map (
            O => \N__8649\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__1872\ : InMux
    port map (
            O => \N__8646\,
            I => \N__8643\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__8643\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1870\ : InMux
    port map (
            O => \N__8640\,
            I => \N__8634\
        );

    \I__1869\ : InMux
    port map (
            O => \N__8639\,
            I => \N__8634\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__8634\,
            I => \N__8631\
        );

    \I__1867\ : Span4Mux_h
    port map (
            O => \N__8631\,
            I => \N__8628\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__8628\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__1865\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8622\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__8622\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__1863\ : InMux
    port map (
            O => \N__8619\,
            I => \N__8615\
        );

    \I__1862\ : InMux
    port map (
            O => \N__8618\,
            I => \N__8610\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__8615\,
            I => \N__8607\
        );

    \I__1860\ : InMux
    port map (
            O => \N__8614\,
            I => \N__8604\
        );

    \I__1859\ : InMux
    port map (
            O => \N__8613\,
            I => \N__8601\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__8610\,
            I => \N__8598\
        );

    \I__1857\ : Span4Mux_h
    port map (
            O => \N__8607\,
            I => \N__8591\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__8604\,
            I => \N__8591\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__8601\,
            I => \N__8591\
        );

    \I__1854\ : Span4Mux_h
    port map (
            O => \N__8598\,
            I => \N__8586\
        );

    \I__1853\ : Span4Mux_h
    port map (
            O => \N__8591\,
            I => \N__8586\
        );

    \I__1852\ : Span4Mux_v
    port map (
            O => \N__8586\,
            I => \N__8583\
        );

    \I__1851\ : Span4Mux_v
    port map (
            O => \N__8583\,
            I => \N__8580\
        );

    \I__1850\ : Span4Mux_v
    port map (
            O => \N__8580\,
            I => \N__8577\
        );

    \I__1849\ : Span4Mux_v
    port map (
            O => \N__8577\,
            I => \N__8574\
        );

    \I__1848\ : Odrv4
    port map (
            O => \N__8574\,
            I => \CLK40_PLL_i\
        );

    \I__1847\ : IoInMux
    port map (
            O => \N__8571\,
            I => \N__8566\
        );

    \I__1846\ : IoInMux
    port map (
            O => \N__8570\,
            I => \N__8563\
        );

    \I__1845\ : IoInMux
    port map (
            O => \N__8569\,
            I => \N__8560\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__8566\,
            I => \N__8557\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__8563\,
            I => \N__8554\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__8560\,
            I => \N__8551\
        );

    \I__1841\ : IoSpan4Mux
    port map (
            O => \N__8557\,
            I => \N__8548\
        );

    \I__1840\ : Span4Mux_s3_v
    port map (
            O => \N__8554\,
            I => \N__8545\
        );

    \I__1839\ : Span4Mux_s2_h
    port map (
            O => \N__8551\,
            I => \N__8542\
        );

    \I__1838\ : IoSpan4Mux
    port map (
            O => \N__8548\,
            I => \N__8539\
        );

    \I__1837\ : Span4Mux_h
    port map (
            O => \N__8545\,
            I => \N__8536\
        );

    \I__1836\ : Span4Mux_v
    port map (
            O => \N__8542\,
            I => \N__8533\
        );

    \I__1835\ : Sp12to4
    port map (
            O => \N__8539\,
            I => \N__8528\
        );

    \I__1834\ : Sp12to4
    port map (
            O => \N__8536\,
            I => \N__8528\
        );

    \I__1833\ : Sp12to4
    port map (
            O => \N__8533\,
            I => \N__8525\
        );

    \I__1832\ : Span12Mux_v
    port map (
            O => \N__8528\,
            I => \N__8520\
        );

    \I__1831\ : Span12Mux_h
    port map (
            O => \N__8525\,
            I => \N__8520\
        );

    \I__1830\ : Odrv12
    port map (
            O => \N__8520\,
            I => \CLK40_PLL_i_i\
        );

    \I__1829\ : IoInMux
    port map (
            O => \N__8517\,
            I => \N__8514\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__8514\,
            I => \N__8511\
        );

    \I__1827\ : Span4Mux_s2_v
    port map (
            O => \N__8511\,
            I => \N__8508\
        );

    \I__1826\ : Span4Mux_h
    port map (
            O => \N__8508\,
            I => \N__8505\
        );

    \I__1825\ : Span4Mux_v
    port map (
            O => \N__8505\,
            I => \N__8502\
        );

    \I__1824\ : Odrv4
    port map (
            O => \N__8502\,
            I => \UMBEn_c\
        );

    \I__1823\ : CascadeMux
    port map (
            O => \N__8499\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8496\,
            I => \N__8493\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__8493\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i\
        );

    \I__1820\ : InMux
    port map (
            O => \N__8490\,
            I => \N__8487\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__8487\,
            I => \N__8483\
        );

    \I__1818\ : InMux
    port map (
            O => \N__8486\,
            I => \N__8475\
        );

    \I__1817\ : Span4Mux_h
    port map (
            O => \N__8483\,
            I => \N__8472\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8482\,
            I => \N__8465\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8481\,
            I => \N__8465\
        );

    \I__1814\ : InMux
    port map (
            O => \N__8480\,
            I => \N__8465\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8479\,
            I => \N__8460\
        );

    \I__1812\ : InMux
    port map (
            O => \N__8478\,
            I => \N__8460\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__8475\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1810\ : Odrv4
    port map (
            O => \N__8472\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__8465\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__8460\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1807\ : InMux
    port map (
            O => \N__8451\,
            I => \N__8448\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__8448\,
            I => \N__8444\
        );

    \I__1805\ : InMux
    port map (
            O => \N__8447\,
            I => \N__8441\
        );

    \I__1804\ : Span4Mux_h
    port map (
            O => \N__8444\,
            I => \N__8436\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__8441\,
            I => \N__8436\
        );

    \I__1802\ : Span4Mux_h
    port map (
            O => \N__8436\,
            I => \N__8431\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8435\,
            I => \N__8426\
        );

    \I__1800\ : InMux
    port map (
            O => \N__8434\,
            I => \N__8426\
        );

    \I__1799\ : Odrv4
    port map (
            O => \N__8431\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__8426\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__8421\,
            I => \U712_REG_SM.N_236_cascade_\
        );

    \I__1796\ : CascadeMux
    port map (
            O => \N__8418\,
            I => \N__8415\
        );

    \I__1795\ : InMux
    port map (
            O => \N__8415\,
            I => \N__8409\
        );

    \I__1794\ : InMux
    port map (
            O => \N__8414\,
            I => \N__8404\
        );

    \I__1793\ : InMux
    port map (
            O => \N__8413\,
            I => \N__8404\
        );

    \I__1792\ : InMux
    port map (
            O => \N__8412\,
            I => \N__8401\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__8409\,
            I => \N__8389\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__8404\,
            I => \N__8389\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__8401\,
            I => \N__8386\
        );

    \I__1788\ : InMux
    port map (
            O => \N__8400\,
            I => \N__8379\
        );

    \I__1787\ : InMux
    port map (
            O => \N__8399\,
            I => \N__8379\
        );

    \I__1786\ : InMux
    port map (
            O => \N__8398\,
            I => \N__8379\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8397\,
            I => \N__8376\
        );

    \I__1784\ : InMux
    port map (
            O => \N__8396\,
            I => \N__8373\
        );

    \I__1783\ : InMux
    port map (
            O => \N__8395\,
            I => \N__8368\
        );

    \I__1782\ : InMux
    port map (
            O => \N__8394\,
            I => \N__8368\
        );

    \I__1781\ : Span4Mux_h
    port map (
            O => \N__8389\,
            I => \N__8365\
        );

    \I__1780\ : Odrv4
    port map (
            O => \N__8386\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__8379\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__8376\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__8373\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__8368\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1775\ : Odrv4
    port map (
            O => \N__8365\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__8352\,
            I => \N__8348\
        );

    \I__1773\ : CascadeMux
    port map (
            O => \N__8351\,
            I => \N__8343\
        );

    \I__1772\ : InMux
    port map (
            O => \N__8348\,
            I => \N__8338\
        );

    \I__1771\ : InMux
    port map (
            O => \N__8347\,
            I => \N__8335\
        );

    \I__1770\ : InMux
    port map (
            O => \N__8346\,
            I => \N__8332\
        );

    \I__1769\ : InMux
    port map (
            O => \N__8343\,
            I => \N__8327\
        );

    \I__1768\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8327\
        );

    \I__1767\ : InMux
    port map (
            O => \N__8341\,
            I => \N__8324\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__8338\,
            I => \N__8317\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__8335\,
            I => \N__8317\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8332\,
            I => \N__8317\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__8327\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__8324\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1761\ : Odrv12
    port map (
            O => \N__8317\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1760\ : CascadeMux
    port map (
            O => \N__8310\,
            I => \N__8297\
        );

    \I__1759\ : InMux
    port map (
            O => \N__8309\,
            I => \N__8291\
        );

    \I__1758\ : InMux
    port map (
            O => \N__8308\,
            I => \N__8291\
        );

    \I__1757\ : CascadeMux
    port map (
            O => \N__8307\,
            I => \N__8288\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__8306\,
            I => \N__8285\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8305\,
            I => \N__8282\
        );

    \I__1754\ : InMux
    port map (
            O => \N__8304\,
            I => \N__8277\
        );

    \I__1753\ : InMux
    port map (
            O => \N__8303\,
            I => \N__8277\
        );

    \I__1752\ : InMux
    port map (
            O => \N__8302\,
            I => \N__8273\
        );

    \I__1751\ : InMux
    port map (
            O => \N__8301\,
            I => \N__8264\
        );

    \I__1750\ : InMux
    port map (
            O => \N__8300\,
            I => \N__8264\
        );

    \I__1749\ : InMux
    port map (
            O => \N__8297\,
            I => \N__8264\
        );

    \I__1748\ : InMux
    port map (
            O => \N__8296\,
            I => \N__8264\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__8291\,
            I => \N__8261\
        );

    \I__1746\ : InMux
    port map (
            O => \N__8288\,
            I => \N__8258\
        );

    \I__1745\ : InMux
    port map (
            O => \N__8285\,
            I => \N__8255\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__8282\,
            I => \N__8250\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__8277\,
            I => \N__8250\
        );

    \I__1742\ : InMux
    port map (
            O => \N__8276\,
            I => \N__8247\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__8273\,
            I => \N__8242\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__8264\,
            I => \N__8242\
        );

    \I__1739\ : Span4Mux_v
    port map (
            O => \N__8261\,
            I => \N__8239\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__8258\,
            I => \N__8232\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__8255\,
            I => \N__8232\
        );

    \I__1736\ : Span4Mux_v
    port map (
            O => \N__8250\,
            I => \N__8232\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__8247\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1734\ : Odrv4
    port map (
            O => \N__8242\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1733\ : Odrv4
    port map (
            O => \N__8239\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1732\ : Odrv4
    port map (
            O => \N__8232\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1731\ : InMux
    port map (
            O => \N__8223\,
            I => \N__8220\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__8220\,
            I => \U712_REG_SM.N_273\
        );

    \I__1729\ : InMux
    port map (
            O => \N__8217\,
            I => \N__8208\
        );

    \I__1728\ : InMux
    port map (
            O => \N__8216\,
            I => \N__8208\
        );

    \I__1727\ : InMux
    port map (
            O => \N__8215\,
            I => \N__8203\
        );

    \I__1726\ : InMux
    port map (
            O => \N__8214\,
            I => \N__8203\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__8213\,
            I => \N__8199\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__8208\,
            I => \N__8181\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__8203\,
            I => \N__8181\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8202\,
            I => \N__8176\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8199\,
            I => \N__8176\
        );

    \I__1720\ : InMux
    port map (
            O => \N__8198\,
            I => \N__8173\
        );

    \I__1719\ : InMux
    port map (
            O => \N__8197\,
            I => \N__8168\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8196\,
            I => \N__8168\
        );

    \I__1717\ : InMux
    port map (
            O => \N__8195\,
            I => \N__8165\
        );

    \I__1716\ : InMux
    port map (
            O => \N__8194\,
            I => \N__8162\
        );

    \I__1715\ : InMux
    port map (
            O => \N__8193\,
            I => \N__8156\
        );

    \I__1714\ : InMux
    port map (
            O => \N__8192\,
            I => \N__8156\
        );

    \I__1713\ : InMux
    port map (
            O => \N__8191\,
            I => \N__8153\
        );

    \I__1712\ : InMux
    port map (
            O => \N__8190\,
            I => \N__8148\
        );

    \I__1711\ : InMux
    port map (
            O => \N__8189\,
            I => \N__8148\
        );

    \I__1710\ : InMux
    port map (
            O => \N__8188\,
            I => \N__8141\
        );

    \I__1709\ : InMux
    port map (
            O => \N__8187\,
            I => \N__8141\
        );

    \I__1708\ : InMux
    port map (
            O => \N__8186\,
            I => \N__8141\
        );

    \I__1707\ : Span4Mux_v
    port map (
            O => \N__8181\,
            I => \N__8132\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__8176\,
            I => \N__8132\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__8173\,
            I => \N__8132\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__8168\,
            I => \N__8132\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__8165\,
            I => \N__8122\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__8162\,
            I => \N__8119\
        );

    \I__1701\ : InMux
    port map (
            O => \N__8161\,
            I => \N__8116\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8156\,
            I => \N__8104\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__8153\,
            I => \N__8104\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__8148\,
            I => \N__8104\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__8141\,
            I => \N__8104\
        );

    \I__1696\ : Span4Mux_v
    port map (
            O => \N__8132\,
            I => \N__8104\
        );

    \I__1695\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8101\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8130\,
            I => \N__8096\
        );

    \I__1693\ : InMux
    port map (
            O => \N__8129\,
            I => \N__8096\
        );

    \I__1692\ : InMux
    port map (
            O => \N__8128\,
            I => \N__8092\
        );

    \I__1691\ : InMux
    port map (
            O => \N__8127\,
            I => \N__8085\
        );

    \I__1690\ : InMux
    port map (
            O => \N__8126\,
            I => \N__8085\
        );

    \I__1689\ : InMux
    port map (
            O => \N__8125\,
            I => \N__8085\
        );

    \I__1688\ : Span4Mux_v
    port map (
            O => \N__8122\,
            I => \N__8078\
        );

    \I__1687\ : Span4Mux_v
    port map (
            O => \N__8119\,
            I => \N__8078\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__8116\,
            I => \N__8078\
        );

    \I__1685\ : InMux
    port map (
            O => \N__8115\,
            I => \N__8075\
        );

    \I__1684\ : Span4Mux_v
    port map (
            O => \N__8104\,
            I => \N__8067\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__8101\,
            I => \N__8064\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__8096\,
            I => \N__8061\
        );

    \I__1681\ : InMux
    port map (
            O => \N__8095\,
            I => \N__8058\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__8092\,
            I => \N__8049\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__8085\,
            I => \N__8049\
        );

    \I__1678\ : Span4Mux_h
    port map (
            O => \N__8078\,
            I => \N__8049\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__8075\,
            I => \N__8049\
        );

    \I__1676\ : InMux
    port map (
            O => \N__8074\,
            I => \N__8044\
        );

    \I__1675\ : InMux
    port map (
            O => \N__8073\,
            I => \N__8044\
        );

    \I__1674\ : InMux
    port map (
            O => \N__8072\,
            I => \N__8037\
        );

    \I__1673\ : InMux
    port map (
            O => \N__8071\,
            I => \N__8037\
        );

    \I__1672\ : InMux
    port map (
            O => \N__8070\,
            I => \N__8037\
        );

    \I__1671\ : Span4Mux_h
    port map (
            O => \N__8067\,
            I => \N__8030\
        );

    \I__1670\ : Span4Mux_v
    port map (
            O => \N__8064\,
            I => \N__8030\
        );

    \I__1669\ : Span4Mux_v
    port map (
            O => \N__8061\,
            I => \N__8030\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__8058\,
            I => \N__8021\
        );

    \I__1667\ : Sp12to4
    port map (
            O => \N__8049\,
            I => \N__8021\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__8044\,
            I => \N__8021\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__8037\,
            I => \N__8021\
        );

    \I__1664\ : Span4Mux_h
    port map (
            O => \N__8030\,
            I => \N__8018\
        );

    \I__1663\ : Span12Mux_v
    port map (
            O => \N__8021\,
            I => \N__8015\
        );

    \I__1662\ : Span4Mux_h
    port map (
            O => \N__8018\,
            I => \N__8012\
        );

    \I__1661\ : Span12Mux_h
    port map (
            O => \N__8015\,
            I => \N__8009\
        );

    \I__1660\ : Span4Mux_h
    port map (
            O => \N__8012\,
            I => \N__8006\
        );

    \I__1659\ : Odrv12
    port map (
            O => \N__8009\,
            I => \RESETn_c\
        );

    \I__1658\ : Odrv4
    port map (
            O => \N__8006\,
            I => \RESETn_c\
        );

    \I__1657\ : InMux
    port map (
            O => \N__8001\,
            I => \N__7995\
        );

    \I__1656\ : InMux
    port map (
            O => \N__8000\,
            I => \N__7995\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__7995\,
            I => \N__7992\
        );

    \I__1654\ : Odrv12
    port map (
            O => \N__7992\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1653\ : InMux
    port map (
            O => \N__7989\,
            I => \N__7986\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__7986\,
            I => \N__7983\
        );

    \I__1651\ : Span4Mux_v
    port map (
            O => \N__7983\,
            I => \N__7980\
        );

    \I__1650\ : Sp12to4
    port map (
            O => \N__7980\,
            I => \N__7977\
        );

    \I__1649\ : Span12Mux_h
    port map (
            O => \N__7977\,
            I => \N__7974\
        );

    \I__1648\ : Span12Mux_v
    port map (
            O => \N__7974\,
            I => \N__7971\
        );

    \I__1647\ : Odrv12
    port map (
            O => \N__7971\,
            I => \A_c_19\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__7968\,
            I => \N__7965\
        );

    \I__1645\ : InMux
    port map (
            O => \N__7965\,
            I => \N__7961\
        );

    \I__1644\ : InMux
    port map (
            O => \N__7964\,
            I => \N__7958\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__7961\,
            I => \N__7952\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__7958\,
            I => \N__7952\
        );

    \I__1641\ : CascadeMux
    port map (
            O => \N__7957\,
            I => \N__7949\
        );

    \I__1640\ : Span4Mux_h
    port map (
            O => \N__7952\,
            I => \N__7945\
        );

    \I__1639\ : InMux
    port map (
            O => \N__7949\,
            I => \N__7940\
        );

    \I__1638\ : InMux
    port map (
            O => \N__7948\,
            I => \N__7940\
        );

    \I__1637\ : Odrv4
    port map (
            O => \N__7945\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__7940\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1635\ : IoInMux
    port map (
            O => \N__7935\,
            I => \N__7932\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__7932\,
            I => \N__7929\
        );

    \I__1633\ : IoSpan4Mux
    port map (
            O => \N__7929\,
            I => \N__7926\
        );

    \I__1632\ : IoSpan4Mux
    port map (
            O => \N__7926\,
            I => \N__7923\
        );

    \I__1631\ : Span4Mux_s3_h
    port map (
            O => \N__7923\,
            I => \N__7920\
        );

    \I__1630\ : Sp12to4
    port map (
            O => \N__7920\,
            I => \N__7917\
        );

    \I__1629\ : Odrv12
    port map (
            O => \N__7917\,
            I => \CMA_c_9\
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__7914\,
            I => \N__7911\
        );

    \I__1627\ : InMux
    port map (
            O => \N__7911\,
            I => \N__7908\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__7908\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\
        );

    \I__1625\ : InMux
    port map (
            O => \N__7905\,
            I => \N__7902\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__7902\,
            I => \N__7899\
        );

    \I__1623\ : Sp12to4
    port map (
            O => \N__7899\,
            I => \N__7896\
        );

    \I__1622\ : Span12Mux_v
    port map (
            O => \N__7896\,
            I => \N__7893\
        );

    \I__1621\ : Span12Mux_h
    port map (
            O => \N__7893\,
            I => \N__7890\
        );

    \I__1620\ : Odrv12
    port map (
            O => \N__7890\,
            I => \A_c_16\
        );

    \I__1619\ : InMux
    port map (
            O => \N__7887\,
            I => \N__7884\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__7884\,
            I => \N__7881\
        );

    \I__1617\ : Sp12to4
    port map (
            O => \N__7881\,
            I => \N__7878\
        );

    \I__1616\ : Span12Mux_v
    port map (
            O => \N__7878\,
            I => \N__7875\
        );

    \I__1615\ : Span12Mux_h
    port map (
            O => \N__7875\,
            I => \N__7872\
        );

    \I__1614\ : Odrv12
    port map (
            O => \N__7872\,
            I => \A_c_18\
        );

    \I__1613\ : CascadeMux
    port map (
            O => \N__7869\,
            I => \N__7866\
        );

    \I__1612\ : InMux
    port map (
            O => \N__7866\,
            I => \N__7863\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__7863\,
            I => \N__7860\
        );

    \I__1610\ : Odrv12
    port map (
            O => \N__7860\,
            I => \U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0\
        );

    \I__1609\ : InMux
    port map (
            O => \N__7857\,
            I => \N__7854\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__7854\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1607\ : InMux
    port map (
            O => \N__7851\,
            I => \N__7848\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__7848\,
            I => \N__7845\
        );

    \I__1605\ : Span4Mux_v
    port map (
            O => \N__7845\,
            I => \N__7842\
        );

    \I__1604\ : Sp12to4
    port map (
            O => \N__7842\,
            I => \N__7839\
        );

    \I__1603\ : Span12Mux_h
    port map (
            O => \N__7839\,
            I => \N__7836\
        );

    \I__1602\ : Odrv12
    port map (
            O => \N__7836\,
            I => \A_c_6\
        );

    \I__1601\ : InMux
    port map (
            O => \N__7833\,
            I => \N__7830\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__7830\,
            I => \N__7827\
        );

    \I__1599\ : Span4Mux_v
    port map (
            O => \N__7827\,
            I => \N__7824\
        );

    \I__1598\ : Span4Mux_v
    port map (
            O => \N__7824\,
            I => \N__7821\
        );

    \I__1597\ : Sp12to4
    port map (
            O => \N__7821\,
            I => \N__7818\
        );

    \I__1596\ : Span12Mux_h
    port map (
            O => \N__7818\,
            I => \N__7815\
        );

    \I__1595\ : Odrv12
    port map (
            O => \N__7815\,
            I => \A_c_13\
        );

    \I__1594\ : InMux
    port map (
            O => \N__7812\,
            I => \N__7809\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__7809\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\
        );

    \I__1592\ : InMux
    port map (
            O => \N__7806\,
            I => \N__7803\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__7803\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__1590\ : InMux
    port map (
            O => \N__7800\,
            I => \N__7797\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__7797\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__1588\ : IoInMux
    port map (
            O => \N__7794\,
            I => \N__7791\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__7791\,
            I => \N__7788\
        );

    \I__1586\ : Span12Mux_s4_v
    port map (
            O => \N__7788\,
            I => \N__7785\
        );

    \I__1585\ : Span12Mux_v
    port map (
            O => \N__7785\,
            I => \N__7782\
        );

    \I__1584\ : Odrv12
    port map (
            O => \N__7782\,
            I => \CMA_c_2\
        );

    \I__1583\ : InMux
    port map (
            O => \N__7779\,
            I => \N__7776\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__7776\,
            I => \N__7773\
        );

    \I__1581\ : Span4Mux_v
    port map (
            O => \N__7773\,
            I => \N__7770\
        );

    \I__1580\ : Sp12to4
    port map (
            O => \N__7770\,
            I => \N__7767\
        );

    \I__1579\ : Span12Mux_h
    port map (
            O => \N__7767\,
            I => \N__7764\
        );

    \I__1578\ : Odrv12
    port map (
            O => \N__7764\,
            I => \A_c_5\
        );

    \I__1577\ : InMux
    port map (
            O => \N__7761\,
            I => \N__7758\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__7758\,
            I => \N__7755\
        );

    \I__1575\ : Sp12to4
    port map (
            O => \N__7755\,
            I => \N__7752\
        );

    \I__1574\ : Span12Mux_v
    port map (
            O => \N__7752\,
            I => \N__7749\
        );

    \I__1573\ : Span12Mux_h
    port map (
            O => \N__7749\,
            I => \N__7746\
        );

    \I__1572\ : Odrv12
    port map (
            O => \N__7746\,
            I => \A_c_12\
        );

    \I__1571\ : InMux
    port map (
            O => \N__7743\,
            I => \N__7740\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__7740\,
            I => \U712_BYTE_ENABLE.N_314\
        );

    \I__1569\ : CascadeMux
    port map (
            O => \N__7737\,
            I => \N__7734\
        );

    \I__1568\ : InMux
    port map (
            O => \N__7734\,
            I => \N__7731\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__7731\,
            I => \N__7728\
        );

    \I__1566\ : Span4Mux_v
    port map (
            O => \N__7728\,
            I => \N__7725\
        );

    \I__1565\ : Odrv4
    port map (
            O => \N__7725\,
            I => \U712_BYTE_ENABLE.UUBE\
        );

    \I__1564\ : IoInMux
    port map (
            O => \N__7722\,
            I => \N__7719\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__7719\,
            I => \N__7716\
        );

    \I__1562\ : Odrv12
    port map (
            O => \N__7716\,
            I => \RESETn_c_i\
        );

    \I__1561\ : IoInMux
    port map (
            O => \N__7713\,
            I => \N__7710\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__7710\,
            I => \N__7707\
        );

    \I__1559\ : Span12Mux_s3_h
    port map (
            O => \N__7707\,
            I => \N__7704\
        );

    \I__1558\ : Span12Mux_h
    port map (
            O => \N__7704\,
            I => \N__7701\
        );

    \I__1557\ : Odrv12
    port map (
            O => \N__7701\,
            I => \WEn_c\
        );

    \I__1556\ : IoInMux
    port map (
            O => \N__7698\,
            I => \N__7695\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__7695\,
            I => \N__7692\
        );

    \I__1554\ : Span4Mux_s2_v
    port map (
            O => \N__7692\,
            I => \N__7689\
        );

    \I__1553\ : Span4Mux_v
    port map (
            O => \N__7689\,
            I => \N__7686\
        );

    \I__1552\ : Sp12to4
    port map (
            O => \N__7686\,
            I => \N__7683\
        );

    \I__1551\ : Span12Mux_h
    port map (
            O => \N__7683\,
            I => \N__7680\
        );

    \I__1550\ : Odrv12
    port map (
            O => \N__7680\,
            I => \RASn_c\
        );

    \I__1549\ : InMux
    port map (
            O => \N__7677\,
            I => \N__7673\
        );

    \I__1548\ : InMux
    port map (
            O => \N__7676\,
            I => \N__7670\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__7673\,
            I => \N__7667\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__7670\,
            I => \N__7664\
        );

    \I__1545\ : Span4Mux_h
    port map (
            O => \N__7667\,
            I => \N__7658\
        );

    \I__1544\ : Span4Mux_h
    port map (
            O => \N__7664\,
            I => \N__7655\
        );

    \I__1543\ : InMux
    port map (
            O => \N__7663\,
            I => \N__7652\
        );

    \I__1542\ : CascadeMux
    port map (
            O => \N__7662\,
            I => \N__7648\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7661\,
            I => \N__7644\
        );

    \I__1540\ : Span4Mux_v
    port map (
            O => \N__7658\,
            I => \N__7641\
        );

    \I__1539\ : Span4Mux_v
    port map (
            O => \N__7655\,
            I => \N__7638\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7652\,
            I => \N__7635\
        );

    \I__1537\ : InMux
    port map (
            O => \N__7651\,
            I => \N__7630\
        );

    \I__1536\ : InMux
    port map (
            O => \N__7648\,
            I => \N__7630\
        );

    \I__1535\ : InMux
    port map (
            O => \N__7647\,
            I => \N__7627\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__7644\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__7641\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1532\ : Odrv4
    port map (
            O => \N__7638\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1531\ : Odrv4
    port map (
            O => \N__7635\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__7630\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__7627\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7614\,
            I => \N__7609\
        );

    \I__1527\ : InMux
    port map (
            O => \N__7613\,
            I => \N__7606\
        );

    \I__1526\ : InMux
    port map (
            O => \N__7612\,
            I => \N__7603\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__7609\,
            I => \N__7598\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__7606\,
            I => \N__7598\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__7603\,
            I => \N__7595\
        );

    \I__1522\ : Span4Mux_v
    port map (
            O => \N__7598\,
            I => \N__7588\
        );

    \I__1521\ : Span4Mux_h
    port map (
            O => \N__7595\,
            I => \N__7585\
        );

    \I__1520\ : InMux
    port map (
            O => \N__7594\,
            I => \N__7578\
        );

    \I__1519\ : InMux
    port map (
            O => \N__7593\,
            I => \N__7578\
        );

    \I__1518\ : InMux
    port map (
            O => \N__7592\,
            I => \N__7578\
        );

    \I__1517\ : InMux
    port map (
            O => \N__7591\,
            I => \N__7575\
        );

    \I__1516\ : Odrv4
    port map (
            O => \N__7588\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1515\ : Odrv4
    port map (
            O => \N__7585\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__7578\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__7575\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1512\ : IoInMux
    port map (
            O => \N__7566\,
            I => \N__7563\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__7563\,
            I => \N__7560\
        );

    \I__1510\ : Span4Mux_s0_v
    port map (
            O => \N__7560\,
            I => \N__7557\
        );

    \I__1509\ : Sp12to4
    port map (
            O => \N__7557\,
            I => \N__7554\
        );

    \I__1508\ : Span12Mux_h
    port map (
            O => \N__7554\,
            I => \N__7551\
        );

    \I__1507\ : Span12Mux_v
    port map (
            O => \N__7551\,
            I => \N__7548\
        );

    \I__1506\ : Odrv12
    port map (
            O => \N__7548\,
            I => \CMA_c_10\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7545\,
            I => \N__7542\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__7542\,
            I => \N__7539\
        );

    \I__1503\ : Span4Mux_v
    port map (
            O => \N__7539\,
            I => \N__7536\
        );

    \I__1502\ : Span4Mux_v
    port map (
            O => \N__7536\,
            I => \N__7533\
        );

    \I__1501\ : Sp12to4
    port map (
            O => \N__7533\,
            I => \N__7530\
        );

    \I__1500\ : Span12Mux_h
    port map (
            O => \N__7530\,
            I => \N__7527\
        );

    \I__1499\ : Odrv12
    port map (
            O => \N__7527\,
            I => \A_c_17\
        );

    \I__1498\ : IoInMux
    port map (
            O => \N__7524\,
            I => \N__7521\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__7521\,
            I => \N__7518\
        );

    \I__1496\ : IoSpan4Mux
    port map (
            O => \N__7518\,
            I => \N__7515\
        );

    \I__1495\ : Span4Mux_s1_h
    port map (
            O => \N__7515\,
            I => \N__7512\
        );

    \I__1494\ : Sp12to4
    port map (
            O => \N__7512\,
            I => \N__7509\
        );

    \I__1493\ : Span12Mux_h
    port map (
            O => \N__7509\,
            I => \N__7506\
        );

    \I__1492\ : Odrv12
    port map (
            O => \N__7506\,
            I => \CMA_c_8\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7503\,
            I => \N__7500\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__7500\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__1489\ : CascadeMux
    port map (
            O => \N__7497\,
            I => \U712_REG_SM.N_235_cascade_\
        );

    \I__1488\ : SRMux
    port map (
            O => \N__7494\,
            I => \N__7491\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__7491\,
            I => \N__7488\
        );

    \I__1486\ : Span4Mux_h
    port map (
            O => \N__7488\,
            I => \N__7485\
        );

    \I__1485\ : Odrv4
    port map (
            O => \N__7485\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7482\,
            I => \N__7479\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7479\,
            I => \U712_REG_SM.N_281\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7476\,
            I => \N__7473\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__7473\,
            I => \U712_REG_SM.N_235\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7470\,
            I => \N__7467\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7467\,
            I => \N__7463\
        );

    \I__1478\ : InMux
    port map (
            O => \N__7466\,
            I => \N__7460\
        );

    \I__1477\ : Odrv4
    port map (
            O => \N__7463\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__7460\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7455\,
            I => \N__7452\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7452\,
            I => \N__7446\
        );

    \I__1473\ : InMux
    port map (
            O => \N__7451\,
            I => \N__7443\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7450\,
            I => \N__7440\
        );

    \I__1471\ : InMux
    port map (
            O => \N__7449\,
            I => \N__7437\
        );

    \I__1470\ : Odrv12
    port map (
            O => \N__7446\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__7443\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__7440\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__7437\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1466\ : CascadeMux
    port map (
            O => \N__7428\,
            I => \N__7425\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7425\,
            I => \N__7422\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__7422\,
            I => \N__7419\
        );

    \I__1463\ : Odrv12
    port map (
            O => \N__7419\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\
        );

    \I__1462\ : InMux
    port map (
            O => \N__7416\,
            I => \N__7412\
        );

    \I__1461\ : CascadeMux
    port map (
            O => \N__7415\,
            I => \N__7409\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__7412\,
            I => \N__7405\
        );

    \I__1459\ : InMux
    port map (
            O => \N__7409\,
            I => \N__7402\
        );

    \I__1458\ : InMux
    port map (
            O => \N__7408\,
            I => \N__7399\
        );

    \I__1457\ : Span4Mux_h
    port map (
            O => \N__7405\,
            I => \N__7396\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__7402\,
            I => \N__7393\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__7399\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1454\ : Odrv4
    port map (
            O => \N__7396\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1453\ : Odrv4
    port map (
            O => \N__7393\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1452\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7382\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7385\,
            I => \N__7379\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__7382\,
            I => \N__7374\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__7379\,
            I => \N__7371\
        );

    \I__1448\ : InMux
    port map (
            O => \N__7378\,
            I => \N__7366\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7377\,
            I => \N__7366\
        );

    \I__1446\ : Span12Mux_v
    port map (
            O => \N__7374\,
            I => \N__7363\
        );

    \I__1445\ : Span4Mux_v
    port map (
            O => \N__7371\,
            I => \N__7360\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__7366\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1443\ : Odrv12
    port map (
            O => \N__7363\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__7360\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1441\ : InMux
    port map (
            O => \N__7353\,
            I => \N__7349\
        );

    \I__1440\ : InMux
    port map (
            O => \N__7352\,
            I => \N__7345\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__7349\,
            I => \N__7342\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7348\,
            I => \N__7339\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__7345\,
            I => \U712_REG_SM.N_212\
        );

    \I__1436\ : Odrv12
    port map (
            O => \N__7342\,
            I => \U712_REG_SM.N_212\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__7339\,
            I => \U712_REG_SM.N_212\
        );

    \I__1434\ : InMux
    port map (
            O => \N__7332\,
            I => \N__7329\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__7329\,
            I => \U712_REG_SM.REG_TACK_RNOZ0Z_0\
        );

    \I__1432\ : CascadeMux
    port map (
            O => \N__7326\,
            I => \N__7323\
        );

    \I__1431\ : InMux
    port map (
            O => \N__7323\,
            I => \N__7318\
        );

    \I__1430\ : InMux
    port map (
            O => \N__7322\,
            I => \N__7313\
        );

    \I__1429\ : InMux
    port map (
            O => \N__7321\,
            I => \N__7313\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__7318\,
            I => \REG_TACK\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__7313\,
            I => \REG_TACK\
        );

    \I__1426\ : IoInMux
    port map (
            O => \N__7308\,
            I => \N__7305\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__7305\,
            I => \N__7302\
        );

    \I__1424\ : IoSpan4Mux
    port map (
            O => \N__7302\,
            I => \N__7299\
        );

    \I__1423\ : Span4Mux_s3_h
    port map (
            O => \N__7299\,
            I => \N__7296\
        );

    \I__1422\ : Span4Mux_v
    port map (
            O => \N__7296\,
            I => \N__7293\
        );

    \I__1421\ : Span4Mux_v
    port map (
            O => \N__7293\,
            I => \N__7289\
        );

    \I__1420\ : InMux
    port map (
            O => \N__7292\,
            I => \N__7286\
        );

    \I__1419\ : Sp12to4
    port map (
            O => \N__7289\,
            I => \N__7283\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__7286\,
            I => \N__7280\
        );

    \I__1417\ : Span12Mux_h
    port map (
            O => \N__7283\,
            I => \N__7275\
        );

    \I__1416\ : Span12Mux_v
    port map (
            O => \N__7280\,
            I => \N__7275\
        );

    \I__1415\ : Span12Mux_h
    port map (
            O => \N__7275\,
            I => \N__7272\
        );

    \I__1414\ : Odrv12
    port map (
            O => \N__7272\,
            I => \C3_c\
        );

    \I__1413\ : InMux
    port map (
            O => \N__7269\,
            I => \N__7266\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__7266\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7263\,
            I => \N__7260\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__7260\,
            I => \N__7256\
        );

    \I__1409\ : InMux
    port map (
            O => \N__7259\,
            I => \N__7253\
        );

    \I__1408\ : Span4Mux_v
    port map (
            O => \N__7256\,
            I => \N__7250\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__7253\,
            I => \N__7247\
        );

    \I__1406\ : Odrv4
    port map (
            O => \N__7250\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0Z0Z_0\
        );

    \I__1405\ : Odrv4
    port map (
            O => \N__7247\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0Z0Z_0\
        );

    \I__1404\ : CascadeMux
    port map (
            O => \N__7242\,
            I => \U712_BYTE_ENABLE.N_220_cascade_\
        );

    \I__1403\ : IoInMux
    port map (
            O => \N__7239\,
            I => \N__7236\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__7236\,
            I => \N__7233\
        );

    \I__1401\ : IoSpan4Mux
    port map (
            O => \N__7233\,
            I => \N__7230\
        );

    \I__1400\ : IoSpan4Mux
    port map (
            O => \N__7230\,
            I => \N__7227\
        );

    \I__1399\ : Span4Mux_s3_h
    port map (
            O => \N__7227\,
            I => \N__7224\
        );

    \I__1398\ : Sp12to4
    port map (
            O => \N__7224\,
            I => \N__7221\
        );

    \I__1397\ : Span12Mux_h
    port map (
            O => \N__7221\,
            I => \N__7218\
        );

    \I__1396\ : Span12Mux_v
    port map (
            O => \N__7218\,
            I => \N__7215\
        );

    \I__1395\ : Odrv12
    port map (
            O => \N__7215\,
            I => \N_151_i\
        );

    \I__1394\ : InMux
    port map (
            O => \N__7212\,
            I => \N__7209\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__7209\,
            I => \N__7205\
        );

    \I__1392\ : InMux
    port map (
            O => \N__7208\,
            I => \N__7201\
        );

    \I__1391\ : Span4Mux_h
    port map (
            O => \N__7205\,
            I => \N__7198\
        );

    \I__1390\ : InMux
    port map (
            O => \N__7204\,
            I => \N__7195\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__7201\,
            I => \N__7192\
        );

    \I__1388\ : Odrv4
    port map (
            O => \N__7198\,
            I => \U712_CHIP_RAM.N_386\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__7195\,
            I => \U712_CHIP_RAM.N_386\
        );

    \I__1386\ : Odrv4
    port map (
            O => \N__7192\,
            I => \U712_CHIP_RAM.N_386\
        );

    \I__1385\ : CascadeMux
    port map (
            O => \N__7185\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNO_0Z0Z_3_cascade_\
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__7182\,
            I => \N__7176\
        );

    \I__1383\ : InMux
    port map (
            O => \N__7181\,
            I => \N__7170\
        );

    \I__1382\ : InMux
    port map (
            O => \N__7180\,
            I => \N__7167\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7179\,
            I => \N__7164\
        );

    \I__1380\ : InMux
    port map (
            O => \N__7176\,
            I => \N__7159\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7175\,
            I => \N__7159\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7174\,
            I => \N__7149\
        );

    \I__1377\ : CascadeMux
    port map (
            O => \N__7173\,
            I => \N__7146\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__7170\,
            I => \N__7139\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__7167\,
            I => \N__7139\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__7164\,
            I => \N__7134\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__7159\,
            I => \N__7134\
        );

    \I__1372\ : InMux
    port map (
            O => \N__7158\,
            I => \N__7130\
        );

    \I__1371\ : InMux
    port map (
            O => \N__7157\,
            I => \N__7125\
        );

    \I__1370\ : InMux
    port map (
            O => \N__7156\,
            I => \N__7125\
        );

    \I__1369\ : InMux
    port map (
            O => \N__7155\,
            I => \N__7122\
        );

    \I__1368\ : InMux
    port map (
            O => \N__7154\,
            I => \N__7119\
        );

    \I__1367\ : InMux
    port map (
            O => \N__7153\,
            I => \N__7114\
        );

    \I__1366\ : InMux
    port map (
            O => \N__7152\,
            I => \N__7114\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__7149\,
            I => \N__7111\
        );

    \I__1364\ : InMux
    port map (
            O => \N__7146\,
            I => \N__7108\
        );

    \I__1363\ : InMux
    port map (
            O => \N__7145\,
            I => \N__7105\
        );

    \I__1362\ : InMux
    port map (
            O => \N__7144\,
            I => \N__7102\
        );

    \I__1361\ : Span4Mux_v
    port map (
            O => \N__7139\,
            I => \N__7097\
        );

    \I__1360\ : Span4Mux_v
    port map (
            O => \N__7134\,
            I => \N__7097\
        );

    \I__1359\ : InMux
    port map (
            O => \N__7133\,
            I => \N__7094\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__7130\,
            I => \N__7091\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7125\,
            I => \N__7088\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__7122\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__7119\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__7114\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1353\ : Odrv4
    port map (
            O => \N__7111\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__7108\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__7105\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__7102\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1349\ : Odrv4
    port map (
            O => \N__7097\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__7094\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1347\ : Odrv4
    port map (
            O => \N__7091\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1346\ : Odrv4
    port map (
            O => \N__7088\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__7065\,
            I => \N__7061\
        );

    \I__1344\ : CascadeMux
    port map (
            O => \N__7064\,
            I => \N__7055\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7061\,
            I => \N__7052\
        );

    \I__1342\ : InMux
    port map (
            O => \N__7060\,
            I => \N__7046\
        );

    \I__1341\ : InMux
    port map (
            O => \N__7059\,
            I => \N__7040\
        );

    \I__1340\ : InMux
    port map (
            O => \N__7058\,
            I => \N__7034\
        );

    \I__1339\ : InMux
    port map (
            O => \N__7055\,
            I => \N__7034\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__7052\,
            I => \N__7031\
        );

    \I__1337\ : InMux
    port map (
            O => \N__7051\,
            I => \N__7026\
        );

    \I__1336\ : InMux
    port map (
            O => \N__7050\,
            I => \N__7026\
        );

    \I__1335\ : InMux
    port map (
            O => \N__7049\,
            I => \N__7015\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__7046\,
            I => \N__7012\
        );

    \I__1333\ : InMux
    port map (
            O => \N__7045\,
            I => \N__7009\
        );

    \I__1332\ : InMux
    port map (
            O => \N__7044\,
            I => \N__7004\
        );

    \I__1331\ : InMux
    port map (
            O => \N__7043\,
            I => \N__7004\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__7040\,
            I => \N__7001\
        );

    \I__1329\ : InMux
    port map (
            O => \N__7039\,
            I => \N__6998\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__7034\,
            I => \N__6995\
        );

    \I__1327\ : Span4Mux_v
    port map (
            O => \N__7031\,
            I => \N__6990\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__7026\,
            I => \N__6990\
        );

    \I__1325\ : InMux
    port map (
            O => \N__7025\,
            I => \N__6985\
        );

    \I__1324\ : InMux
    port map (
            O => \N__7024\,
            I => \N__6985\
        );

    \I__1323\ : InMux
    port map (
            O => \N__7023\,
            I => \N__6976\
        );

    \I__1322\ : InMux
    port map (
            O => \N__7022\,
            I => \N__6976\
        );

    \I__1321\ : InMux
    port map (
            O => \N__7021\,
            I => \N__6976\
        );

    \I__1320\ : InMux
    port map (
            O => \N__7020\,
            I => \N__6976\
        );

    \I__1319\ : InMux
    port map (
            O => \N__7019\,
            I => \N__6971\
        );

    \I__1318\ : InMux
    port map (
            O => \N__7018\,
            I => \N__6971\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__7015\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1316\ : Odrv4
    port map (
            O => \N__7012\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__7009\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__7004\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1313\ : Odrv4
    port map (
            O => \N__7001\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__6998\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1311\ : Odrv12
    port map (
            O => \N__6995\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1310\ : Odrv4
    port map (
            O => \N__6990\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__6985\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__6976\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__6971\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1306\ : CascadeMux
    port map (
            O => \N__6948\,
            I => \N__6944\
        );

    \I__1305\ : InMux
    port map (
            O => \N__6947\,
            I => \N__6938\
        );

    \I__1304\ : InMux
    port map (
            O => \N__6944\,
            I => \N__6934\
        );

    \I__1303\ : CascadeMux
    port map (
            O => \N__6943\,
            I => \N__6931\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6942\,
            I => \N__6926\
        );

    \I__1301\ : InMux
    port map (
            O => \N__6941\,
            I => \N__6926\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__6938\,
            I => \N__6923\
        );

    \I__1299\ : InMux
    port map (
            O => \N__6937\,
            I => \N__6918\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__6934\,
            I => \N__6915\
        );

    \I__1297\ : InMux
    port map (
            O => \N__6931\,
            I => \N__6912\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__6926\,
            I => \N__6909\
        );

    \I__1295\ : Span4Mux_h
    port map (
            O => \N__6923\,
            I => \N__6906\
        );

    \I__1294\ : InMux
    port map (
            O => \N__6922\,
            I => \N__6901\
        );

    \I__1293\ : InMux
    port map (
            O => \N__6921\,
            I => \N__6901\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__6918\,
            I => \U712_CHIP_RAM.N_338\
        );

    \I__1291\ : Odrv4
    port map (
            O => \N__6915\,
            I => \U712_CHIP_RAM.N_338\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__6912\,
            I => \U712_CHIP_RAM.N_338\
        );

    \I__1289\ : Odrv4
    port map (
            O => \N__6909\,
            I => \U712_CHIP_RAM.N_338\
        );

    \I__1288\ : Odrv4
    port map (
            O => \N__6906\,
            I => \U712_CHIP_RAM.N_338\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__6901\,
            I => \U712_CHIP_RAM.N_338\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6888\,
            I => \N__6884\
        );

    \I__1285\ : InMux
    port map (
            O => \N__6887\,
            I => \N__6881\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__6884\,
            I => \N__6876\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__6881\,
            I => \N__6876\
        );

    \I__1282\ : Span4Mux_h
    port map (
            O => \N__6876\,
            I => \N__6873\
        );

    \I__1281\ : Odrv4
    port map (
            O => \N__6873\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_1_2\
        );

    \I__1280\ : InMux
    port map (
            O => \N__6870\,
            I => \N__6865\
        );

    \I__1279\ : InMux
    port map (
            O => \N__6869\,
            I => \N__6862\
        );

    \I__1278\ : InMux
    port map (
            O => \N__6868\,
            I => \N__6859\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6865\,
            I => \N__6856\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__6862\,
            I => \N__6850\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__6859\,
            I => \N__6850\
        );

    \I__1274\ : Span4Mux_h
    port map (
            O => \N__6856\,
            I => \N__6847\
        );

    \I__1273\ : InMux
    port map (
            O => \N__6855\,
            I => \N__6844\
        );

    \I__1272\ : Span4Mux_h
    port map (
            O => \N__6850\,
            I => \N__6841\
        );

    \I__1271\ : Odrv4
    port map (
            O => \N__6847\,
            I => \U712_CHIP_RAM.N_342\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__6844\,
            I => \U712_CHIP_RAM.N_342\
        );

    \I__1269\ : Odrv4
    port map (
            O => \N__6841\,
            I => \U712_CHIP_RAM.N_342\
        );

    \I__1268\ : CascadeMux
    port map (
            O => \N__6834\,
            I => \U712_CHIP_RAM.N_293_cascade_\
        );

    \I__1267\ : InMux
    port map (
            O => \N__6831\,
            I => \N__6828\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__6828\,
            I => \U712_CHIP_RAM.N_294\
        );

    \I__1265\ : CascadeMux
    port map (
            O => \N__6825\,
            I => \N__6820\
        );

    \I__1264\ : InMux
    port map (
            O => \N__6824\,
            I => \N__6817\
        );

    \I__1263\ : InMux
    port map (
            O => \N__6823\,
            I => \N__6814\
        );

    \I__1262\ : InMux
    port map (
            O => \N__6820\,
            I => \N__6811\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__6817\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__6814\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__6811\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__1258\ : InMux
    port map (
            O => \N__6804\,
            I => \N__6801\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__6801\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_3\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6798\,
            I => \N__6795\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__6795\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_2\
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__6792\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\
        );

    \I__1253\ : CascadeMux
    port map (
            O => \N__6789\,
            I => \N__6783\
        );

    \I__1252\ : InMux
    port map (
            O => \N__6788\,
            I => \N__6779\
        );

    \I__1251\ : InMux
    port map (
            O => \N__6787\,
            I => \N__6776\
        );

    \I__1250\ : InMux
    port map (
            O => \N__6786\,
            I => \N__6773\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6783\,
            I => \N__6768\
        );

    \I__1248\ : InMux
    port map (
            O => \N__6782\,
            I => \N__6768\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__6779\,
            I => \N__6763\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__6776\,
            I => \N__6763\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__6773\,
            I => \N__6760\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__6768\,
            I => \N__6757\
        );

    \I__1243\ : Span4Mux_v
    port map (
            O => \N__6763\,
            I => \N__6752\
        );

    \I__1242\ : Span4Mux_h
    port map (
            O => \N__6760\,
            I => \N__6752\
        );

    \I__1241\ : Span4Mux_v
    port map (
            O => \N__6757\,
            I => \N__6749\
        );

    \I__1240\ : Odrv4
    port map (
            O => \N__6752\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1239\ : Odrv4
    port map (
            O => \N__6749\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1238\ : InMux
    port map (
            O => \N__6744\,
            I => \N__6741\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__6741\,
            I => \N__6738\
        );

    \I__1236\ : Odrv4
    port map (
            O => \N__6738\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_1_0\
        );

    \I__1235\ : InMux
    port map (
            O => \N__6735\,
            I => \N__6725\
        );

    \I__1234\ : InMux
    port map (
            O => \N__6734\,
            I => \N__6725\
        );

    \I__1233\ : InMux
    port map (
            O => \N__6733\,
            I => \N__6719\
        );

    \I__1232\ : InMux
    port map (
            O => \N__6732\,
            I => \N__6719\
        );

    \I__1231\ : InMux
    port map (
            O => \N__6731\,
            I => \N__6714\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6730\,
            I => \N__6714\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__6725\,
            I => \N__6711\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6724\,
            I => \N__6708\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__6719\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__6714\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1225\ : Odrv4
    port map (
            O => \N__6711\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__6708\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1223\ : InMux
    port map (
            O => \N__6699\,
            I => \N__6694\
        );

    \I__1222\ : InMux
    port map (
            O => \N__6698\,
            I => \N__6691\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6697\,
            I => \N__6688\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6694\,
            I => \U712_CHIP_RAM.N_207\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__6691\,
            I => \U712_CHIP_RAM.N_207\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__6688\,
            I => \U712_CHIP_RAM.N_207\
        );

    \I__1217\ : InMux
    port map (
            O => \N__6681\,
            I => \N__6676\
        );

    \I__1216\ : CascadeMux
    port map (
            O => \N__6680\,
            I => \N__6670\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6679\,
            I => \N__6667\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__6676\,
            I => \N__6663\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6655\
        );

    \I__1212\ : InMux
    port map (
            O => \N__6674\,
            I => \N__6652\
        );

    \I__1211\ : InMux
    port map (
            O => \N__6673\,
            I => \N__6649\
        );

    \I__1210\ : InMux
    port map (
            O => \N__6670\,
            I => \N__6646\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__6667\,
            I => \N__6643\
        );

    \I__1208\ : InMux
    port map (
            O => \N__6666\,
            I => \N__6640\
        );

    \I__1207\ : Span4Mux_h
    port map (
            O => \N__6663\,
            I => \N__6637\
        );

    \I__1206\ : InMux
    port map (
            O => \N__6662\,
            I => \N__6634\
        );

    \I__1205\ : InMux
    port map (
            O => \N__6661\,
            I => \N__6629\
        );

    \I__1204\ : InMux
    port map (
            O => \N__6660\,
            I => \N__6629\
        );

    \I__1203\ : InMux
    port map (
            O => \N__6659\,
            I => \N__6624\
        );

    \I__1202\ : InMux
    port map (
            O => \N__6658\,
            I => \N__6624\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__6655\,
            I => \N__6615\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__6652\,
            I => \N__6615\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__6649\,
            I => \N__6615\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__6646\,
            I => \N__6615\
        );

    \I__1197\ : Odrv4
    port map (
            O => \N__6643\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__6640\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1195\ : Odrv4
    port map (
            O => \N__6637\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__6634\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__6629\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__6624\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1191\ : Odrv4
    port map (
            O => \N__6615\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1190\ : CascadeMux
    port map (
            O => \N__6600\,
            I => \N__6595\
        );

    \I__1189\ : CascadeMux
    port map (
            O => \N__6599\,
            I => \N__6592\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6598\,
            I => \N__6587\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6595\,
            I => \N__6584\
        );

    \I__1186\ : InMux
    port map (
            O => \N__6592\,
            I => \N__6576\
        );

    \I__1185\ : InMux
    port map (
            O => \N__6591\,
            I => \N__6576\
        );

    \I__1184\ : InMux
    port map (
            O => \N__6590\,
            I => \N__6576\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__6587\,
            I => \N__6572\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__6584\,
            I => \N__6569\
        );

    \I__1181\ : CascadeMux
    port map (
            O => \N__6583\,
            I => \N__6566\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6576\,
            I => \N__6560\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6575\,
            I => \N__6557\
        );

    \I__1178\ : Span4Mux_v
    port map (
            O => \N__6572\,
            I => \N__6552\
        );

    \I__1177\ : Span4Mux_v
    port map (
            O => \N__6569\,
            I => \N__6552\
        );

    \I__1176\ : InMux
    port map (
            O => \N__6566\,
            I => \N__6547\
        );

    \I__1175\ : InMux
    port map (
            O => \N__6565\,
            I => \N__6547\
        );

    \I__1174\ : InMux
    port map (
            O => \N__6564\,
            I => \N__6542\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6563\,
            I => \N__6542\
        );

    \I__1172\ : Span4Mux_h
    port map (
            O => \N__6560\,
            I => \N__6539\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__6557\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1170\ : Odrv4
    port map (
            O => \N__6552\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__6547\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__6542\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1167\ : Odrv4
    port map (
            O => \N__6539\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1166\ : InMux
    port map (
            O => \N__6528\,
            I => \N__6525\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6525\,
            I => \U712_CHIP_RAM.N_262\
        );

    \I__1164\ : CascadeMux
    port map (
            O => \N__6522\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_0_cascade_\
        );

    \I__1163\ : InMux
    port map (
            O => \N__6519\,
            I => \N__6516\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__6516\,
            I => \N__6513\
        );

    \I__1161\ : Odrv4
    port map (
            O => \N__6513\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_0\
        );

    \I__1160\ : CascadeMux
    port map (
            O => \N__6510\,
            I => \N__6507\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6507\,
            I => \N__6504\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__6504\,
            I => \U712_CHIP_RAM.N_237\
        );

    \I__1157\ : CascadeMux
    port map (
            O => \N__6501\,
            I => \N__6497\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__6500\,
            I => \N__6493\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6497\,
            I => \N__6487\
        );

    \I__1154\ : InMux
    port map (
            O => \N__6496\,
            I => \N__6482\
        );

    \I__1153\ : InMux
    port map (
            O => \N__6493\,
            I => \N__6482\
        );

    \I__1152\ : InMux
    port map (
            O => \N__6492\,
            I => \N__6476\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6491\,
            I => \N__6471\
        );

    \I__1150\ : InMux
    port map (
            O => \N__6490\,
            I => \N__6471\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__6487\,
            I => \N__6465\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__6482\,
            I => \N__6465\
        );

    \I__1147\ : InMux
    port map (
            O => \N__6481\,
            I => \N__6460\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6480\,
            I => \N__6457\
        );

    \I__1145\ : InMux
    port map (
            O => \N__6479\,
            I => \N__6454\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__6476\,
            I => \N__6451\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__6471\,
            I => \N__6448\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6470\,
            I => \N__6445\
        );

    \I__1141\ : Span4Mux_h
    port map (
            O => \N__6465\,
            I => \N__6442\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6464\,
            I => \N__6439\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6463\,
            I => \N__6436\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__6460\,
            I => \N__6431\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__6457\,
            I => \N__6431\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6454\,
            I => \N__6428\
        );

    \I__1135\ : Span4Mux_h
    port map (
            O => \N__6451\,
            I => \N__6423\
        );

    \I__1134\ : Span4Mux_v
    port map (
            O => \N__6448\,
            I => \N__6423\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6445\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1132\ : Odrv4
    port map (
            O => \N__6442\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__6439\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__6436\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1129\ : Odrv4
    port map (
            O => \N__6431\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1128\ : Odrv12
    port map (
            O => \N__6428\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1127\ : Odrv4
    port map (
            O => \N__6423\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1126\ : InMux
    port map (
            O => \N__6408\,
            I => \N__6405\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6405\,
            I => \N__6402\
        );

    \I__1124\ : Span4Mux_v
    port map (
            O => \N__6402\,
            I => \N__6399\
        );

    \I__1123\ : Span4Mux_h
    port map (
            O => \N__6399\,
            I => \N__6396\
        );

    \I__1122\ : Span4Mux_h
    port map (
            O => \N__6396\,
            I => \N__6393\
        );

    \I__1121\ : Sp12to4
    port map (
            O => \N__6393\,
            I => \N__6390\
        );

    \I__1120\ : Odrv12
    port map (
            O => \N__6390\,
            I => \A_c_4\
        );

    \I__1119\ : InMux
    port map (
            O => \N__6387\,
            I => \N__6384\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6384\,
            I => \N__6381\
        );

    \I__1117\ : Span12Mux_v
    port map (
            O => \N__6381\,
            I => \N__6378\
        );

    \I__1116\ : Span12Mux_h
    port map (
            O => \N__6378\,
            I => \N__6375\
        );

    \I__1115\ : Odrv12
    port map (
            O => \N__6375\,
            I => \A_c_11\
        );

    \I__1114\ : CascadeMux
    port map (
            O => \N__6372\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\
        );

    \I__1113\ : CascadeMux
    port map (
            O => \N__6369\,
            I => \N__6365\
        );

    \I__1112\ : CascadeMux
    port map (
            O => \N__6368\,
            I => \N__6356\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6365\,
            I => \N__6352\
        );

    \I__1110\ : InMux
    port map (
            O => \N__6364\,
            I => \N__6347\
        );

    \I__1109\ : InMux
    port map (
            O => \N__6363\,
            I => \N__6347\
        );

    \I__1108\ : InMux
    port map (
            O => \N__6362\,
            I => \N__6344\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6361\,
            I => \N__6339\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__6360\,
            I => \N__6336\
        );

    \I__1105\ : InMux
    port map (
            O => \N__6359\,
            I => \N__6333\
        );

    \I__1104\ : InMux
    port map (
            O => \N__6356\,
            I => \N__6328\
        );

    \I__1103\ : InMux
    port map (
            O => \N__6355\,
            I => \N__6325\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__6352\,
            I => \N__6318\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__6347\,
            I => \N__6318\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__6344\,
            I => \N__6318\
        );

    \I__1099\ : InMux
    port map (
            O => \N__6343\,
            I => \N__6315\
        );

    \I__1098\ : InMux
    port map (
            O => \N__6342\,
            I => \N__6312\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__6339\,
            I => \N__6309\
        );

    \I__1096\ : InMux
    port map (
            O => \N__6336\,
            I => \N__6306\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__6333\,
            I => \N__6303\
        );

    \I__1094\ : InMux
    port map (
            O => \N__6332\,
            I => \N__6298\
        );

    \I__1093\ : InMux
    port map (
            O => \N__6331\,
            I => \N__6298\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__6328\,
            I => \N__6295\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__6325\,
            I => \N__6290\
        );

    \I__1090\ : Span4Mux_v
    port map (
            O => \N__6318\,
            I => \N__6290\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__6315\,
            I => \N__6287\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__6312\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1087\ : Odrv4
    port map (
            O => \N__6309\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__6306\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1085\ : Odrv12
    port map (
            O => \N__6303\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__6298\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1083\ : Odrv4
    port map (
            O => \N__6295\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1082\ : Odrv4
    port map (
            O => \N__6290\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1081\ : Odrv12
    port map (
            O => \N__6287\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1080\ : InMux
    port map (
            O => \N__6270\,
            I => \N__6267\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__6267\,
            I => \N__6264\
        );

    \I__1078\ : Span4Mux_v
    port map (
            O => \N__6264\,
            I => \N__6260\
        );

    \I__1077\ : InMux
    port map (
            O => \N__6263\,
            I => \N__6257\
        );

    \I__1076\ : Odrv4
    port map (
            O => \N__6260\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_a2_0\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__6257\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_a2_0\
        );

    \I__1074\ : CascadeMux
    port map (
            O => \N__6252\,
            I => \N__6249\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6249\,
            I => \N__6243\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6248\,
            I => \N__6240\
        );

    \I__1071\ : InMux
    port map (
            O => \N__6247\,
            I => \N__6237\
        );

    \I__1070\ : CascadeMux
    port map (
            O => \N__6246\,
            I => \N__6229\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__6243\,
            I => \N__6226\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__6240\,
            I => \N__6221\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__6237\,
            I => \N__6221\
        );

    \I__1066\ : InMux
    port map (
            O => \N__6236\,
            I => \N__6218\
        );

    \I__1065\ : InMux
    port map (
            O => \N__6235\,
            I => \N__6215\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6234\,
            I => \N__6210\
        );

    \I__1063\ : InMux
    port map (
            O => \N__6233\,
            I => \N__6210\
        );

    \I__1062\ : InMux
    port map (
            O => \N__6232\,
            I => \N__6207\
        );

    \I__1061\ : InMux
    port map (
            O => \N__6229\,
            I => \N__6204\
        );

    \I__1060\ : Span4Mux_h
    port map (
            O => \N__6226\,
            I => \N__6199\
        );

    \I__1059\ : Span4Mux_h
    port map (
            O => \N__6221\,
            I => \N__6199\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__6218\,
            I => \U712_CHIP_RAM.N_335\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__6215\,
            I => \U712_CHIP_RAM.N_335\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__6210\,
            I => \U712_CHIP_RAM.N_335\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__6207\,
            I => \U712_CHIP_RAM.N_335\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__6204\,
            I => \U712_CHIP_RAM.N_335\
        );

    \I__1053\ : Odrv4
    port map (
            O => \N__6199\,
            I => \U712_CHIP_RAM.N_335\
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__6186\,
            I => \N__6182\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6185\,
            I => \N__6179\
        );

    \I__1050\ : InMux
    port map (
            O => \N__6182\,
            I => \N__6176\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__6179\,
            I => \U712_CHIP_RAM.N_261\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__6176\,
            I => \U712_CHIP_RAM.N_261\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6167\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6170\,
            I => \N__6163\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__6167\,
            I => \N__6156\
        );

    \I__1044\ : InMux
    port map (
            O => \N__6166\,
            I => \N__6153\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__6163\,
            I => \N__6149\
        );

    \I__1042\ : InMux
    port map (
            O => \N__6162\,
            I => \N__6146\
        );

    \I__1041\ : CascadeMux
    port map (
            O => \N__6161\,
            I => \N__6137\
        );

    \I__1040\ : InMux
    port map (
            O => \N__6160\,
            I => \N__6131\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6159\,
            I => \N__6128\
        );

    \I__1038\ : Span4Mux_v
    port map (
            O => \N__6156\,
            I => \N__6123\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__6153\,
            I => \N__6123\
        );

    \I__1036\ : InMux
    port map (
            O => \N__6152\,
            I => \N__6120\
        );

    \I__1035\ : Span4Mux_h
    port map (
            O => \N__6149\,
            I => \N__6115\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__6146\,
            I => \N__6115\
        );

    \I__1033\ : InMux
    port map (
            O => \N__6145\,
            I => \N__6110\
        );

    \I__1032\ : InMux
    port map (
            O => \N__6144\,
            I => \N__6110\
        );

    \I__1031\ : InMux
    port map (
            O => \N__6143\,
            I => \N__6103\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6142\,
            I => \N__6103\
        );

    \I__1029\ : InMux
    port map (
            O => \N__6141\,
            I => \N__6103\
        );

    \I__1028\ : InMux
    port map (
            O => \N__6140\,
            I => \N__6098\
        );

    \I__1027\ : InMux
    port map (
            O => \N__6137\,
            I => \N__6098\
        );

    \I__1026\ : InMux
    port map (
            O => \N__6136\,
            I => \N__6095\
        );

    \I__1025\ : InMux
    port map (
            O => \N__6135\,
            I => \N__6090\
        );

    \I__1024\ : InMux
    port map (
            O => \N__6134\,
            I => \N__6090\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__6131\,
            I => \U712_CHIP_RAM.N_180\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__6128\,
            I => \U712_CHIP_RAM.N_180\
        );

    \I__1021\ : Odrv4
    port map (
            O => \N__6123\,
            I => \U712_CHIP_RAM.N_180\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__6120\,
            I => \U712_CHIP_RAM.N_180\
        );

    \I__1019\ : Odrv4
    port map (
            O => \N__6115\,
            I => \U712_CHIP_RAM.N_180\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__6110\,
            I => \U712_CHIP_RAM.N_180\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__6103\,
            I => \U712_CHIP_RAM.N_180\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__6098\,
            I => \U712_CHIP_RAM.N_180\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__6095\,
            I => \U712_CHIP_RAM.N_180\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__6090\,
            I => \U712_CHIP_RAM.N_180\
        );

    \I__1013\ : InMux
    port map (
            O => \N__6069\,
            I => \N__6066\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__6066\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_0\
        );

    \I__1011\ : CascadeMux
    port map (
            O => \N__6063\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_0_cascade_\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6060\,
            I => \N__6057\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__6057\,
            I => \U712_BYTE_ENABLE.N_319\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__6054\,
            I => \N__6048\
        );

    \I__1007\ : InMux
    port map (
            O => \N__6053\,
            I => \N__6042\
        );

    \I__1006\ : InMux
    port map (
            O => \N__6052\,
            I => \N__6042\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6038\
        );

    \I__1004\ : InMux
    port map (
            O => \N__6048\,
            I => \N__6033\
        );

    \I__1003\ : InMux
    port map (
            O => \N__6047\,
            I => \N__6033\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__6042\,
            I => \N__6030\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6041\,
            I => \N__6027\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__6038\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__6033\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__998\ : Odrv4
    port map (
            O => \N__6030\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__6027\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__996\ : InMux
    port map (
            O => \N__6018\,
            I => \N__6015\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__6015\,
            I => \U712_REG_SM.un1_STATE_COUNT_4_i_i_0\
        );

    \I__994\ : InMux
    port map (
            O => \N__6012\,
            I => \N__6009\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__6009\,
            I => \U712_REG_SM.N_26\
        );

    \I__992\ : CascadeMux
    port map (
            O => \N__6006\,
            I => \N__6003\
        );

    \I__991\ : InMux
    port map (
            O => \N__6003\,
            I => \N__6000\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__6000\,
            I => \U712_REG_SM.N_274\
        );

    \I__989\ : IoInMux
    port map (
            O => \N__5997\,
            I => \N__5994\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__5994\,
            I => \N__5991\
        );

    \I__987\ : IoSpan4Mux
    port map (
            O => \N__5991\,
            I => \N__5988\
        );

    \I__986\ : Span4Mux_s2_v
    port map (
            O => \N__5988\,
            I => \N__5985\
        );

    \I__985\ : Span4Mux_v
    port map (
            O => \N__5985\,
            I => \N__5982\
        );

    \I__984\ : Span4Mux_h
    port map (
            O => \N__5982\,
            I => \N__5979\
        );

    \I__983\ : Odrv4
    port map (
            O => \N__5979\,
            I => \DMA_LATCH_EN_c\
        );

    \I__982\ : IoInMux
    port map (
            O => \N__5976\,
            I => \N__5973\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__5973\,
            I => \N__5970\
        );

    \I__980\ : Span12Mux_s6_v
    port map (
            O => \N__5970\,
            I => \N__5967\
        );

    \I__979\ : Odrv12
    port map (
            O => \N__5967\,
            I => \CONSTANT_ONE_NET\
        );

    \I__978\ : InMux
    port map (
            O => \N__5964\,
            I => \N__5961\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__5961\,
            I => \N__5958\
        );

    \I__976\ : Span12Mux_v
    port map (
            O => \N__5958\,
            I => \N__5955\
        );

    \I__975\ : Span12Mux_h
    port map (
            O => \N__5955\,
            I => \N__5952\
        );

    \I__974\ : Odrv12
    port map (
            O => \N__5952\,
            I => \A_c_15\
        );

    \I__973\ : InMux
    port map (
            O => \N__5949\,
            I => \N__5946\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__5946\,
            I => \N__5943\
        );

    \I__971\ : Span4Mux_v
    port map (
            O => \N__5943\,
            I => \N__5940\
        );

    \I__970\ : Sp12to4
    port map (
            O => \N__5940\,
            I => \N__5937\
        );

    \I__969\ : Span12Mux_h
    port map (
            O => \N__5937\,
            I => \N__5934\
        );

    \I__968\ : Odrv12
    port map (
            O => \N__5934\,
            I => \A_c_8\
        );

    \I__967\ : InMux
    port map (
            O => \N__5931\,
            I => \N__5928\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5928\,
            I => \N__5925\
        );

    \I__965\ : Span12Mux_v
    port map (
            O => \N__5925\,
            I => \N__5922\
        );

    \I__964\ : Span12Mux_h
    port map (
            O => \N__5922\,
            I => \N__5919\
        );

    \I__963\ : Odrv12
    port map (
            O => \N__5919\,
            I => \A_c_2\
        );

    \I__962\ : InMux
    port map (
            O => \N__5916\,
            I => \N__5913\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__5913\,
            I => \N__5910\
        );

    \I__960\ : Span12Mux_h
    port map (
            O => \N__5910\,
            I => \N__5907\
        );

    \I__959\ : Odrv12
    port map (
            O => \N__5907\,
            I => \A_c_9\
        );

    \I__958\ : InMux
    port map (
            O => \N__5904\,
            I => \N__5901\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__5901\,
            I => \N__5898\
        );

    \I__956\ : Span4Mux_v
    port map (
            O => \N__5898\,
            I => \N__5895\
        );

    \I__955\ : Odrv4
    port map (
            O => \N__5895\,
            I => \U712_REG_SM.N_383\
        );

    \I__954\ : CascadeMux
    port map (
            O => \N__5892\,
            I => \U712_REG_SM.N_383_cascade_\
        );

    \I__953\ : InMux
    port map (
            O => \N__5889\,
            I => \N__5885\
        );

    \I__952\ : InMux
    port map (
            O => \N__5888\,
            I => \N__5873\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__5885\,
            I => \N__5870\
        );

    \I__950\ : InMux
    port map (
            O => \N__5884\,
            I => \N__5867\
        );

    \I__949\ : InMux
    port map (
            O => \N__5883\,
            I => \N__5864\
        );

    \I__948\ : InMux
    port map (
            O => \N__5882\,
            I => \N__5861\
        );

    \I__947\ : InMux
    port map (
            O => \N__5881\,
            I => \N__5858\
        );

    \I__946\ : InMux
    port map (
            O => \N__5880\,
            I => \N__5853\
        );

    \I__945\ : InMux
    port map (
            O => \N__5879\,
            I => \N__5853\
        );

    \I__944\ : InMux
    port map (
            O => \N__5878\,
            I => \N__5846\
        );

    \I__943\ : InMux
    port map (
            O => \N__5877\,
            I => \N__5846\
        );

    \I__942\ : InMux
    port map (
            O => \N__5876\,
            I => \N__5846\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__5873\,
            I => \N__5843\
        );

    \I__940\ : Odrv4
    port map (
            O => \N__5870\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__5867\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__5864\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__5861\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__5858\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__5853\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5846\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__933\ : Odrv4
    port map (
            O => \N__5843\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__932\ : CascadeMux
    port map (
            O => \N__5826\,
            I => \U712_CYCLE_TERM.N_321_cascade_\
        );

    \I__931\ : CascadeMux
    port map (
            O => \N__5823\,
            I => \N__5820\
        );

    \I__930\ : InMux
    port map (
            O => \N__5820\,
            I => \N__5816\
        );

    \I__929\ : InMux
    port map (
            O => \N__5819\,
            I => \N__5813\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__5816\,
            I => \N__5808\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__5813\,
            I => \N__5808\
        );

    \I__926\ : Odrv12
    port map (
            O => \N__5808\,
            I => \CPU_TACKm\
        );

    \I__925\ : IoInMux
    port map (
            O => \N__5805\,
            I => \N__5802\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__5802\,
            I => \N__5799\
        );

    \I__923\ : IoSpan4Mux
    port map (
            O => \N__5799\,
            I => \N__5796\
        );

    \I__922\ : Sp12to4
    port map (
            O => \N__5796\,
            I => \N__5793\
        );

    \I__921\ : Span12Mux_s7_v
    port map (
            O => \N__5793\,
            I => \N__5790\
        );

    \I__920\ : Span12Mux_v
    port map (
            O => \N__5790\,
            I => \N__5787\
        );

    \I__919\ : Odrv12
    port map (
            O => \N__5787\,
            I => \N_156_i\
        );

    \I__918\ : InMux
    port map (
            O => \N__5784\,
            I => \N__5781\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__5781\,
            I => \N__5777\
        );

    \I__916\ : InMux
    port map (
            O => \N__5780\,
            I => \N__5774\
        );

    \I__915\ : Odrv12
    port map (
            O => \N__5777\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1Z0Z_0\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__5774\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1Z0Z_0\
        );

    \I__913\ : IoInMux
    port map (
            O => \N__5769\,
            I => \N__5766\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__5766\,
            I => \N__5763\
        );

    \I__911\ : Span12Mux_s5_h
    port map (
            O => \N__5763\,
            I => \N__5760\
        );

    \I__910\ : Span12Mux_h
    port map (
            O => \N__5760\,
            I => \N__5757\
        );

    \I__909\ : Span12Mux_v
    port map (
            O => \N__5757\,
            I => \N__5754\
        );

    \I__908\ : Odrv12
    port map (
            O => \N__5754\,
            I => \N_126_i\
        );

    \I__907\ : CascadeMux
    port map (
            O => \N__5751\,
            I => \N__5748\
        );

    \I__906\ : InMux
    port map (
            O => \N__5748\,
            I => \N__5742\
        );

    \I__905\ : InMux
    port map (
            O => \N__5747\,
            I => \N__5742\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__5742\,
            I => \U712_BYTE_ENABLE.N_315\
        );

    \I__903\ : CascadeMux
    port map (
            O => \N__5739\,
            I => \U712_CHIP_RAM.N_184_cascade_\
        );

    \I__902\ : InMux
    port map (
            O => \N__5736\,
            I => \N__5733\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__5733\,
            I => \N__5730\
        );

    \I__900\ : Odrv4
    port map (
            O => \N__5730\,
            I => \U712_CHIP_RAM.N_304\
        );

    \I__899\ : InMux
    port map (
            O => \N__5727\,
            I => \N__5724\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__5724\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERlde_0_0_a2_0\
        );

    \I__897\ : CascadeMux
    port map (
            O => \N__5721\,
            I => \U712_CHIP_RAM.N_392_cascade_\
        );

    \I__896\ : CEMux
    port map (
            O => \N__5718\,
            I => \N__5714\
        );

    \I__895\ : CEMux
    port map (
            O => \N__5717\,
            I => \N__5710\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__5714\,
            I => \N__5707\
        );

    \I__893\ : CEMux
    port map (
            O => \N__5713\,
            I => \N__5704\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__5710\,
            I => \N__5701\
        );

    \I__891\ : Span4Mux_h
    port map (
            O => \N__5707\,
            I => \N__5696\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__5704\,
            I => \N__5696\
        );

    \I__889\ : Sp12to4
    port map (
            O => \N__5701\,
            I => \N__5693\
        );

    \I__888\ : Sp12to4
    port map (
            O => \N__5696\,
            I => \N__5690\
        );

    \I__887\ : Odrv12
    port map (
            O => \N__5693\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__886\ : Odrv12
    port map (
            O => \N__5690\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__885\ : InMux
    port map (
            O => \N__5685\,
            I => \N__5682\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__5682\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_0\
        );

    \I__883\ : CascadeMux
    port map (
            O => \N__5679\,
            I => \N__5676\
        );

    \I__882\ : InMux
    port map (
            O => \N__5676\,
            I => \N__5672\
        );

    \I__881\ : InMux
    port map (
            O => \N__5675\,
            I => \N__5669\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__5672\,
            I => \N__5664\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__5669\,
            I => \N__5664\
        );

    \I__878\ : Odrv4
    port map (
            O => \N__5664\,
            I => \U712_REG_SM.N_196\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__5661\,
            I => \N__5656\
        );

    \I__876\ : InMux
    port map (
            O => \N__5660\,
            I => \N__5653\
        );

    \I__875\ : InMux
    port map (
            O => \N__5659\,
            I => \N__5650\
        );

    \I__874\ : InMux
    port map (
            O => \N__5656\,
            I => \N__5647\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__5653\,
            I => \U712_CHIP_RAM.N_333\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__5650\,
            I => \U712_CHIP_RAM.N_333\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__5647\,
            I => \U712_CHIP_RAM.N_333\
        );

    \I__870\ : CascadeMux
    port map (
            O => \N__5640\,
            I => \U712_CHIP_RAM.N_310_cascade_\
        );

    \I__869\ : CascadeMux
    port map (
            O => \N__5637\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_\
        );

    \I__868\ : CEMux
    port map (
            O => \N__5634\,
            I => \N__5631\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__5631\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0\
        );

    \I__866\ : InMux
    port map (
            O => \N__5628\,
            I => \N__5624\
        );

    \I__865\ : InMux
    port map (
            O => \N__5627\,
            I => \N__5620\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__5624\,
            I => \N__5617\
        );

    \I__863\ : InMux
    port map (
            O => \N__5623\,
            I => \N__5614\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__5620\,
            I => \N__5606\
        );

    \I__861\ : Span4Mux_v
    port map (
            O => \N__5617\,
            I => \N__5606\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__5614\,
            I => \N__5606\
        );

    \I__859\ : InMux
    port map (
            O => \N__5613\,
            I => \N__5603\
        );

    \I__858\ : Span4Mux_h
    port map (
            O => \N__5606\,
            I => \N__5599\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__5603\,
            I => \N__5596\
        );

    \I__856\ : InMux
    port map (
            O => \N__5602\,
            I => \N__5593\
        );

    \I__855\ : Odrv4
    port map (
            O => \N__5599\,
            I => \DMA_CYCLEm\
        );

    \I__854\ : Odrv4
    port map (
            O => \N__5596\,
            I => \DMA_CYCLEm\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5593\,
            I => \DMA_CYCLEm\
        );

    \I__852\ : IoInMux
    port map (
            O => \N__5586\,
            I => \N__5583\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__5583\,
            I => \N__5580\
        );

    \I__850\ : Span4Mux_s3_v
    port map (
            O => \N__5580\,
            I => \N__5575\
        );

    \I__849\ : InMux
    port map (
            O => \N__5579\,
            I => \N__5572\
        );

    \I__848\ : InMux
    port map (
            O => \N__5578\,
            I => \N__5569\
        );

    \I__847\ : Span4Mux_h
    port map (
            O => \N__5575\,
            I => \N__5566\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__5572\,
            I => \N__5563\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__5569\,
            I => \N__5560\
        );

    \I__844\ : Sp12to4
    port map (
            O => \N__5566\,
            I => \N__5556\
        );

    \I__843\ : Span4Mux_v
    port map (
            O => \N__5563\,
            I => \N__5553\
        );

    \I__842\ : Span4Mux_h
    port map (
            O => \N__5560\,
            I => \N__5550\
        );

    \I__841\ : InMux
    port map (
            O => \N__5559\,
            I => \N__5547\
        );

    \I__840\ : Odrv12
    port map (
            O => \N__5556\,
            I => \DBENn_c\
        );

    \I__839\ : Odrv4
    port map (
            O => \N__5553\,
            I => \DBENn_c\
        );

    \I__838\ : Odrv4
    port map (
            O => \N__5550\,
            I => \DBENn_c\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__5547\,
            I => \DBENn_c\
        );

    \I__836\ : InMux
    port map (
            O => \N__5538\,
            I => \N__5535\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__5535\,
            I => \N__5531\
        );

    \I__834\ : InMux
    port map (
            O => \N__5534\,
            I => \N__5528\
        );

    \I__833\ : Odrv4
    port map (
            O => \N__5531\,
            I => \U712_CHIP_RAM.N_334\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__5528\,
            I => \U712_CHIP_RAM.N_334\
        );

    \I__831\ : InMux
    port map (
            O => \N__5523\,
            I => \N__5520\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__5520\,
            I => \U712_CHIP_RAM.N_297\
        );

    \I__829\ : InMux
    port map (
            O => \N__5517\,
            I => \N__5514\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__5514\,
            I => \N__5510\
        );

    \I__827\ : InMux
    port map (
            O => \N__5513\,
            I => \N__5507\
        );

    \I__826\ : Span4Mux_v
    port map (
            O => \N__5510\,
            I => \N__5502\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__5507\,
            I => \N__5502\
        );

    \I__824\ : Odrv4
    port map (
            O => \N__5502\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_0_0\
        );

    \I__823\ : InMux
    port map (
            O => \N__5499\,
            I => \N__5495\
        );

    \I__822\ : InMux
    port map (
            O => \N__5498\,
            I => \N__5492\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5495\,
            I => \U712_CHIP_RAM.N_202\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__5492\,
            I => \U712_CHIP_RAM.N_202\
        );

    \I__819\ : InMux
    port map (
            O => \N__5487\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__818\ : InMux
    port map (
            O => \N__5484\,
            I => \N__5480\
        );

    \I__817\ : InMux
    port map (
            O => \N__5483\,
            I => \N__5477\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__5480\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__5477\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__814\ : ClkMux
    port map (
            O => \N__5472\,
            I => \N__5445\
        );

    \I__813\ : ClkMux
    port map (
            O => \N__5471\,
            I => \N__5445\
        );

    \I__812\ : ClkMux
    port map (
            O => \N__5470\,
            I => \N__5445\
        );

    \I__811\ : ClkMux
    port map (
            O => \N__5469\,
            I => \N__5445\
        );

    \I__810\ : ClkMux
    port map (
            O => \N__5468\,
            I => \N__5445\
        );

    \I__809\ : ClkMux
    port map (
            O => \N__5467\,
            I => \N__5445\
        );

    \I__808\ : ClkMux
    port map (
            O => \N__5466\,
            I => \N__5445\
        );

    \I__807\ : ClkMux
    port map (
            O => \N__5465\,
            I => \N__5445\
        );

    \I__806\ : ClkMux
    port map (
            O => \N__5464\,
            I => \N__5445\
        );

    \I__805\ : GlobalMux
    port map (
            O => \N__5445\,
            I => \N__5442\
        );

    \I__804\ : gio2CtrlBuf
    port map (
            O => \N__5442\,
            I => \C1_c_g\
        );

    \I__803\ : InMux
    port map (
            O => \N__5439\,
            I => \N__5436\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__5436\,
            I => \U712_CHIP_RAM.N_134\
        );

    \I__801\ : InMux
    port map (
            O => \N__5433\,
            I => \N__5430\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__5430\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\
        );

    \I__799\ : IoInMux
    port map (
            O => \N__5427\,
            I => \N__5424\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__5424\,
            I => \N__5421\
        );

    \I__797\ : IoSpan4Mux
    port map (
            O => \N__5421\,
            I => \N__5418\
        );

    \I__796\ : IoSpan4Mux
    port map (
            O => \N__5418\,
            I => \N__5415\
        );

    \I__795\ : Span4Mux_s2_h
    port map (
            O => \N__5415\,
            I => \N__5412\
        );

    \I__794\ : Sp12to4
    port map (
            O => \N__5412\,
            I => \N__5409\
        );

    \I__793\ : Span12Mux_s9_h
    port map (
            O => \N__5409\,
            I => \N__5406\
        );

    \I__792\ : Odrv12
    port map (
            O => \N__5406\,
            I => \N_116_i\
        );

    \I__791\ : CascadeMux
    port map (
            O => \N__5403\,
            I => \U712_CHIP_RAM.N_207_cascade_\
        );

    \I__790\ : CascadeMux
    port map (
            O => \N__5400\,
            I => \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_1_cascade_\
        );

    \I__789\ : CascadeMux
    port map (
            O => \N__5397\,
            I => \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_2_cascade_\
        );

    \I__788\ : CascadeMux
    port map (
            O => \N__5394\,
            I => \U712_REG_SM.N_284_cascade_\
        );

    \I__787\ : InMux
    port map (
            O => \N__5391\,
            I => \N__5387\
        );

    \I__786\ : InMux
    port map (
            O => \N__5390\,
            I => \N__5384\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__5387\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__5384\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__783\ : InMux
    port map (
            O => \N__5379\,
            I => \bfn_10_15_0_\
        );

    \I__782\ : InMux
    port map (
            O => \N__5376\,
            I => \N__5372\
        );

    \I__781\ : InMux
    port map (
            O => \N__5375\,
            I => \N__5369\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__5372\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5369\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__778\ : InMux
    port map (
            O => \N__5364\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__777\ : InMux
    port map (
            O => \N__5361\,
            I => \N__5357\
        );

    \I__776\ : InMux
    port map (
            O => \N__5360\,
            I => \N__5354\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5357\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__5354\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__773\ : InMux
    port map (
            O => \N__5349\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__772\ : InMux
    port map (
            O => \N__5346\,
            I => \N__5342\
        );

    \I__771\ : InMux
    port map (
            O => \N__5345\,
            I => \N__5339\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__5342\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__5339\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__768\ : InMux
    port map (
            O => \N__5334\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__767\ : CascadeMux
    port map (
            O => \N__5331\,
            I => \N__5327\
        );

    \I__766\ : InMux
    port map (
            O => \N__5330\,
            I => \N__5324\
        );

    \I__765\ : InMux
    port map (
            O => \N__5327\,
            I => \N__5321\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5324\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__5321\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__762\ : InMux
    port map (
            O => \N__5316\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__761\ : InMux
    port map (
            O => \N__5313\,
            I => \N__5309\
        );

    \I__760\ : InMux
    port map (
            O => \N__5312\,
            I => \N__5306\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__5309\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5306\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__757\ : InMux
    port map (
            O => \N__5301\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__756\ : InMux
    port map (
            O => \N__5298\,
            I => \N__5294\
        );

    \I__755\ : InMux
    port map (
            O => \N__5297\,
            I => \N__5291\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__5294\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__5291\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__752\ : InMux
    port map (
            O => \N__5286\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__751\ : InMux
    port map (
            O => \N__5283\,
            I => \N__5280\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__5280\,
            I => \N__5277\
        );

    \I__749\ : Odrv4
    port map (
            O => \N__5277\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER18\
        );

    \I__748\ : InMux
    port map (
            O => \N__5274\,
            I => \N__5264\
        );

    \I__747\ : InMux
    port map (
            O => \N__5273\,
            I => \N__5264\
        );

    \I__746\ : InMux
    port map (
            O => \N__5272\,
            I => \N__5264\
        );

    \I__745\ : InMux
    port map (
            O => \N__5271\,
            I => \N__5261\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__5264\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__5261\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__742\ : InMux
    port map (
            O => \N__5256\,
            I => \N__5253\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__5253\,
            I => \U712_REG_SM.STATE_COUNT_srsts_i_0_a2_0_0_0\
        );

    \I__740\ : InMux
    port map (
            O => \N__5250\,
            I => \N__5247\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__5247\,
            I => \U712_REG_SM.N_222\
        );

    \I__738\ : CascadeMux
    port map (
            O => \N__5244\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_\
        );

    \I__737\ : CascadeMux
    port map (
            O => \N__5241\,
            I => \N__5236\
        );

    \I__736\ : InMux
    port map (
            O => \N__5240\,
            I => \N__5231\
        );

    \I__735\ : InMux
    port map (
            O => \N__5239\,
            I => \N__5231\
        );

    \I__734\ : InMux
    port map (
            O => \N__5236\,
            I => \N__5228\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__5231\,
            I => \N__5225\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__5228\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__731\ : Odrv4
    port map (
            O => \N__5225\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__730\ : InMux
    port map (
            O => \N__5220\,
            I => \N__5216\
        );

    \I__729\ : InMux
    port map (
            O => \N__5219\,
            I => \N__5213\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__5216\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__5213\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__726\ : InMux
    port map (
            O => \N__5208\,
            I => \N__5205\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__5205\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__724\ : InMux
    port map (
            O => \N__5202\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__723\ : InMux
    port map (
            O => \N__5199\,
            I => \N__5195\
        );

    \I__722\ : InMux
    port map (
            O => \N__5198\,
            I => \N__5192\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__5195\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__5192\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__719\ : InMux
    port map (
            O => \N__5187\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__718\ : InMux
    port map (
            O => \N__5184\,
            I => \N__5180\
        );

    \I__717\ : InMux
    port map (
            O => \N__5183\,
            I => \N__5177\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__5180\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__5177\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__714\ : InMux
    port map (
            O => \N__5172\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__713\ : CascadeMux
    port map (
            O => \N__5169\,
            I => \N__5166\
        );

    \I__712\ : InMux
    port map (
            O => \N__5166\,
            I => \N__5162\
        );

    \I__711\ : InMux
    port map (
            O => \N__5165\,
            I => \N__5153\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__5162\,
            I => \N__5150\
        );

    \I__709\ : InMux
    port map (
            O => \N__5161\,
            I => \N__5141\
        );

    \I__708\ : InMux
    port map (
            O => \N__5160\,
            I => \N__5141\
        );

    \I__707\ : InMux
    port map (
            O => \N__5159\,
            I => \N__5141\
        );

    \I__706\ : InMux
    port map (
            O => \N__5158\,
            I => \N__5141\
        );

    \I__705\ : InMux
    port map (
            O => \N__5157\,
            I => \N__5136\
        );

    \I__704\ : InMux
    port map (
            O => \N__5156\,
            I => \N__5136\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__5153\,
            I => \N__5133\
        );

    \I__702\ : Odrv4
    port map (
            O => \N__5150\,
            I => \U712_CHIP_RAM.N_46\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__5141\,
            I => \U712_CHIP_RAM.N_46\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__5136\,
            I => \U712_CHIP_RAM.N_46\
        );

    \I__699\ : Odrv4
    port map (
            O => \N__5133\,
            I => \U712_CHIP_RAM.N_46\
        );

    \I__698\ : InMux
    port map (
            O => \N__5124\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__697\ : InMux
    port map (
            O => \N__5121\,
            I => \N__5117\
        );

    \I__696\ : InMux
    port map (
            O => \N__5120\,
            I => \N__5114\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__5117\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__5114\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__693\ : InMux
    port map (
            O => \N__5109\,
            I => \N__5106\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__5106\,
            I => \U712_CYCLE_TERM.N_217_i_0_en\
        );

    \I__691\ : InMux
    port map (
            O => \N__5103\,
            I => \N__5100\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__5100\,
            I => \U712_REG_SM.START_RST_0_sqmuxa\
        );

    \I__689\ : InMux
    port map (
            O => \N__5097\,
            I => \N__5091\
        );

    \I__688\ : InMux
    port map (
            O => \N__5096\,
            I => \N__5091\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__5091\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__686\ : CascadeMux
    port map (
            O => \N__5088\,
            I => \U712_REG_SM.N_285_cascade_\
        );

    \I__685\ : CascadeMux
    port map (
            O => \N__5085\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER18_cascade_\
        );

    \I__684\ : InMux
    port map (
            O => \N__5082\,
            I => \N__5079\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__5079\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_0\
        );

    \I__682\ : InMux
    port map (
            O => \N__5076\,
            I => \N__5073\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__5073\,
            I => \U712_CHIP_RAM.N_239\
        );

    \I__680\ : InMux
    port map (
            O => \N__5070\,
            I => \N__5067\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__5067\,
            I => \U712_CHIP_RAM.N_269\
        );

    \I__678\ : CascadeMux
    port map (
            O => \N__5064\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_0_0_a2_1_1_cascade_\
        );

    \I__677\ : InMux
    port map (
            O => \N__5061\,
            I => \N__5058\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__5058\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__675\ : InMux
    port map (
            O => \N__5055\,
            I => \bfn_10_12_0_\
        );

    \I__674\ : InMux
    port map (
            O => \N__5052\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__673\ : InMux
    port map (
            O => \N__5049\,
            I => \N__5046\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__5046\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__671\ : InMux
    port map (
            O => \N__5043\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__670\ : InMux
    port map (
            O => \N__5040\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__669\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5034\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__5034\,
            I => \N__5031\
        );

    \I__667\ : Span4Mux_v
    port map (
            O => \N__5031\,
            I => \N__5028\
        );

    \I__666\ : Odrv4
    port map (
            O => \N__5028\,
            I => \U712_CHIP_RAM.BANK0_RNOZ0Z_3\
        );

    \I__665\ : CascadeMux
    port map (
            O => \N__5025\,
            I => \N__5021\
        );

    \I__664\ : InMux
    port map (
            O => \N__5024\,
            I => \N__5018\
        );

    \I__663\ : InMux
    port map (
            O => \N__5021\,
            I => \N__5015\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__5018\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__5015\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\
        );

    \I__660\ : InMux
    port map (
            O => \N__5010\,
            I => \N__5006\
        );

    \I__659\ : InMux
    port map (
            O => \N__5009\,
            I => \N__5003\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__5006\,
            I => \N__5000\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__5003\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__656\ : Odrv4
    port map (
            O => \N__5000\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__655\ : InMux
    port map (
            O => \N__4995\,
            I => \N__4992\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__4992\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__653\ : CascadeMux
    port map (
            O => \N__4989\,
            I => \U712_CHIP_RAM.BANK0_RNOZ0Z_1_cascade_\
        );

    \I__652\ : IoInMux
    port map (
            O => \N__4986\,
            I => \N__4983\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__4983\,
            I => \N__4980\
        );

    \I__650\ : Span4Mux_s3_v
    port map (
            O => \N__4980\,
            I => \N__4977\
        );

    \I__649\ : Span4Mux_v
    port map (
            O => \N__4977\,
            I => \N__4974\
        );

    \I__648\ : Span4Mux_v
    port map (
            O => \N__4974\,
            I => \N__4971\
        );

    \I__647\ : Span4Mux_v
    port map (
            O => \N__4971\,
            I => \N__4967\
        );

    \I__646\ : InMux
    port map (
            O => \N__4970\,
            I => \N__4964\
        );

    \I__645\ : Odrv4
    port map (
            O => \N__4967\,
            I => \BANK0_c\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__4964\,
            I => \BANK0_c\
        );

    \I__643\ : InMux
    port map (
            O => \N__4959\,
            I => \N__4956\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__4956\,
            I => \U712_CHIP_RAM.BANK0_RNOZ0Z_4\
        );

    \I__641\ : InMux
    port map (
            O => \N__4953\,
            I => \N__4949\
        );

    \I__640\ : InMux
    port map (
            O => \N__4952\,
            I => \N__4946\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__4949\,
            I => \U712_CHIP_RAM.N_186\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__4946\,
            I => \U712_CHIP_RAM.N_186\
        );

    \I__637\ : CascadeMux
    port map (
            O => \N__4941\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_0_a2_0_0_cascade_\
        );

    \I__636\ : InMux
    port map (
            O => \N__4938\,
            I => \N__4935\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__4935\,
            I => \U712_CHIP_RAM.N_306\
        );

    \I__634\ : CascadeMux
    port map (
            O => \N__4932\,
            I => \U712_CHIP_RAM.N_333_cascade_\
        );

    \I__633\ : CascadeMux
    port map (
            O => \N__4929\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_0_0_a2_1_0_cascade_\
        );

    \I__632\ : InMux
    port map (
            O => \N__4926\,
            I => \N__4922\
        );

    \I__631\ : IoInMux
    port map (
            O => \N__4925\,
            I => \N__4919\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4922\,
            I => \N__4916\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__4919\,
            I => \N__4913\
        );

    \I__628\ : Span4Mux_v
    port map (
            O => \N__4916\,
            I => \N__4910\
        );

    \I__627\ : IoSpan4Mux
    port map (
            O => \N__4913\,
            I => \N__4907\
        );

    \I__626\ : Sp12to4
    port map (
            O => \N__4910\,
            I => \N__4904\
        );

    \I__625\ : IoSpan4Mux
    port map (
            O => \N__4907\,
            I => \N__4901\
        );

    \I__624\ : Span12Mux_h
    port map (
            O => \N__4904\,
            I => \N__4898\
        );

    \I__623\ : IoSpan4Mux
    port map (
            O => \N__4901\,
            I => \N__4895\
        );

    \I__622\ : Odrv12
    port map (
            O => \N__4898\,
            I => \C1_c\
        );

    \I__621\ : Odrv4
    port map (
            O => \N__4895\,
            I => \C1_c\
        );

    \I__620\ : InMux
    port map (
            O => \N__4890\,
            I => \N__4887\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__4887\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__618\ : InMux
    port map (
            O => \N__4884\,
            I => \N__4880\
        );

    \I__617\ : InMux
    port map (
            O => \N__4883\,
            I => \N__4877\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__4880\,
            I => \N__4874\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__4877\,
            I => \N__4871\
        );

    \I__614\ : Span4Mux_v
    port map (
            O => \N__4874\,
            I => \N__4868\
        );

    \I__613\ : Span4Mux_h
    port map (
            O => \N__4871\,
            I => \N__4865\
        );

    \I__612\ : Sp12to4
    port map (
            O => \N__4868\,
            I => \N__4862\
        );

    \I__611\ : Span4Mux_v
    port map (
            O => \N__4865\,
            I => \N__4859\
        );

    \I__610\ : Span12Mux_h
    port map (
            O => \N__4862\,
            I => \N__4856\
        );

    \I__609\ : IoSpan4Mux
    port map (
            O => \N__4859\,
            I => \N__4853\
        );

    \I__608\ : Odrv12
    port map (
            O => \N__4856\,
            I => \TSn_c\
        );

    \I__607\ : Odrv4
    port map (
            O => \N__4853\,
            I => \TSn_c\
        );

    \I__606\ : InMux
    port map (
            O => \N__4848\,
            I => \N__4845\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__4845\,
            I => \N__4842\
        );

    \I__604\ : Span4Mux_h
    port map (
            O => \N__4842\,
            I => \N__4839\
        );

    \I__603\ : Span4Mux_v
    port map (
            O => \N__4839\,
            I => \N__4836\
        );

    \I__602\ : Odrv4
    port map (
            O => \N__4836\,
            I => \RAMSPACEn_c\
        );

    \I__601\ : InMux
    port map (
            O => \N__4833\,
            I => \N__4830\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__4830\,
            I => \N__4827\
        );

    \I__599\ : Span12Mux_v
    port map (
            O => \N__4827\,
            I => \N__4824\
        );

    \I__598\ : Odrv12
    port map (
            O => \N__4824\,
            I => \U712_CHIP_RAM.N_289\
        );

    \I__597\ : IoInMux
    port map (
            O => \N__4821\,
            I => \N__4818\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__4818\,
            I => \N__4815\
        );

    \I__595\ : Span4Mux_s1_v
    port map (
            O => \N__4815\,
            I => \N__4812\
        );

    \I__594\ : Span4Mux_v
    port map (
            O => \N__4812\,
            I => \N__4809\
        );

    \I__593\ : Span4Mux_v
    port map (
            O => \N__4809\,
            I => \N__4806\
        );

    \I__592\ : Span4Mux_v
    port map (
            O => \N__4806\,
            I => \N__4803\
        );

    \I__591\ : Odrv4
    port map (
            O => \N__4803\,
            I => \CMA_c_1\
        );

    \I__590\ : InMux
    port map (
            O => \N__4800\,
            I => \N__4797\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__4797\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\
        );

    \I__588\ : InMux
    port map (
            O => \N__4794\,
            I => \N__4791\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__4791\,
            I => \N__4788\
        );

    \I__586\ : Span12Mux_v
    port map (
            O => \N__4788\,
            I => \N__4785\
        );

    \I__585\ : Span12Mux_h
    port map (
            O => \N__4785\,
            I => \N__4782\
        );

    \I__584\ : Odrv12
    port map (
            O => \N__4782\,
            I => \A_c_3\
        );

    \I__583\ : InMux
    port map (
            O => \N__4779\,
            I => \N__4776\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__4776\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__581\ : CascadeMux
    port map (
            O => \N__4773\,
            I => \N__4770\
        );

    \I__580\ : InMux
    port map (
            O => \N__4770\,
            I => \N__4764\
        );

    \I__579\ : InMux
    port map (
            O => \N__4769\,
            I => \N__4764\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__4764\,
            I => \N__4761\
        );

    \I__577\ : Span12Mux_v
    port map (
            O => \N__4761\,
            I => \N__4758\
        );

    \I__576\ : Span12Mux_h
    port map (
            O => \N__4758\,
            I => \N__4755\
        );

    \I__575\ : Odrv12
    port map (
            O => \N__4755\,
            I => \A_c_10\
        );

    \I__574\ : InMux
    port map (
            O => \N__4752\,
            I => \N__4749\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__4749\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__572\ : InMux
    port map (
            O => \N__4746\,
            I => \N__4741\
        );

    \I__571\ : InMux
    port map (
            O => \N__4745\,
            I => \N__4736\
        );

    \I__570\ : InMux
    port map (
            O => \N__4744\,
            I => \N__4736\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__4741\,
            I => \U712_CHIP_RAM.N_208\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__4736\,
            I => \U712_CHIP_RAM.N_208\
        );

    \I__567\ : CEMux
    port map (
            O => \N__4731\,
            I => \N__4728\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__4728\,
            I => \N__4725\
        );

    \I__565\ : Odrv4
    port map (
            O => \N__4725\,
            I => \U712_CYCLE_TERM.N_217_i_0_en_0\
        );

    \I__564\ : IoInMux
    port map (
            O => \N__4722\,
            I => \N__4719\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__4719\,
            I => \N__4715\
        );

    \I__562\ : IoInMux
    port map (
            O => \N__4718\,
            I => \N__4712\
        );

    \I__561\ : Span12Mux_s1_v
    port map (
            O => \N__4715\,
            I => \N__4709\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__4712\,
            I => \N__4706\
        );

    \I__559\ : Span12Mux_v
    port map (
            O => \N__4709\,
            I => \N__4703\
        );

    \I__558\ : Span12Mux_s1_v
    port map (
            O => \N__4706\,
            I => \N__4700\
        );

    \I__557\ : Span12Mux_h
    port map (
            O => \N__4703\,
            I => \N__4694\
        );

    \I__556\ : Span12Mux_v
    port map (
            O => \N__4700\,
            I => \N__4694\
        );

    \I__555\ : InMux
    port map (
            O => \N__4699\,
            I => \N__4691\
        );

    \I__554\ : Odrv12
    port map (
            O => \N__4694\,
            I => \ASn_c\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__4691\,
            I => \ASn_c\
        );

    \I__552\ : InMux
    port map (
            O => \N__4686\,
            I => \N__4682\
        );

    \I__551\ : InMux
    port map (
            O => \N__4685\,
            I => \N__4679\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__4682\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4679\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__548\ : IoInMux
    port map (
            O => \N__4674\,
            I => \N__4671\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4671\,
            I => \N__4667\
        );

    \I__546\ : InMux
    port map (
            O => \N__4670\,
            I => \N__4664\
        );

    \I__545\ : Span4Mux_s1_v
    port map (
            O => \N__4667\,
            I => \N__4661\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__4664\,
            I => \N__4658\
        );

    \I__543\ : Sp12to4
    port map (
            O => \N__4661\,
            I => \N__4655\
        );

    \I__542\ : Span4Mux_v
    port map (
            O => \N__4658\,
            I => \N__4652\
        );

    \I__541\ : Span12Mux_h
    port map (
            O => \N__4655\,
            I => \N__4649\
        );

    \I__540\ : Sp12to4
    port map (
            O => \N__4652\,
            I => \N__4646\
        );

    \I__539\ : Span12Mux_v
    port map (
            O => \N__4649\,
            I => \N__4641\
        );

    \I__538\ : Span12Mux_h
    port map (
            O => \N__4646\,
            I => \N__4641\
        );

    \I__537\ : Span12Mux_v
    port map (
            O => \N__4641\,
            I => \N__4638\
        );

    \I__536\ : Odrv12
    port map (
            O => \N__4638\,
            I => \RAMENn_c\
        );

    \I__535\ : CascadeMux
    port map (
            O => \N__4635\,
            I => \U712_REG_SM.N_270_cascade_\
        );

    \I__534\ : InMux
    port map (
            O => \N__4632\,
            I => \N__4629\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__4629\,
            I => \N__4626\
        );

    \I__532\ : Odrv12
    port map (
            O => \N__4626\,
            I => \U712_CHIP_RAM.CLK_EN_6_0_a2_2\
        );

    \I__531\ : CascadeMux
    port map (
            O => \N__4623\,
            I => \N__4620\
        );

    \I__530\ : InMux
    port map (
            O => \N__4620\,
            I => \N__4617\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__4617\,
            I => \N__4614\
        );

    \I__528\ : Odrv4
    port map (
            O => \N__4614\,
            I => \U712_CHIP_RAM.CLK_EN_6_0_a2_1\
        );

    \I__527\ : CascadeMux
    port map (
            O => \N__4611\,
            I => \U712_CHIP_RAM.CLK_EN_6_0_cascade_\
        );

    \I__526\ : IoInMux
    port map (
            O => \N__4608\,
            I => \N__4605\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__4605\,
            I => \N__4602\
        );

    \I__524\ : Span12Mux_s7_h
    port map (
            O => \N__4602\,
            I => \N__4599\
        );

    \I__523\ : Span12Mux_h
    port map (
            O => \N__4599\,
            I => \N__4595\
        );

    \I__522\ : InMux
    port map (
            O => \N__4598\,
            I => \N__4592\
        );

    \I__521\ : Odrv12
    port map (
            O => \N__4595\,
            I => \CLK_EN_c\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__4592\,
            I => \CLK_EN_c\
        );

    \I__519\ : InMux
    port map (
            O => \N__4587\,
            I => \N__4584\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__4584\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0\
        );

    \I__517\ : InMux
    port map (
            O => \N__4581\,
            I => \N__4578\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__4578\,
            I => \U712_CHIP_RAM.N_385\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__4575\,
            I => \U712_CHIP_RAM.N_338_cascade_\
        );

    \I__514\ : CascadeMux
    port map (
            O => \N__4572\,
            I => \U712_CHIP_RAM.N_305_cascade_\
        );

    \I__513\ : CascadeMux
    port map (
            O => \N__4569\,
            I => \U712_CHIP_RAM.N_239_cascade_\
        );

    \I__512\ : CascadeMux
    port map (
            O => \N__4566\,
            I => \N__4563\
        );

    \I__511\ : InMux
    port map (
            O => \N__4563\,
            I => \N__4559\
        );

    \I__510\ : InMux
    port map (
            O => \N__4562\,
            I => \N__4556\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__4559\,
            I => \N__4553\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__4556\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__507\ : Odrv4
    port map (
            O => \N__4553\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__506\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4543\
        );

    \I__505\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4540\
        );

    \I__504\ : InMux
    port map (
            O => \N__4546\,
            I => \N__4537\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4543\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__4540\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__4537\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\
        );

    \I__500\ : InMux
    port map (
            O => \N__4530\,
            I => \N__4527\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4527\,
            I => \U712_CHIP_RAM.N_387\
        );

    \I__498\ : CascadeMux
    port map (
            O => \N__4524\,
            I => \U712_CHIP_RAM.N_385_cascade_\
        );

    \I__497\ : CascadeMux
    port map (
            O => \N__4521\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_cascade_\
        );

    \I__496\ : CascadeMux
    port map (
            O => \N__4518\,
            I => \N__4515\
        );

    \I__495\ : InMux
    port map (
            O => \N__4515\,
            I => \N__4512\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4512\,
            I => \U712_CHIP_RAM.N_223\
        );

    \I__493\ : CascadeMux
    port map (
            O => \N__4509\,
            I => \U712_CHIP_RAM.N_335_cascade_\
        );

    \I__492\ : CascadeMux
    port map (
            O => \N__4506\,
            I => \U712_CHIP_RAM.N_342_cascade_\
        );

    \I__491\ : InMux
    port map (
            O => \N__4503\,
            I => \N__4500\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__4500\,
            I => \N__4497\
        );

    \I__489\ : Span4Mux_v
    port map (
            O => \N__4497\,
            I => \N__4494\
        );

    \I__488\ : Span4Mux_h
    port map (
            O => \N__4494\,
            I => \N__4491\
        );

    \I__487\ : Odrv4
    port map (
            O => \N__4491\,
            I => \TACK_EN_i_ess\
        );

    \I__486\ : IoInMux
    port map (
            O => \N__4488\,
            I => \N__4485\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__4485\,
            I => \N__4482\
        );

    \I__484\ : IoSpan4Mux
    port map (
            O => \N__4482\,
            I => \N__4479\
        );

    \I__483\ : Span4Mux_s0_h
    port map (
            O => \N__4479\,
            I => \N__4476\
        );

    \I__482\ : Sp12to4
    port map (
            O => \N__4476\,
            I => \N__4473\
        );

    \I__481\ : Span12Mux_s11_h
    port map (
            O => \N__4473\,
            I => \N__4469\
        );

    \I__480\ : InMux
    port map (
            O => \N__4472\,
            I => \N__4466\
        );

    \I__479\ : Odrv12
    port map (
            O => \N__4469\,
            I => \TACK_OUTn\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__4466\,
            I => \TACK_OUTn\
        );

    \I__477\ : InMux
    port map (
            O => \N__4461\,
            I => \N__4458\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__4458\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\
        );

    \I__475\ : InMux
    port map (
            O => \N__4455\,
            I => \N__4452\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4452\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\
        );

    \I__473\ : IoInMux
    port map (
            O => \N__4449\,
            I => \N__4446\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__4446\,
            I => \N__4443\
        );

    \I__471\ : Span12Mux_s7_h
    port map (
            O => \N__4443\,
            I => \N__4440\
        );

    \I__470\ : Span12Mux_h
    port map (
            O => \N__4440\,
            I => \N__4437\
        );

    \I__469\ : Odrv12
    port map (
            O => \N__4437\,
            I => \CMA_c_5\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__4434\,
            I => \U712_CHIP_RAM.N_387_cascade_\
        );

    \I__467\ : InMux
    port map (
            O => \N__4431\,
            I => \N__4428\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__4428\,
            I => \N__4424\
        );

    \I__465\ : InMux
    port map (
            O => \N__4427\,
            I => \N__4421\
        );

    \I__464\ : Span4Mux_h
    port map (
            O => \N__4424\,
            I => \N__4416\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__4421\,
            I => \N__4416\
        );

    \I__462\ : Span4Mux_v
    port map (
            O => \N__4416\,
            I => \N__4413\
        );

    \I__461\ : Span4Mux_h
    port map (
            O => \N__4413\,
            I => \N__4410\
        );

    \I__460\ : Sp12to4
    port map (
            O => \N__4410\,
            I => \N__4407\
        );

    \I__459\ : Odrv12
    port map (
            O => \N__4407\,
            I => \AWEn_c\
        );

    \I__458\ : InMux
    port map (
            O => \N__4404\,
            I => \N__4395\
        );

    \I__457\ : InMux
    port map (
            O => \N__4403\,
            I => \N__4395\
        );

    \I__456\ : InMux
    port map (
            O => \N__4402\,
            I => \N__4395\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__4395\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__454\ : CascadeMux
    port map (
            O => \N__4392\,
            I => \U712_CHIP_RAM.N_186_cascade_\
        );

    \I__453\ : InMux
    port map (
            O => \N__4389\,
            I => \N__4386\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__4386\,
            I => \N__4383\
        );

    \I__451\ : Odrv4
    port map (
            O => \N__4383\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__450\ : InMux
    port map (
            O => \N__4380\,
            I => \N__4377\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__4377\,
            I => \U712_CHIP_RAM.DBENn_8_0\
        );

    \I__448\ : InMux
    port map (
            O => \N__4374\,
            I => \N__4371\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__4371\,
            I => \N__4368\
        );

    \I__446\ : Odrv4
    port map (
            O => \N__4368\,
            I => \U712_CHIP_RAM.N_341\
        );

    \I__445\ : CascadeMux
    port map (
            O => \N__4365\,
            I => \U712_CHIP_RAM.N_341_cascade_\
        );

    \I__444\ : InMux
    port map (
            O => \N__4362\,
            I => \N__4359\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__4359\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_a2_0\
        );

    \I__442\ : InMux
    port map (
            O => \N__4356\,
            I => \N__4352\
        );

    \I__441\ : InMux
    port map (
            O => \N__4355\,
            I => \N__4349\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__4352\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__4349\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0\
        );

    \I__438\ : CEMux
    port map (
            O => \N__4344\,
            I => \N__4341\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__4341\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0\
        );

    \I__436\ : InMux
    port map (
            O => \N__4338\,
            I => \N__4335\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__4335\,
            I => \N__4332\
        );

    \I__434\ : Span4Mux_h
    port map (
            O => \N__4332\,
            I => \N__4329\
        );

    \I__433\ : Span4Mux_v
    port map (
            O => \N__4329\,
            I => \N__4326\
        );

    \I__432\ : Sp12to4
    port map (
            O => \N__4326\,
            I => \N__4323\
        );

    \I__431\ : Odrv12
    port map (
            O => \N__4323\,
            I => \A_c_20\
        );

    \I__430\ : InMux
    port map (
            O => \N__4320\,
            I => \N__4316\
        );

    \I__429\ : CascadeMux
    port map (
            O => \N__4319\,
            I => \N__4313\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__4316\,
            I => \N__4310\
        );

    \I__427\ : InMux
    port map (
            O => \N__4313\,
            I => \N__4307\
        );

    \I__426\ : Span4Mux_h
    port map (
            O => \N__4310\,
            I => \N__4304\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__4307\,
            I => \N__4301\
        );

    \I__424\ : Odrv4
    port map (
            O => \N__4304\,
            I => \DBRn_c_i\
        );

    \I__423\ : Odrv4
    port map (
            O => \N__4301\,
            I => \DBRn_c_i\
        );

    \I__422\ : IoInMux
    port map (
            O => \N__4296\,
            I => \N__4293\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__4293\,
            I => \N__4290\
        );

    \I__420\ : Span12Mux_s11_v
    port map (
            O => \N__4290\,
            I => \N__4287\
        );

    \I__419\ : Odrv12
    port map (
            O => \N__4287\,
            I => \VBENn_c\
        );

    \I__418\ : InMux
    port map (
            O => \N__4284\,
            I => \N__4281\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__4281\,
            I => \N__4278\
        );

    \I__416\ : Span4Mux_h
    port map (
            O => \N__4278\,
            I => \N__4275\
        );

    \I__415\ : Sp12to4
    port map (
            O => \N__4275\,
            I => \N__4272\
        );

    \I__414\ : Span12Mux_v
    port map (
            O => \N__4272\,
            I => \N__4269\
        );

    \I__413\ : Odrv12
    port map (
            O => \N__4269\,
            I => \A_c_14\
        );

    \I__412\ : InMux
    port map (
            O => \N__4266\,
            I => \N__4263\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__4263\,
            I => \N__4260\
        );

    \I__410\ : Span4Mux_h
    port map (
            O => \N__4260\,
            I => \N__4257\
        );

    \I__409\ : Span4Mux_v
    port map (
            O => \N__4257\,
            I => \N__4254\
        );

    \I__408\ : Sp12to4
    port map (
            O => \N__4254\,
            I => \N__4251\
        );

    \I__407\ : Odrv12
    port map (
            O => \N__4251\,
            I => \A_c_7\
        );

    \I__406\ : CascadeMux
    port map (
            O => \N__4248\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5_cascade_\
        );

    \I__405\ : CascadeMux
    port map (
            O => \N__4245\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_\
        );

    \I__404\ : IoInMux
    port map (
            O => \N__4242\,
            I => \N__4239\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__4239\,
            I => \N__4236\
        );

    \I__402\ : Span4Mux_s3_v
    port map (
            O => \N__4236\,
            I => \N__4233\
        );

    \I__401\ : Span4Mux_v
    port map (
            O => \N__4233\,
            I => \N__4230\
        );

    \I__400\ : Sp12to4
    port map (
            O => \N__4230\,
            I => \N__4227\
        );

    \I__399\ : Span12Mux_s11_h
    port map (
            O => \N__4227\,
            I => \N__4223\
        );

    \I__398\ : InMux
    port map (
            O => \N__4226\,
            I => \N__4220\
        );

    \I__397\ : Odrv12
    port map (
            O => \N__4223\,
            I => \LATCH_CLK_c\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__4220\,
            I => \LATCH_CLK_c\
        );

    \I__395\ : InMux
    port map (
            O => \N__4215\,
            I => \N__4212\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__4212\,
            I => \U712_CHIP_RAM.LATCH_CLK_RNOZ0Z_0\
        );

    \I__393\ : IoInMux
    port map (
            O => \N__4209\,
            I => \N__4206\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__4206\,
            I => \N__4203\
        );

    \I__391\ : Span4Mux_s3_v
    port map (
            O => \N__4203\,
            I => \N__4200\
        );

    \I__390\ : Span4Mux_v
    port map (
            O => \N__4200\,
            I => \N__4197\
        );

    \I__389\ : Span4Mux_v
    port map (
            O => \N__4197\,
            I => \N__4194\
        );

    \I__388\ : Span4Mux_v
    port map (
            O => \N__4194\,
            I => \N__4190\
        );

    \I__387\ : InMux
    port map (
            O => \N__4193\,
            I => \N__4187\
        );

    \I__386\ : Odrv4
    port map (
            O => \N__4190\,
            I => \DBDIR_c\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__4187\,
            I => \DBDIR_c\
        );

    \I__384\ : IoInMux
    port map (
            O => \N__4182\,
            I => \N__4179\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__4179\,
            I => \N__4176\
        );

    \I__382\ : Odrv12
    port map (
            O => \N__4176\,
            I => \DBRn_c_i_0\
        );

    \I__381\ : IoInMux
    port map (
            O => \N__4173\,
            I => \N__4170\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__4170\,
            I => \N__4167\
        );

    \I__379\ : Span4Mux_s3_v
    port map (
            O => \N__4167\,
            I => \N__4164\
        );

    \I__378\ : Span4Mux_h
    port map (
            O => \N__4164\,
            I => \N__4161\
        );

    \I__377\ : Odrv4
    port map (
            O => \N__4161\,
            I => \CLK80_PLL_i_i\
        );

    \I__376\ : IoInMux
    port map (
            O => \N__4158\,
            I => \N__4155\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__4155\,
            I => \N__4152\
        );

    \I__374\ : Span4Mux_s2_h
    port map (
            O => \N__4152\,
            I => \N__4149\
        );

    \I__373\ : Span4Mux_h
    port map (
            O => \N__4149\,
            I => \N__4146\
        );

    \I__372\ : Span4Mux_v
    port map (
            O => \N__4146\,
            I => \N__4143\
        );

    \I__371\ : Odrv4
    port map (
            O => \N__4143\,
            I => \N_861_i\
        );

    \I__370\ : InMux
    port map (
            O => \N__4140\,
            I => \N__4136\
        );

    \I__369\ : InMux
    port map (
            O => \N__4139\,
            I => \N__4133\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__4136\,
            I => \N__4128\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__4133\,
            I => \N__4128\
        );

    \I__366\ : Span4Mux_v
    port map (
            O => \N__4128\,
            I => \N__4125\
        );

    \I__365\ : Span4Mux_h
    port map (
            O => \N__4125\,
            I => \N__4122\
        );

    \I__364\ : Sp12to4
    port map (
            O => \N__4122\,
            I => \N__4119\
        );

    \I__363\ : Span12Mux_v
    port map (
            O => \N__4119\,
            I => \N__4116\
        );

    \I__362\ : Odrv12
    port map (
            O => \N__4116\,
            I => \DBRn_c\
        );

    \I__361\ : IoInMux
    port map (
            O => \N__4113\,
            I => \N__4110\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__4110\,
            I => \N__4107\
        );

    \I__359\ : Span4Mux_s0_v
    port map (
            O => \N__4107\,
            I => \N__4104\
        );

    \I__358\ : Span4Mux_v
    port map (
            O => \N__4104\,
            I => \N__4101\
        );

    \I__357\ : Sp12to4
    port map (
            O => \N__4101\,
            I => \N__4098\
        );

    \I__356\ : Span12Mux_h
    port map (
            O => \N__4098\,
            I => \N__4095\
        );

    \I__355\ : Span12Mux_v
    port map (
            O => \N__4095\,
            I => \N__4092\
        );

    \I__354\ : Odrv12
    port map (
            O => \N__4092\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            I => \N__5467\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__5469\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            I => \N__5470\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            I => \N__5465\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            I => \N__5466\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            I => \N__5468\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__5471\
        );

    \INVU712_CHIP_RAM.DMA_A20C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A20C_net\,
            I => \N__5472\
        );

    \IN_MUX_bfv_10_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_12_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_15_0_\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4925\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7722\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4182\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7308\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10017\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4320\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_3_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10707\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_obuft_RNO_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4503\,
            lcout => \N_861_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBRn_ibuf_RNIBAB_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4139\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_0_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4140\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10693\,
            ce => 'H',
            sr => \N__9991\
        );

    \U712_CHIP_RAM.DMA_A20_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__10325\,
            in1 => \N__9212\,
            in2 => \N__4319\,
            in3 => \N__5009\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A20C_net\,
            ce => 'H',
            sr => \N__9984\
        );

    \U712_BUFFERS.un1_VBENn_0_a2_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8821\,
            in2 => \_gnd_net_\,
            in3 => \N__9842\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4284\,
            in1 => \N__4266\,
            in2 => \_gnd_net_\,
            in3 => \N__9396\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9397\,
            in1 => \N__8820\,
            in2 => \N__4248\,
            in3 => \N__8937\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__4547\,
            in1 => \N__4374\,
            in2 => \N__6948\,
            in3 => \N__6270\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100010101000"
        )
    port map (
            in0 => \N__8194\,
            in1 => \N__4226\,
            in2 => \N__4245\,
            in3 => \N__4215\,
            lcout => \LATCH_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10679\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7179\,
            in2 => \_gnd_net_\,
            in3 => \N__5613\,
            lcout => \U712_CHIP_RAM.LATCH_CLK_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001001010"
        )
    port map (
            in0 => \N__10802\,
            in1 => \N__10952\,
            in2 => \N__9402\,
            in3 => \N__8787\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBDIR_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__4427\,
            in1 => \N__4193\,
            in2 => \_gnd_net_\,
            in3 => \N__4548\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10684\,
            ce => 'H',
            sr => \N__9978\
        );

    \U712_CHIP_RAM.DBENn_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__5559\,
            in1 => \N__4356\,
            in2 => \_gnd_net_\,
            in3 => \N__4380\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10684\,
            ce => 'H',
            sr => \N__9978\
        );

    \DBR_SYNC_1_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4389\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10684\,
            ce => 'H',
            sr => \N__9978\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10016\,
            in2 => \_gnd_net_\,
            in3 => \N__4355\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6236\,
            in1 => \N__6166\,
            in2 => \_gnd_net_\,
            in3 => \N__8922\,
            lcout => \U712_CHIP_RAM.DBENn_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_0_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__7175\,
            in1 => \N__7050\,
            in2 => \N__6360\,
            in3 => \N__11096\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI8MK44_1_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__4746\,
            in1 => \N__7051\,
            in2 => \N__7182\,
            in3 => \N__6921\,
            lcout => \U712_CHIP_RAM.N_341\,
            ltout => \U712_CHIP_RAM.N_341_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIBTHEC_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__6922\,
            in1 => \N__4546\,
            in2 => \N__4365\,
            in3 => \N__4362\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6171\,
            in1 => \N__6492\,
            in2 => \N__6252\,
            in3 => \N__6598\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10694\,
            ce => \N__4344\,
            sr => \N__9965\
        );

    \U712_CHIP_RAM.BANK0_RNO_3_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10326\,
            in2 => \_gnd_net_\,
            in3 => \N__4338\,
            lcout => \U712_CHIP_RAM.BANK0_RNOZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__8195\,
            in1 => \N__7386\,
            in2 => \_gnd_net_\,
            in3 => \N__7416\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10698\,
            ce => \N__4731\,
            sr => \N__9958\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111100011111010"
        )
    port map (
            in0 => \N__4472\,
            in1 => \N__8619\,
            in2 => \N__5241\,
            in3 => \N__7455\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10701\,
            ce => 'H',
            sr => \N__9950\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4800\,
            in1 => \N__4461\,
            in2 => \_gnd_net_\,
            in3 => \N__4455\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10669\,
            ce => \N__10565\,
            sr => \N__9985\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__6591\,
            in1 => \N__4403\,
            in2 => \N__6789\,
            in3 => \N__8435\,
            lcout => \U712_CHIP_RAM.N_387\,
            ltout => \U712_CHIP_RAM.N_387_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIURFN4_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6235\,
            in2 => \N__4434\,
            in3 => \N__6162\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010100110101"
        )
    port map (
            in0 => \N__11341\,
            in1 => \N__4431\,
            in2 => \N__6599\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_223\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011100000"
        )
    port map (
            in0 => \N__4404\,
            in1 => \N__4833\,
            in2 => \N__8213\,
            in3 => \N__8778\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10674\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4402\,
            in2 => \_gnd_net_\,
            in3 => \N__8434\,
            lcout => \U712_CHIP_RAM.N_186\,
            ltout => \U712_CHIP_RAM.N_186_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIHJRU1_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__8202\,
            in1 => \N__6590\,
            in2 => \N__4392\,
            in3 => \N__6782\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_3_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__8777\,
            in1 => \N__7174\,
            in2 => \_gnd_net_\,
            in3 => \N__7059\,
            lcout => \U712_CHIP_RAM.CLK_EN_6_0_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_2_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__11100\,
            in1 => \N__6674\,
            in2 => \_gnd_net_\,
            in3 => \N__6361\,
            lcout => \U712_CHIP_RAM.CLK_EN_6_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6563\,
            in1 => \N__6491\,
            in2 => \N__6246\,
            in3 => \N__6135\,
            lcout => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010100000"
        )
    port map (
            in0 => \N__7157\,
            in1 => \N__7019\,
            in2 => \N__6368\,
            in3 => \N__11094\,
            lcout => \U712_CHIP_RAM.N_385\,
            ltout => \U712_CHIP_RAM.N_385_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__4530\,
            in1 => \N__6855\,
            in2 => \N__4524\,
            in3 => \N__6937\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__8196\,
            in1 => \N__8788\,
            in2 => \N__4521\,
            in3 => \N__5024\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__11095\,
            in1 => \N__8197\,
            in2 => \N__4518\,
            in3 => \N__4562\,
            lcout => \WRITE_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_3_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7156\,
            in1 => \N__6343\,
            in2 => \N__6680\,
            in3 => \N__7018\,
            lcout => \U712_CHIP_RAM.N_335\,
            ltout => \U712_CHIP_RAM.N_335_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU2TJ3_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6490\,
            in2 => \N__4509\,
            in3 => \N__6134\,
            lcout => \U712_CHIP_RAM.N_342\,
            ltout => \U712_CHIP_RAM.N_342_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIPCS25_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011010000"
        )
    port map (
            in0 => \N__4953\,
            in1 => \N__6564\,
            in2 => \N__4506\,
            in3 => \N__6787\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5880\,
            in1 => \N__4632\,
            in2 => \N__4623\,
            in3 => \N__6140\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CLK_EN_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000111110101010"
        )
    port map (
            in0 => \N__4598\,
            in1 => \_gnd_net_\,
            in2 => \N__4611\,
            in3 => \N__4587\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10685\,
            ce => 'H',
            sr => \N__9966\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7155\,
            in1 => \N__4745\,
            in2 => \N__6943\,
            in3 => \N__7044\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5O1M2_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__6662\,
            in1 => \N__5879\,
            in2 => \N__6161\,
            in3 => \N__6480\,
            lcout => \U712_CHIP_RAM.N_338\,
            ltout => \U712_CHIP_RAM.N_338_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITIV55_0_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011100000"
        )
    port map (
            in0 => \N__4581\,
            in1 => \N__7043\,
            in2 => \N__4575\,
            in3 => \N__4744\,
            lcout => \U712_CHIP_RAM.N_305\,
            ltout => \U712_CHIP_RAM.N_305_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSRL5_0_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4572\,
            in3 => \N__8161\,
            lcout => \U712_CHIP_RAM.N_239\,
            ltout => \U712_CHIP_RAM.N_239_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQVN9G_3_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__5082\,
            in1 => \N__5659\,
            in2 => \N__4569\,
            in3 => \N__5538\,
            lcout => \U712_CHIP_RAM.N_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIL1QU_2_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8188\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6332\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__5165\,
            in1 => \N__5049\,
            in2 => \N__4566\,
            in3 => \N__8187\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10690\,
            ce => \N__5717\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8HNG_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5602\,
            in2 => \_gnd_net_\,
            in3 => \N__6331\,
            lcout => \U712_CHIP_RAM.N_208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7060\,
            in1 => \N__8186\,
            in2 => \_gnd_net_\,
            in3 => \N__7208\,
            lcout => \U712_CHIP_RAM.N_304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6342\,
            in1 => \N__5883\,
            in2 => \_gnd_net_\,
            in3 => \N__5499\,
            lcout => \U712_CHIP_RAM.N_269\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10015\,
            in2 => \_gnd_net_\,
            in3 => \N__5109\,
            lcout => \U712_CYCLE_TERM.N_217_i_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010001000100011"
        )
    port map (
            in0 => \N__5256\,
            in1 => \N__7353\,
            in2 => \N__8352\,
            in3 => \N__5675\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10695\,
            ce => 'H',
            sr => \N__9951\
        );

    \U712_REG_SM.ASn_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101100001000"
        )
    port map (
            in0 => \N__8302\,
            in1 => \N__5250\,
            in2 => \N__8418\,
            in3 => \N__4699\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10695\,
            ce => 'H',
            sr => \N__9951\
        );

    \U712_REG_SM.START_RST_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__4686\,
            in1 => \N__5103\,
            in2 => \_gnd_net_\,
            in3 => \N__6051\,
            lcout => \U712_REG_SM.START_RSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10695\,
            ce => 'H',
            sr => \N__9951\
        );

    \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4685\,
            in2 => \_gnd_net_\,
            in3 => \N__5271\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_270_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100010"
        )
    port map (
            in0 => \N__8217\,
            in1 => \N__4670\,
            in2 => \N__4635\,
            in3 => \N__4884\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10699\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8216\,
            in2 => \_gnd_net_\,
            in3 => \N__5220\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10699\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_1_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4890\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10702\,
            ce => 'H',
            sr => \N__9945\
        );

    \U712_REG_SM.C1_SYNC_0_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4926\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10703\,
            ce => 'H',
            sr => \N__9944\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4883\,
            in2 => \_gnd_net_\,
            in3 => \N__4848\,
            lcout => \U712_CHIP_RAM.N_289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4752\,
            in1 => \N__4779\,
            in2 => \_gnd_net_\,
            in3 => \N__5433\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10666\,
            ce => \N__10556\,
            sr => \N__9979\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011111111"
        )
    port map (
            in0 => \N__8774\,
            in1 => \N__10956\,
            in2 => \N__10819\,
            in3 => \N__9398\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4794\,
            in1 => \N__8773\,
            in2 => \_gnd_net_\,
            in3 => \N__8658\,
            lcout => \U712_CHIP_RAM.N_134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__8775\,
            in1 => \N__4769\,
            in2 => \N__7957\,
            in3 => \N__8639\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011101100"
        )
    port map (
            in0 => \N__8198\,
            in1 => \N__6575\,
            in2 => \N__7869\,
            in3 => \N__5623\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10670\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110111011"
        )
    port map (
            in0 => \N__8640\,
            in1 => \N__7948\,
            in2 => \N__4773\,
            in3 => \N__8776\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_1_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101010000"
        )
    port map (
            in0 => \N__5037\,
            in1 => \N__4959\,
            in2 => \N__5025\,
            in3 => \N__5010\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.BANK0_RNOZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__4970\,
            in1 => \N__4995\,
            in2 => \N__4989\,
            in3 => \N__4938\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10675\,
            ce => 'H',
            sr => \N__9967\
        );

    \U712_CHIP_RAM.BANK0_RNO_4_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__6233\,
            in1 => \N__6152\,
            in2 => \_gnd_net_\,
            in3 => \N__6565\,
            lcout => \U712_CHIP_RAM.BANK0_RNOZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_2_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000100"
        )
    port map (
            in0 => \N__4952\,
            in1 => \N__6234\,
            in2 => \N__6583\,
            in3 => \N__6788\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_0_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_0_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4941\,
            in3 => \N__5660\,
            lcout => \U712_CHIP_RAM.N_306\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5888\,
            in1 => \N__6479\,
            in2 => \_gnd_net_\,
            in3 => \N__6136\,
            lcout => \U712_CHIP_RAM.N_333\,
            ltout => \U712_CHIP_RAM.N_333_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI27TJ3_3_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6697\,
            in2 => \N__4932\,
            in3 => \N__6673\,
            lcout => \U712_CHIP_RAM.N_386\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6661\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7025\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_0_0_a2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_4_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6698\,
            in1 => \N__5881\,
            in2 => \N__4929\,
            in3 => \N__6142\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER18\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI7UUV6_4_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110000"
        )
    port map (
            in0 => \N__6143\,
            in1 => \_gnd_net_\,
            in2 => \N__5085\,
            in3 => \N__6232\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000111010"
        )
    port map (
            in0 => \N__5061\,
            in1 => \N__5076\,
            in2 => \N__5169\,
            in3 => \N__5070\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10681\,
            ce => \N__5713\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6660\,
            in1 => \N__7144\,
            in2 => \_gnd_net_\,
            in3 => \N__7024\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_0_0_a2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQGOH4_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__6481\,
            in1 => \N__5534\,
            in2 => \N__5064\,
            in3 => \N__6141\,
            lcout => \U712_CHIP_RAM.N_202\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__5120\,
            in1 => \N__5183\,
            in2 => \_gnd_net_\,
            in3 => \N__5198\,
            lcout => \U712_CHIP_RAM.N_180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7045\,
            in2 => \_gnd_net_\,
            in3 => \N__5055\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \bfn_10_12_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5158\,
            in1 => \N__7154\,
            in2 => \_gnd_net_\,
            in3 => \N__5052\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__10686\,
            ce => \N__5718\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6355\,
            in2 => \_gnd_net_\,
            in3 => \N__5043\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5159\,
            in1 => \N__6675\,
            in2 => \_gnd_net_\,
            in3 => \N__5040\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__10686\,
            ce => \N__5718\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5156\,
            in1 => \N__5884\,
            in2 => \_gnd_net_\,
            in3 => \N__5202\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__10686\,
            ce => \N__5718\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5160\,
            in1 => \N__5199\,
            in2 => \_gnd_net_\,
            in3 => \N__5187\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__10686\,
            ce => \N__5718\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5157\,
            in1 => \N__5184\,
            in2 => \_gnd_net_\,
            in3 => \N__5172\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__10686\,
            ce => \N__5718\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5161\,
            in1 => \N__5121\,
            in2 => \_gnd_net_\,
            in3 => \N__5124\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10686\,
            ce => \N__5718\,
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010101010"
        )
    port map (
            in0 => \N__7466\,
            in1 => \N__8190\,
            in2 => \N__7415\,
            in3 => \N__7385\,
            lcout => \U712_CYCLE_TERM.N_217_i_0_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.START_RST_RNO_0_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5097\,
            in1 => \N__5273\,
            in2 => \N__8310\,
            in3 => \N__8413\,
            lcout => \U712_REG_SM.START_RST_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__5272\,
            in1 => \N__5096\,
            in2 => \N__6054\,
            in3 => \N__8300\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_285_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__8301\,
            in1 => \N__8191\,
            in2 => \N__5088\,
            in3 => \N__8414\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10691\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__5283\,
            in1 => \N__8189\,
            in2 => \_gnd_net_\,
            in3 => \N__6470\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10691\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6732\,
            in1 => \N__5274\,
            in2 => \_gnd_net_\,
            in3 => \N__8346\,
            lcout => \U712_REG_SM.STATE_COUNT_srsts_i_0_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_RNO_0_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6047\,
            in1 => \N__6733\,
            in2 => \_gnd_net_\,
            in3 => \N__8296\,
            lcout => \U712_REG_SM.N_222\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__8613\,
            in1 => \N__8193\,
            in2 => \_gnd_net_\,
            in3 => \N__7451\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5240\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8214\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5484\,
            in1 => \N__5297\,
            in2 => \_gnd_net_\,
            in3 => \N__5312\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101010001010"
        )
    port map (
            in0 => \N__8192\,
            in1 => \N__5345\,
            in2 => \N__5244\,
            in3 => \N__5208\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5239\,
            in2 => \_gnd_net_\,
            in3 => \N__5219\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__5360\,
            in1 => \N__5390\,
            in2 => \N__5331\,
            in3 => \N__5375\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__8412\,
            in1 => \N__8486\,
            in2 => \_gnd_net_\,
            in3 => \N__8276\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_284_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__7348\,
            in1 => \N__5904\,
            in2 => \N__5394\,
            in3 => \N__8215\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5391\,
            in2 => \_gnd_net_\,
            in3 => \N__5379\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__5464\,
            ce => 'H',
            sr => \N__7494\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5376\,
            in2 => \_gnd_net_\,
            in3 => \N__5364\,
            lcout => \U712_CHIP_RAM.REFRESH5lto1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__5464\,
            ce => 'H',
            sr => \N__7494\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5361\,
            in2 => \_gnd_net_\,
            in3 => \N__5349\,
            lcout => \U712_CHIP_RAM.REFRESH5lto2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__5464\,
            ce => 'H',
            sr => \N__7494\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5346\,
            in2 => \_gnd_net_\,
            in3 => \N__5334\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__5464\,
            ce => 'H',
            sr => \N__7494\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5330\,
            in2 => \_gnd_net_\,
            in3 => \N__5316\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__5464\,
            ce => 'H',
            sr => \N__7494\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5313\,
            in2 => \_gnd_net_\,
            in3 => \N__5301\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__5464\,
            ce => 'H',
            sr => \N__7494\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5298\,
            in2 => \_gnd_net_\,
            in3 => \N__5286\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__5464\,
            ce => 'H',
            sr => \N__7494\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5483\,
            in2 => \_gnd_net_\,
            in3 => \N__5487\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5464\,
            ce => 'H',
            sr => \N__7494\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__7663\,
            in1 => \N__9362\,
            in2 => \_gnd_net_\,
            in3 => \N__7612\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_0_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5579\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5627\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__9363\,
            in1 => \N__10803\,
            in2 => \_gnd_net_\,
            in3 => \N__5439\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_116_i_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__11286\,
            in1 => \N__5780\,
            in2 => \N__7737\,
            in3 => \N__8810\,
            lcout => \N_116_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_2_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7158\,
            in2 => \_gnd_net_\,
            in3 => \N__6362\,
            lcout => \U712_CHIP_RAM.N_207\,
            ltout => \U712_CHIP_RAM.N_207_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_5_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5403\,
            in3 => \N__8809\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__11132\,
            in1 => \N__6679\,
            in2 => \N__5400\,
            in3 => \N__7049\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__5523\,
            in1 => \N__5889\,
            in2 => \N__5397\,
            in3 => \N__6160\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10671\,
            ce => \N__5634\,
            sr => \N__9959\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__6659\,
            in1 => \N__7022\,
            in2 => \N__5661\,
            in3 => \N__5517\,
            lcout => \U712_CHIP_RAM.N_262\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__7021\,
            in1 => \N__7152\,
            in2 => \N__6369\,
            in3 => \N__6941\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_310_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__6942\,
            in1 => \N__6263\,
            in2 => \N__5640\,
            in3 => \N__7204\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10014\,
            in1 => \_gnd_net_\,
            in2 => \N__5637\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__5628\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5578\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__7023\,
            in1 => \N__11137\,
            in2 => \N__6501\,
            in3 => \N__6159\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_3_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6658\,
            in1 => \N__7133\,
            in2 => \_gnd_net_\,
            in3 => \N__7020\,
            lcout => \U712_CHIP_RAM.N_334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__8830\,
            in1 => \N__11136\,
            in2 => \_gnd_net_\,
            in3 => \N__7153\,
            lcout => \U712_CHIP_RAM.N_297\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIGCGV5_4_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__5878\,
            in1 => \N__5513\,
            in2 => \_gnd_net_\,
            in3 => \N__5498\,
            lcout => \U712_CHIP_RAM.N_294\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNISAAQ_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5876\,
            in2 => \_gnd_net_\,
            in3 => \N__6463\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERlde_0_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001001010000"
        )
    port map (
            in0 => \N__6359\,
            in1 => \N__6666\,
            in2 => \N__7173\,
            in3 => \N__7039\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_184_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_4_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6145\,
            in1 => \N__5685\,
            in2 => \N__5739\,
            in3 => \N__5877\,
            lcout => \U712_CHIP_RAM.N_261\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000001"
        )
    port map (
            in0 => \N__6069\,
            in1 => \N__5736\,
            in2 => \N__6825\,
            in3 => \N__7661\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10682\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_3_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6144\,
            in1 => \N__6247\,
            in2 => \_gnd_net_\,
            in3 => \N__8115\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_392_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4TF5A_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__5727\,
            in1 => \N__6888\,
            in2 => \N__5721\,
            in3 => \N__6869\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__8347\,
            in1 => \N__6731\,
            in2 => \N__5679\,
            in3 => \N__8127\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10687\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8478\,
            in2 => \_gnd_net_\,
            in3 => \N__6041\,
            lcout => \U712_REG_SM.N_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__8126\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6464\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__8304\,
            in1 => \N__6730\,
            in2 => \_gnd_net_\,
            in3 => \N__8395\,
            lcout => \U712_REG_SM.N_196\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI347S_1_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8394\,
            in1 => \N__8303\,
            in2 => \_gnd_net_\,
            in3 => \N__8447\,
            lcout => \U712_REG_SM.N_383\,
            ltout => \U712_REG_SM.N_383_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_0_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__8479\,
            in1 => \_gnd_net_\,
            in2 => \N__5892\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.N_281\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__8125\,
            in1 => \N__5882\,
            in2 => \_gnd_net_\,
            in3 => \N__7145\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010111"
        )
    port map (
            in0 => \N__7377\,
            in1 => \N__7322\,
            in2 => \N__5823\,
            in3 => \N__7449\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_321_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__8614\,
            in1 => \N__8128\,
            in2 => \N__5826\,
            in3 => \N__7378\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10692\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7321\,
            in2 => \_gnd_net_\,
            in3 => \N__5819\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_156_i_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__7259\,
            in1 => \N__6060\,
            in2 => \N__5751\,
            in3 => \N__11209\,
            lcout => \N_156_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_126_i_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__5784\,
            in1 => \N__5747\,
            in2 => \N__11211\,
            in3 => \N__7743\,
            lcout => \N_126_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__8848\,
            in1 => \N__9563\,
            in2 => \_gnd_net_\,
            in3 => \N__9482\,
            lcout => \U712_BYTE_ENABLE.N_315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__9712\,
            in1 => \N__9632\,
            in2 => \N__9564\,
            in3 => \N__8847\,
            lcout => \U712_BYTE_ENABLE.N_319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__11334\,
            in1 => \N__6734\,
            in2 => \_gnd_net_\,
            in3 => \N__8480\,
            lcout => \U712_REG_SM.N_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_2_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__8482\,
            in1 => \N__6052\,
            in2 => \N__8306\,
            in3 => \N__8397\,
            lcout => \U712_REG_SM.un1_STATE_COUNT_4_i_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_1_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__6053\,
            in1 => \N__6735\,
            in2 => \N__8307\,
            in3 => \N__8481\,
            lcout => \U712_REG_SM.N_274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101100000001"
        )
    port map (
            in0 => \N__6018\,
            in1 => \N__6012\,
            in2 => \N__6006\,
            in3 => \N__9743\,
            lcout => \DS_ENm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10700\,
            ce => 'H',
            sr => \N__9942\
        );

    \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__11148\,
            in1 => \N__11266\,
            in2 => \_gnd_net_\,
            in3 => \N__11205\,
            lcout => \DMA_LATCH_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9333\,
            in1 => \N__5964\,
            in2 => \_gnd_net_\,
            in3 => \N__5949\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5931\,
            in1 => \N__5916\,
            in2 => \_gnd_net_\,
            in3 => \N__9332\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111001010"
        )
    port map (
            in0 => \N__7058\,
            in1 => \N__6699\,
            in2 => \N__6500\,
            in3 => \N__6681\,
            lcout => \U712_CHIP_RAM.N_237\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__6744\,
            in1 => \N__6870\,
            in2 => \N__6600\,
            in3 => \N__6185\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110100000001"
        )
    port map (
            in0 => \N__6528\,
            in1 => \N__6824\,
            in2 => \N__6522\,
            in3 => \N__9360\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10668\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__6364\,
            in1 => \N__6519\,
            in2 => \N__6510\,
            in3 => \N__6496\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6408\,
            in1 => \N__6387\,
            in2 => \_gnd_net_\,
            in3 => \N__9358\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9359\,
            in1 => \N__8826\,
            in2 => \N__6372\,
            in3 => \N__8913\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_1_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__7180\,
            in1 => \N__6363\,
            in2 => \N__7064\,
            in3 => \N__11123\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIE24B8_4_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__8071\,
            in1 => \N__6248\,
            in2 => \N__6186\,
            in3 => \N__6170\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_0\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8070\,
            in2 => \N__6063\,
            in3 => \N__7212\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6823\,
            in2 => \N__7185\,
            in3 => \N__9030\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10673\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7651\,
            in2 => \_gnd_net_\,
            in3 => \N__7593\,
            lcout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100110001"
        )
    port map (
            in0 => \N__7592\,
            in1 => \N__9029\,
            in2 => \N__7662\,
            in3 => \N__9320\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIMEP34_1_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100000000000"
        )
    port map (
            in0 => \N__7181\,
            in1 => \N__8072\,
            in2 => \N__7065\,
            in3 => \N__6947\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_293_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNILH2MF_1_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__6887\,
            in1 => \N__6868\,
            in2 => \N__6834\,
            in3 => \N__6831\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000001110"
        )
    port map (
            in0 => \N__6804\,
            in1 => \N__6798\,
            in2 => \N__6792\,
            in3 => \N__7594\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10673\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8073\,
            in2 => \_gnd_net_\,
            in3 => \N__6786\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__6724\,
            in1 => \N__8396\,
            in2 => \_gnd_net_\,
            in3 => \N__8305\,
            lcout => \U712_REG_SM.N_235\,
            ltout => \U712_REG_SM.N_235_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11345\,
            in2 => \N__7497\,
            in3 => \N__8341\,
            lcout => \U712_REG_SM.REG_TACK_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__7647\,
            in1 => \N__7591\,
            in2 => \N__9037\,
            in3 => \N__9361\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010111000"
        )
    port map (
            in0 => \N__7482\,
            in1 => \N__8074\,
            in2 => \N__9829\,
            in3 => \N__7476\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001000100010"
        )
    port map (
            in0 => \N__7470\,
            in1 => \N__7450\,
            in2 => \N__7428\,
            in3 => \N__7408\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10683\,
            ce => 'H',
            sr => \N__9943\
        );

    \U712_REG_SM.REG_TACK_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__7352\,
            in1 => \N__7332\,
            in2 => \N__7326\,
            in3 => \N__8223\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10683\,
            ce => 'H',
            sr => \N__9943\
        );

    \U712_REG_SM.C3_SYNC_1_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7269\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10683\,
            ce => 'H',
            sr => \N__9943\
        );

    \U712_REG_SM.C3_SYNC_0_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7292\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10683\,
            ce => 'H',
            sr => \N__9943\
        );

    \U712_BYTE_ENABLE.LMBE_i_o2_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111000111011"
        )
    port map (
            in0 => \N__9713\,
            in1 => \N__9558\,
            in2 => \N__9650\,
            in3 => \N__9483\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_220_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_151_i_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111011101"
        )
    port map (
            in0 => \N__7263\,
            in1 => \N__11279\,
            in2 => \N__7242\,
            in3 => \N__8849\,
            lcout => \N_151_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__9641\,
            in1 => \N__9714\,
            in2 => \N__8853\,
            in3 => \N__9559\,
            lcout => \U712_BYTE_ENABLE.N_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UUBE_0_a2_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__9593\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9702\,
            lcout => \U712_BYTE_ENABLE.UUBE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8095\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WEn_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7613\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10658\,
            ce => 'H',
            sr => \N__9986\
        );

    \U712_CHIP_RAM.RASn_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7677\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10658\,
            ce => 'H',
            sr => \N__9986\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__7676\,
            in1 => \N__9392\,
            in2 => \N__9051\,
            in3 => \N__7614\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10660\,
            ce => \N__10560\,
            sr => \N__9980\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__7964\,
            in1 => \N__7503\,
            in2 => \N__8836\,
            in3 => \N__7545\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10660\,
            ce => \N__10560\,
            sr => \N__9980\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9213\,
            in1 => \N__10315\,
            in2 => \_gnd_net_\,
            in3 => \N__9144\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10098\,
            ce => \N__10059\,
            sr => \N__9971\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7905\,
            in1 => \N__7887\,
            in2 => \_gnd_net_\,
            in3 => \N__9370\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7857\,
            in2 => \_gnd_net_\,
            in3 => \N__8000\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8131\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8001\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10667\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7851\,
            in1 => \N__7833\,
            in2 => \_gnd_net_\,
            in3 => \N__9342\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__8794\,
            in1 => \N__7812\,
            in2 => \N__9380\,
            in3 => \N__8670\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8792\,
            in2 => \_gnd_net_\,
            in3 => \N__9343\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__8793\,
            in1 => \N__7806\,
            in2 => \N__9379\,
            in3 => \N__8646\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__10850\,
            in1 => \N__8865\,
            in2 => \N__10798\,
            in3 => \N__7800\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10676\,
            ce => \N__10543\,
            sr => \N__9952\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7779\,
            in1 => \N__7761\,
            in2 => \_gnd_net_\,
            in3 => \N__9356\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9357\,
            in1 => \N__8825\,
            in2 => \N__8499\,
            in3 => \N__8625\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10013\,
            in2 => \_gnd_net_\,
            in3 => \N__8496\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011110101111"
        )
    port map (
            in0 => \N__8490\,
            in1 => \N__8399\,
            in2 => \N__8351\,
            in3 => \N__8451\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_236_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000100"
        )
    port map (
            in0 => \N__8400\,
            in1 => \N__8130\,
            in2 => \N__8421\,
            in3 => \N__8309\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10688\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__8398\,
            in1 => \N__8342\,
            in2 => \_gnd_net_\,
            in3 => \N__8308\,
            lcout => \U712_REG_SM.N_273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__11210\,
            in1 => \N__8129\,
            in2 => \_gnd_net_\,
            in3 => \N__11272\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10688\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__7989\,
            in1 => \N__8824\,
            in2 => \N__7968\,
            in3 => \N__9156\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10661\,
            ce => \N__10555\,
            sr => \N__9987\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10254\,
            in1 => \N__9208\,
            in2 => \_gnd_net_\,
            in3 => \N__9140\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__10063\,
            sr => \N__9981\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__8822\,
            in1 => \N__8664\,
            in2 => \N__7914\,
            in3 => \N__9400\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9399\,
            in1 => \N__8823\,
            in2 => \N__8685\,
            in3 => \N__8676\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9139\,
            in1 => \N__10253\,
            in2 => \_gnd_net_\,
            in3 => \N__10418\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__10056\,
            sr => \N__9968\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10252\,
            in1 => \N__10464\,
            in2 => \_gnd_net_\,
            in3 => \N__10929\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__10056\,
            sr => \N__9968\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10372\,
            in1 => \N__10251\,
            in2 => \_gnd_net_\,
            in3 => \N__8901\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__10054\,
            sr => \N__9960\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8900\,
            in1 => \N__10250\,
            in2 => \_gnd_net_\,
            in3 => \N__11027\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__10054\,
            sr => \N__9960\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11028\,
            in1 => \N__10310\,
            in2 => \_gnd_net_\,
            in3 => \N__8899\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10096\,
            ce => \N__10057\,
            sr => \N__9953\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10149\,
            in1 => \N__10309\,
            in2 => \_gnd_net_\,
            in3 => \N__10923\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            ce => \N__10060\,
            sr => \N__9946\
        );

    \pll_RNI8MQ3_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8618\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UMBE_0_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111000000"
        )
    port map (
            in0 => \N__9648\,
            in1 => \N__9698\,
            in2 => \N__9528\,
            in3 => \N__9465\,
            lcout => \UMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UUBE_i_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9649\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9699\,
            lcout => \U712_BYTE_ENABLE_UUBE_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CRCSn_LC_15_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9050\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10659\,
            ce => 'H',
            sr => \N__9993\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__10877\,
            in1 => \N__9102\,
            in2 => \N__10827\,
            in3 => \N__8985\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10672\,
            ce => \N__10566\,
            sr => \N__9988\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__10887\,
            in1 => \N__10876\,
            in2 => \N__10826\,
            in3 => \N__8958\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10677\,
            ce => \N__10561\,
            sr => \N__9982\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10311\,
            in1 => \N__10417\,
            in2 => \_gnd_net_\,
            in3 => \N__10463\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__10061\,
            sr => \N__9972\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10986\,
            in1 => \N__10300\,
            in2 => \_gnd_net_\,
            in3 => \N__11023\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10055\,
            sr => \N__9969\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10148\,
            in1 => \N__10308\,
            in2 => \_gnd_net_\,
            in3 => \N__10374\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__10062\,
            sr => \N__9961\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10307\,
            in1 => \N__10373\,
            in2 => \_gnd_net_\,
            in3 => \N__8890\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10097\,
            ce => \N__10064\,
            sr => \N__9954\
        );

    \U712_BYTE_ENABLE.un1_UDSn_i_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__9642\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9755\,
            lcout => \U712_BYTE_ENABLE_un1_UDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_0_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100101010"
        )
    port map (
            in0 => \N__9479\,
            in1 => \N__9700\,
            in2 => \N__9651\,
            in3 => \N__9542\,
            lcout => \LLBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100101111"
        )
    port map (
            in0 => \N__9481\,
            in1 => \N__9647\,
            in2 => \N__9759\,
            in3 => \N__9546\,
            lcout => \N_119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_220_i_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111010000"
        )
    port map (
            in0 => \N__9701\,
            in1 => \N__9646\,
            in2 => \N__9557\,
            in3 => \N__9480\,
            lcout => \N_220_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CASn_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9401\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10662\,
            ce => 'H',
            sr => \N__9994\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9225\,
            in1 => \N__10299\,
            in2 => \_gnd_net_\,
            in3 => \N__9207\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10095\,
            ce => \N__10068\,
            sr => \N__9992\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9129\,
            in1 => \N__10298\,
            in2 => \_gnd_net_\,
            in3 => \N__10419\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10092\,
            ce => \N__10065\,
            sr => \N__9989\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__10866\,
            in1 => \N__10380\,
            in2 => \N__10821\,
            in3 => \N__9096\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10689\,
            ce => \N__10554\,
            sr => \N__9983\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__10865\,
            in1 => \N__10962\,
            in2 => \N__10820\,
            in3 => \N__9072\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10689\,
            ce => \N__10554\,
            sr => \N__9983\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10287\,
            in1 => \N__11022\,
            in2 => \_gnd_net_\,
            in3 => \N__10982\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10093\,
            ce => \N__10058\,
            sr => \N__9973\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10925\,
            in1 => \N__10455\,
            in2 => \_gnd_net_\,
            in3 => \N__10288\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10093\,
            ce => \N__10058\,
            sr => \N__9973\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10146\,
            in1 => \N__10289\,
            in2 => \_gnd_net_\,
            in3 => \N__10924\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10093\,
            ce => \N__10058\,
            sr => \N__9973\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__10878\,
            in1 => \N__10104\,
            in2 => \N__10825\,
            in3 => \N__10737\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10697\,
            ce => \N__10547\,
            sr => \N__9970\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10456\,
            in1 => \N__10297\,
            in2 => \_gnd_net_\,
            in3 => \N__10413\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10091\,
            ce => \N__10066\,
            sr => \N__9990\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10362\,
            in1 => \N__10296\,
            in2 => \_gnd_net_\,
            in3 => \N__10147\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10094\,
            ce => \N__10067\,
            sr => \N__9974\
        );

    \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__11180\,
            in1 => \N__9843\,
            in2 => \_gnd_net_\,
            in3 => \N__11248\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_0_m2_LC_24_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001111111"
        )
    port map (
            in0 => \N__11349\,
            in1 => \N__11247\,
            in2 => \N__11190\,
            in3 => \N__11147\,
            lcout => \N_238\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Feb 19 2025 16:48:39

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    CMA : out std_logic_vector(10 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    A : in std_logic_vector(20 downto 0);
    RAMENn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    DBRn : in std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__11973\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10434\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \N_1062_i\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.N_348\ : std_logic;
signal \DBRn_c_i_cascade_\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_START_RNITO6SZ0Z1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_319\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_cascade_\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A20C_net\ : std_logic;
signal \U712_REG_SM.C1_SYNC_RNIAS4F1Z0Z_1\ : std_logic;
signal \U712_REG_SM.N_346_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_srsts_i_i_0_o2_0_1_3_cascade_\ : std_logic;
signal \U712_REG_SM.N_342\ : std_logic;
signal \U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0_0\ : std_logic;
signal \U712_REG_SM.N_106\ : std_logic;
signal \U712_REG_SM.N_379\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \REGENn_c\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0\ : std_logic;
signal \U712_CHIP_RAM.N_409\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_489_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_361_cascade_\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z20\ : std_logic;
signal \U712_CHIP_RAM.N_416_cascade_\ : std_logic;
signal \U712_CHIP_RAM.BANK0_RNOZ0Z_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_i_i_0\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_410_cascade_\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_RNI4BRHZ0Z_3\ : std_logic;
signal \U712_REG_SM.N_400\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_12_0\ : std_logic;
signal \LATCH_CLK_c\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U712_CHIP_RAM.N_489\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_304\ : std_logic;
signal \U712_CHIP_RAM.N_62_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_452\ : std_logic;
signal \U712_CHIP_RAM.N_452_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_11_cascade_\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.N_288_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_372_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_366_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_15_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_0_0\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_448\ : std_logic;
signal \U712_CHIP_RAM.N_345_cascade_\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_i_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_11_2\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.N_316_i_0_en\ : std_logic;
signal \U712_CYCLE_TERM.N_316_i_0_en_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_282_i\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.N_371_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_0_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_371_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_288\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_329\ : std_logic;
signal \U712_CHIP_RAM.N_414_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_86\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_373\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER15\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_286_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_486\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a2_1\ : std_logic;
signal \U712_CHIP_RAM.N_287_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_436\ : std_logic;
signal \U712_CHIP_RAM.N_283\ : std_logic;
signal \U712_CHIP_RAM.N_347\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_i_0_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_129_i_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_286\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C1_SYNC_RNIAS4F1_0Z0Z_1_cascade_\ : std_logic;
signal \U712_REG_SM.ASn_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a2_0_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.C1_SYNC_RNIAS4F1_0Z0Z_1\ : std_logic;
signal \U712_REG_SM.N_104\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNO_6Z0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1\ : std_logic;
signal \U712_CHIP_RAM.N_287\ : std_logic;
signal \U712_CHIP_RAM.N_388\ : std_logic;
signal \U712_CHIP_RAM.N_370\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUUBEn_i_0_aZ0Z2\ : std_logic;
signal \N_38_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_426_cascade_\ : std_logic;
signal \N_47_i\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLMBEn_i_0_aZ0Z2\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \N_46_i\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2Z0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_431\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2Z0Z_0_cascade_\ : std_logic;
signal \N_45_i\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2Z0Z_0\ : std_logic;
signal \RnW_c\ : std_logic;
signal \N_344\ : std_logic;
signal \DMA_LATCH_EN_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \A_c_8\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.N_62\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.N_434_i\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_201_i_i_a2_3_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \WRITE_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.N_306_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.un3_DMA_CYCLE_START\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8_cascade_\ : std_logic;
signal \A_c_14\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.N_463_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRTZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \A_c_3\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_0\ : std_logic;
signal \A_c_13\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \RASn_c\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \N_357_i\ : std_logic;
signal \N_42\ : std_logic;
signal \N_231\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \N_358_i\ : std_logic;
signal \DS_ENm\ : std_logic;
signal \N_40\ : std_logic;
signal \A_c_1\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \LLBEn_c\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \RAMENn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    RAMENn <= \RAMENn_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__4004\,
            RESETB => \N__5051\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11973\,
            DIN => \N__11972\,
            DOUT => \N__11971\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11973\,
            PADOUT => \N__11972\,
            PADIN => \N__11971\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6233\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11964\,
            DIN => \N__11963\,
            DOUT => \N__11962\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11964\,
            PADOUT => \N__11963\,
            PADIN => \N__11962\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11955\,
            DIN => \N__11954\,
            DOUT => \N__11953\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11955\,
            PADOUT => \N__11954\,
            PADIN => \N__11953\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8921\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11946\,
            DIN => \N__11945\,
            DOUT => \N__11944\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11946\,
            PADOUT => \N__11945\,
            PADIN => \N__11944\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6500\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11937\,
            DIN => \N__11936\,
            DOUT => \N__11935\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11937\,
            PADOUT => \N__11936\,
            PADIN => \N__11935\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11928\,
            DIN => \N__11927\,
            DOUT => \N__11926\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11928\,
            PADOUT => \N__11927\,
            PADIN => \N__11926\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11919\,
            DIN => \N__11918\,
            DOUT => \N__11917\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11919\,
            PADOUT => \N__11918\,
            PADIN => \N__11917\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11910\,
            DIN => \N__11909\,
            DOUT => \N__11908\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11910\,
            PADOUT => \N__11909\,
            PADIN => \N__11908\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11901\,
            DIN => \N__11900\,
            DOUT => \N__11899\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11901\,
            PADOUT => \N__11900\,
            PADIN => \N__11899\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11892\,
            DIN => \N__11891\,
            DOUT => \N__11890\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11892\,
            PADOUT => \N__11891\,
            PADIN => \N__11890\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11883\,
            DIN => \N__11882\,
            DOUT => \N__11881\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11883\,
            PADOUT => \N__11882\,
            PADIN => \N__11881\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6446\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11874\,
            DIN => \N__11873\,
            DOUT => \N__11872\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11874\,
            PADOUT => \N__11873\,
            PADIN => \N__11872\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10664\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11865\,
            DIN => \N__11864\,
            DOUT => \N__11863\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11865\,
            PADOUT => \N__11864\,
            PADIN => \N__11863\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11856\,
            DIN => \N__11855\,
            DOUT => \N__11854\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11856\,
            PADOUT => \N__11855\,
            PADIN => \N__11854\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11847\,
            DIN => \N__11846\,
            DOUT => \N__11845\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11847\,
            PADOUT => \N__11846\,
            PADIN => \N__11845\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11838\,
            DIN => \N__11837\,
            DOUT => \N__11836\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11838\,
            PADOUT => \N__11837\,
            PADIN => \N__11836\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4250\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11829\,
            DIN => \N__11828\,
            DOUT => \N__11827\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11829\,
            PADOUT => \N__11828\,
            PADIN => \N__11827\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11820\,
            DIN => \N__11819\,
            DOUT => \N__11818\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11820\,
            PADOUT => \N__11819\,
            PADIN => \N__11818\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11811\,
            DIN => \N__11810\,
            DOUT => \N__11809\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11811\,
            PADOUT => \N__11810\,
            PADIN => \N__11809\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8894\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11802\,
            DIN => \N__11801\,
            DOUT => \N__11800\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11802\,
            PADOUT => \N__11801\,
            PADIN => \N__11800\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11793\,
            DIN => \N__11792\,
            DOUT => \N__11791\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11793\,
            PADOUT => \N__11792\,
            PADIN => \N__11791\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8057\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11784\,
            DIN => \N__11783\,
            DOUT => \N__11782\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11784\,
            PADOUT => \N__11783\,
            PADIN => \N__11782\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11775\,
            DIN => \N__11774\,
            DOUT => \N__11773\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11775\,
            PADOUT => \N__11774\,
            PADIN => \N__11773\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9980\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11766\,
            DIN => \N__11765\,
            DOUT => \N__11764\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11766\,
            PADOUT => \N__11765\,
            PADIN => \N__11764\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11757\,
            DIN => \N__11756\,
            DOUT => \N__11755\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11757\,
            PADOUT => \N__11756\,
            PADIN => \N__11755\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11748\,
            DIN => \N__11747\,
            DOUT => \N__11746\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11748\,
            PADOUT => \N__11747\,
            PADIN => \N__11746\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11739\,
            DIN => \N__11738\,
            DOUT => \N__11737\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11739\,
            PADOUT => \N__11738\,
            PADIN => \N__11737\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11730\,
            DIN => \N__11729\,
            DOUT => \N__11728\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11730\,
            PADOUT => \N__11729\,
            PADIN => \N__11728\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11721\,
            DIN => \N__11720\,
            DOUT => \N__11719\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11721\,
            PADOUT => \N__11720\,
            PADIN => \N__11719\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6476\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11712\,
            DIN => \N__11711\,
            DOUT => \N__11710\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11712\,
            PADOUT => \N__11711\,
            PADIN => \N__11710\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11703\,
            DIN => \N__11702\,
            DOUT => \N__11701\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11703\,
            PADOUT => \N__11702\,
            PADIN => \N__11701\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11694\,
            DIN => \N__11693\,
            DOUT => \N__11692\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11694\,
            PADOUT => \N__11693\,
            PADIN => \N__11692\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11685\,
            DIN => \N__11684\,
            DOUT => \N__11683\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11685\,
            PADOUT => \N__11684\,
            PADIN => \N__11683\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11676\,
            DIN => \N__11675\,
            DOUT => \N__11674\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11676\,
            PADOUT => \N__11675\,
            PADIN => \N__11674\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11667\,
            DIN => \N__11666\,
            DOUT => \N__11665\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11667\,
            PADOUT => \N__11666\,
            PADIN => \N__11665\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9842\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11658\,
            DIN => \N__11657\,
            DOUT => \N__11656\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11658\,
            PADOUT => \N__11657\,
            PADIN => \N__11656\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11649\,
            DIN => \N__11648\,
            DOUT => \N__11647\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11649\,
            PADOUT => \N__11648\,
            PADIN => \N__11647\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4568\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11640\,
            DIN => \N__11639\,
            DOUT => \N__11638\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11640\,
            PADOUT => \N__11639\,
            PADIN => \N__11638\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8440\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11631\,
            DIN => \N__11630\,
            DOUT => \N__11629\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11631\,
            PADOUT => \N__11630\,
            PADIN => \N__11629\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4055\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11622\,
            DIN => \N__11621\,
            DOUT => \N__11620\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11622\,
            PADOUT => \N__11621\,
            PADIN => \N__11620\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11613\,
            DIN => \N__11612\,
            DOUT => \N__11611\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11613\,
            PADOUT => \N__11612\,
            PADIN => \N__11611\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4232\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11604\,
            DIN => \N__11603\,
            DOUT => \N__11602\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11604\,
            PADOUT => \N__11603\,
            PADIN => \N__11602\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8024\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11595\,
            DIN => \N__11594\,
            DOUT => \N__11593\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11595\,
            PADOUT => \N__11594\,
            PADIN => \N__11593\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11586\,
            DIN => \N__11585\,
            DOUT => \N__11584\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11586\,
            PADOUT => \N__11585\,
            PADIN => \N__11584\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11577\,
            DIN => \N__11576\,
            DOUT => \N__11575\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11577\,
            PADOUT => \N__11576\,
            PADIN => \N__11575\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11568\,
            DIN => \N__11567\,
            DOUT => \N__11566\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11568\,
            PADOUT => \N__11567\,
            PADIN => \N__11566\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11559\,
            DIN => \N__11558\,
            DOUT => \N__11557\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11559\,
            PADOUT => \N__11558\,
            PADIN => \N__11557\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11550\,
            DIN => \N__11549\,
            DOUT => \N__11548\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11550\,
            PADOUT => \N__11549\,
            PADIN => \N__11548\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8834\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11541\,
            DIN => \N__11540\,
            DOUT => \N__11539\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11541\,
            PADOUT => \N__11540\,
            PADIN => \N__11539\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11532\,
            DIN => \N__11531\,
            DOUT => \N__11530\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11532\,
            PADOUT => \N__11531\,
            PADIN => \N__11530\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8415\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11523\,
            DIN => \N__11522\,
            DOUT => \N__11521\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11523\,
            PADOUT => \N__11522\,
            PADIN => \N__11521\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8690\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11514\,
            DIN => \N__11513\,
            DOUT => \N__11512\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11514\,
            PADOUT => \N__11513\,
            PADIN => \N__11512\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8078\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11505\,
            DIN => \N__11504\,
            DOUT => \N__11503\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11505\,
            PADOUT => \N__11504\,
            PADIN => \N__11503\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6587\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11496\,
            DIN => \N__11495\,
            DOUT => \N__11494\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11496\,
            PADOUT => \N__11495\,
            PADIN => \N__11494\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8648\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11487\,
            DIN => \N__11486\,
            DOUT => \N__11485\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11487\,
            PADOUT => \N__11486\,
            PADIN => \N__11485\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4295\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11478\,
            DIN => \N__11477\,
            DOUT => \N__11476\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11478\,
            PADOUT => \N__11477\,
            PADIN => \N__11476\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11469\,
            DIN => \N__11468\,
            DOUT => \N__11467\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11469\,
            PADOUT => \N__11468\,
            PADIN => \N__11467\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11460\,
            DIN => \N__11459\,
            DOUT => \N__11458\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11460\,
            PADOUT => \N__11459\,
            PADIN => \N__11458\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6182\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11451\,
            DIN => \N__11450\,
            DOUT => \N__11449\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11451\,
            PADOUT => \N__11450\,
            PADIN => \N__11449\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9917\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11442\,
            DIN => \N__11441\,
            DOUT => \N__11440\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11442\,
            PADOUT => \N__11441\,
            PADIN => \N__11440\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4712\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11433\,
            DIN => \N__11432\,
            DOUT => \N__11431\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11433\,
            PADOUT => \N__11432\,
            PADIN => \N__11431\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6266\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11424\,
            DIN => \N__11423\,
            DOUT => \N__11422\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11424\,
            PADOUT => \N__11423\,
            PADIN => \N__11422\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11415\,
            DIN => \N__11414\,
            DOUT => \N__11413\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11415\,
            PADOUT => \N__11414\,
            PADIN => \N__11413\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11406\,
            DIN => \N__11405\,
            DOUT => \N__11404\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11406\,
            PADOUT => \N__11405\,
            PADIN => \N__11404\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11397\,
            DIN => \N__11396\,
            DOUT => \N__11395\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11397\,
            PADOUT => \N__11396\,
            PADIN => \N__11395\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11388\,
            DIN => \N__11387\,
            DOUT => \N__11386\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11388\,
            PADOUT => \N__11387\,
            PADIN => \N__11386\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9155\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11379\,
            DIN => \N__11378\,
            DOUT => \N__11377\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11379\,
            PADOUT => \N__11378\,
            PADIN => \N__11377\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10391\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11370\,
            DIN => \N__11369\,
            DOUT => \N__11368\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11370\,
            PADOUT => \N__11369\,
            PADIN => \N__11368\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11361\,
            DIN => \N__11360\,
            DOUT => \N__11359\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11361\,
            PADOUT => \N__11360\,
            PADIN => \N__11359\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6293\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11352\,
            DIN => \N__11351\,
            DOUT => \N__11350\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11352\,
            PADOUT => \N__11351\,
            PADIN => \N__11350\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4067\,
            DIN0 => OPEN,
            DOUT0 => \N__4889\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11343\,
            DIN => \N__11342\,
            DOUT => \N__11341\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11343\,
            PADOUT => \N__11342\,
            PADIN => \N__11341\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7676\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11334\,
            DIN => \N__11333\,
            DOUT => \N__11332\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11334\,
            PADOUT => \N__11333\,
            PADIN => \N__11332\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11325\,
            DIN => \N__11324\,
            DOUT => \N__11323\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11325\,
            PADOUT => \N__11324\,
            PADIN => \N__11323\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11316\,
            DIN => \N__11315\,
            DOUT => \N__11314\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11316\,
            PADOUT => \N__11315\,
            PADIN => \N__11314\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8582\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11307\,
            DIN => \N__11306\,
            DOUT => \N__11305\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11307\,
            PADOUT => \N__11306\,
            PADIN => \N__11305\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11298\,
            DIN => \N__11297\,
            DOUT => \N__11296\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11298\,
            PADOUT => \N__11297\,
            PADIN => \N__11296\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11289\,
            DIN => \N__11288\,
            DOUT => \N__11287\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11289\,
            PADOUT => \N__11288\,
            PADIN => \N__11287\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11280\,
            DIN => \N__11279\,
            DOUT => \N__11278\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11280\,
            PADOUT => \N__11279\,
            PADIN => \N__11278\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11271\,
            DIN => \N__11270\,
            DOUT => \N__11269\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11271\,
            PADOUT => \N__11270\,
            PADIN => \N__11269\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8804\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11262\,
            DIN => \N__11261\,
            DOUT => \N__11260\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11262\,
            PADOUT => \N__11261\,
            PADIN => \N__11260\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10649\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11253\,
            DIN => \N__11252\,
            DOUT => \N__11251\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11253\,
            PADOUT => \N__11252\,
            PADIN => \N__11251\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10631\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11244\,
            DIN => \N__11243\,
            DOUT => \N__11242\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11244\,
            PADOUT => \N__11243\,
            PADIN => \N__11242\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4958\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11235\,
            DIN => \N__11234\,
            DOUT => \N__11233\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11235\,
            PADOUT => \N__11234\,
            PADIN => \N__11233\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11226\,
            DIN => \N__11225\,
            DOUT => \N__11224\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11226\,
            PADOUT => \N__11225\,
            PADIN => \N__11224\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11217\,
            DIN => \N__11216\,
            DOUT => \N__11215\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11217\,
            PADOUT => \N__11216\,
            PADIN => \N__11215\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6692\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11208\,
            DIN => \N__11207\,
            DOUT => \N__11206\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11208\,
            PADOUT => \N__11207\,
            PADIN => \N__11206\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11199\,
            DIN => \N__11198\,
            DOUT => \N__11197\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11199\,
            PADOUT => \N__11198\,
            PADIN => \N__11197\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11190\,
            DIN => \N__11189\,
            DOUT => \N__11188\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11190\,
            PADOUT => \N__11189\,
            PADIN => \N__11188\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4664\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11181\,
            DIN => \N__11180\,
            DOUT => \N__11179\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11181\,
            PADOUT => \N__11180\,
            PADIN => \N__11179\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10346\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11172\,
            DIN => \N__11171\,
            DOUT => \N__11170\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11172\,
            PADOUT => \N__11171\,
            PADIN => \N__11170\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8441\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2732\ : InMux
    port map (
            O => \N__11153\,
            I => \N__11149\
        );

    \I__2731\ : InMux
    port map (
            O => \N__11152\,
            I => \N__11146\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__11149\,
            I => \N__11142\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__11146\,
            I => \N__11139\
        );

    \I__2728\ : InMux
    port map (
            O => \N__11145\,
            I => \N__11136\
        );

    \I__2727\ : Span4Mux_v
    port map (
            O => \N__11142\,
            I => \N__11133\
        );

    \I__2726\ : Span4Mux_h
    port map (
            O => \N__11139\,
            I => \N__11128\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__11136\,
            I => \N__11128\
        );

    \I__2724\ : Span4Mux_v
    port map (
            O => \N__11133\,
            I => \N__11124\
        );

    \I__2723\ : Span4Mux_v
    port map (
            O => \N__11128\,
            I => \N__11121\
        );

    \I__2722\ : InMux
    port map (
            O => \N__11127\,
            I => \N__11118\
        );

    \I__2721\ : Sp12to4
    port map (
            O => \N__11124\,
            I => \N__11115\
        );

    \I__2720\ : Sp12to4
    port map (
            O => \N__11121\,
            I => \N__11112\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__11118\,
            I => \N__11109\
        );

    \I__2718\ : Span12Mux_h
    port map (
            O => \N__11115\,
            I => \N__11106\
        );

    \I__2717\ : Span12Mux_h
    port map (
            O => \N__11112\,
            I => \N__11103\
        );

    \I__2716\ : Span12Mux_v
    port map (
            O => \N__11109\,
            I => \N__11100\
        );

    \I__2715\ : Span12Mux_v
    port map (
            O => \N__11106\,
            I => \N__11097\
        );

    \I__2714\ : Span12Mux_v
    port map (
            O => \N__11103\,
            I => \N__11094\
        );

    \I__2713\ : Span12Mux_v
    port map (
            O => \N__11100\,
            I => \N__11091\
        );

    \I__2712\ : Odrv12
    port map (
            O => \N__11097\,
            I => \DRA_c_9\
        );

    \I__2711\ : Odrv12
    port map (
            O => \N__11094\,
            I => \DRA_c_9\
        );

    \I__2710\ : Odrv12
    port map (
            O => \N__11091\,
            I => \DRA_c_9\
        );

    \I__2709\ : InMux
    port map (
            O => \N__11084\,
            I => \N__11081\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__11081\,
            I => \N__11078\
        );

    \I__2707\ : Odrv12
    port map (
            O => \N__11078\,
            I => \RAS0n_c\
        );

    \I__2706\ : CascadeMux
    port map (
            O => \N__11075\,
            I => \N__11072\
        );

    \I__2705\ : InMux
    port map (
            O => \N__11072\,
            I => \N__11066\
        );

    \I__2704\ : InMux
    port map (
            O => \N__11071\,
            I => \N__11063\
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__11070\,
            I => \N__11056\
        );

    \I__2702\ : CascadeMux
    port map (
            O => \N__11069\,
            I => \N__11050\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__11066\,
            I => \N__11043\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__11063\,
            I => \N__11043\
        );

    \I__2699\ : InMux
    port map (
            O => \N__11062\,
            I => \N__11038\
        );

    \I__2698\ : InMux
    port map (
            O => \N__11061\,
            I => \N__11038\
        );

    \I__2697\ : InMux
    port map (
            O => \N__11060\,
            I => \N__11033\
        );

    \I__2696\ : InMux
    port map (
            O => \N__11059\,
            I => \N__11033\
        );

    \I__2695\ : InMux
    port map (
            O => \N__11056\,
            I => \N__11025\
        );

    \I__2694\ : InMux
    port map (
            O => \N__11055\,
            I => \N__11025\
        );

    \I__2693\ : InMux
    port map (
            O => \N__11054\,
            I => \N__11025\
        );

    \I__2692\ : InMux
    port map (
            O => \N__11053\,
            I => \N__11022\
        );

    \I__2691\ : InMux
    port map (
            O => \N__11050\,
            I => \N__11017\
        );

    \I__2690\ : InMux
    port map (
            O => \N__11049\,
            I => \N__11017\
        );

    \I__2689\ : InMux
    port map (
            O => \N__11048\,
            I => \N__11013\
        );

    \I__2688\ : Span4Mux_h
    port map (
            O => \N__11043\,
            I => \N__11007\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__11038\,
            I => \N__11007\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__11033\,
            I => \N__11004\
        );

    \I__2685\ : CascadeMux
    port map (
            O => \N__11032\,
            I => \N__10997\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__11025\,
            I => \N__10993\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__11022\,
            I => \N__10988\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__11017\,
            I => \N__10988\
        );

    \I__2681\ : InMux
    port map (
            O => \N__11016\,
            I => \N__10985\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__11013\,
            I => \N__10982\
        );

    \I__2679\ : InMux
    port map (
            O => \N__11012\,
            I => \N__10979\
        );

    \I__2678\ : Span4Mux_h
    port map (
            O => \N__11007\,
            I => \N__10974\
        );

    \I__2677\ : Span4Mux_v
    port map (
            O => \N__11004\,
            I => \N__10974\
        );

    \I__2676\ : InMux
    port map (
            O => \N__11003\,
            I => \N__10969\
        );

    \I__2675\ : InMux
    port map (
            O => \N__11002\,
            I => \N__10969\
        );

    \I__2674\ : InMux
    port map (
            O => \N__11001\,
            I => \N__10964\
        );

    \I__2673\ : InMux
    port map (
            O => \N__11000\,
            I => \N__10964\
        );

    \I__2672\ : InMux
    port map (
            O => \N__10997\,
            I => \N__10959\
        );

    \I__2671\ : InMux
    port map (
            O => \N__10996\,
            I => \N__10959\
        );

    \I__2670\ : Span4Mux_v
    port map (
            O => \N__10993\,
            I => \N__10952\
        );

    \I__2669\ : Span4Mux_h
    port map (
            O => \N__10988\,
            I => \N__10952\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__10985\,
            I => \N__10952\
        );

    \I__2667\ : Span4Mux_v
    port map (
            O => \N__10982\,
            I => \N__10949\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__10979\,
            I => \N__10946\
        );

    \I__2665\ : Sp12to4
    port map (
            O => \N__10974\,
            I => \N__10937\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__10969\,
            I => \N__10937\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__10964\,
            I => \N__10937\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__10959\,
            I => \N__10937\
        );

    \I__2661\ : Sp12to4
    port map (
            O => \N__10952\,
            I => \N__10934\
        );

    \I__2660\ : Span4Mux_h
    port map (
            O => \N__10949\,
            I => \N__10931\
        );

    \I__2659\ : Span12Mux_v
    port map (
            O => \N__10946\,
            I => \N__10928\
        );

    \I__2658\ : Span12Mux_h
    port map (
            O => \N__10937\,
            I => \N__10925\
        );

    \I__2657\ : Span12Mux_v
    port map (
            O => \N__10934\,
            I => \N__10922\
        );

    \I__2656\ : Sp12to4
    port map (
            O => \N__10931\,
            I => \N__10919\
        );

    \I__2655\ : Span12Mux_h
    port map (
            O => \N__10928\,
            I => \N__10914\
        );

    \I__2654\ : Span12Mux_v
    port map (
            O => \N__10925\,
            I => \N__10914\
        );

    \I__2653\ : Span12Mux_h
    port map (
            O => \N__10922\,
            I => \N__10911\
        );

    \I__2652\ : Span12Mux_v
    port map (
            O => \N__10919\,
            I => \N__10908\
        );

    \I__2651\ : Odrv12
    port map (
            O => \N__10914\,
            I => \AGNUS_REV_c\
        );

    \I__2650\ : Odrv12
    port map (
            O => \N__10911\,
            I => \AGNUS_REV_c\
        );

    \I__2649\ : Odrv12
    port map (
            O => \N__10908\,
            I => \AGNUS_REV_c\
        );

    \I__2648\ : InMux
    port map (
            O => \N__10901\,
            I => \N__10898\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__10898\,
            I => \N__10895\
        );

    \I__2646\ : Span12Mux_h
    port map (
            O => \N__10895\,
            I => \N__10892\
        );

    \I__2645\ : Odrv12
    port map (
            O => \N__10892\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2644\ : ClkMux
    port map (
            O => \N__10889\,
            I => \N__10868\
        );

    \I__2643\ : ClkMux
    port map (
            O => \N__10888\,
            I => \N__10868\
        );

    \I__2642\ : ClkMux
    port map (
            O => \N__10887\,
            I => \N__10868\
        );

    \I__2641\ : ClkMux
    port map (
            O => \N__10886\,
            I => \N__10868\
        );

    \I__2640\ : ClkMux
    port map (
            O => \N__10885\,
            I => \N__10868\
        );

    \I__2639\ : ClkMux
    port map (
            O => \N__10884\,
            I => \N__10868\
        );

    \I__2638\ : ClkMux
    port map (
            O => \N__10883\,
            I => \N__10868\
        );

    \I__2637\ : GlobalMux
    port map (
            O => \N__10868\,
            I => \N__10865\
        );

    \I__2636\ : gio2CtrlBuf
    port map (
            O => \N__10865\,
            I => \C3_c_g\
        );

    \I__2635\ : CEMux
    port map (
            O => \N__10862\,
            I => \N__10832\
        );

    \I__2634\ : CEMux
    port map (
            O => \N__10861\,
            I => \N__10832\
        );

    \I__2633\ : CEMux
    port map (
            O => \N__10860\,
            I => \N__10832\
        );

    \I__2632\ : CEMux
    port map (
            O => \N__10859\,
            I => \N__10832\
        );

    \I__2631\ : CEMux
    port map (
            O => \N__10858\,
            I => \N__10832\
        );

    \I__2630\ : CEMux
    port map (
            O => \N__10857\,
            I => \N__10832\
        );

    \I__2629\ : CEMux
    port map (
            O => \N__10856\,
            I => \N__10832\
        );

    \I__2628\ : CEMux
    port map (
            O => \N__10855\,
            I => \N__10832\
        );

    \I__2627\ : CEMux
    port map (
            O => \N__10854\,
            I => \N__10832\
        );

    \I__2626\ : CEMux
    port map (
            O => \N__10853\,
            I => \N__10832\
        );

    \I__2625\ : GlobalMux
    port map (
            O => \N__10832\,
            I => \N__10829\
        );

    \I__2624\ : gio2CtrlBuf
    port map (
            O => \N__10829\,
            I => \DBRn_c_i_0_g\
        );

    \I__2623\ : InMux
    port map (
            O => \N__10826\,
            I => \N__10817\
        );

    \I__2622\ : InMux
    port map (
            O => \N__10825\,
            I => \N__10817\
        );

    \I__2621\ : InMux
    port map (
            O => \N__10824\,
            I => \N__10814\
        );

    \I__2620\ : InMux
    port map (
            O => \N__10823\,
            I => \N__10811\
        );

    \I__2619\ : InMux
    port map (
            O => \N__10822\,
            I => \N__10808\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__10817\,
            I => \N__10797\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__10814\,
            I => \N__10790\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__10811\,
            I => \N__10772\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__10808\,
            I => \N__10763\
        );

    \I__2614\ : SRMux
    port map (
            O => \N__10807\,
            I => \N__10670\
        );

    \I__2613\ : SRMux
    port map (
            O => \N__10806\,
            I => \N__10670\
        );

    \I__2612\ : SRMux
    port map (
            O => \N__10805\,
            I => \N__10670\
        );

    \I__2611\ : SRMux
    port map (
            O => \N__10804\,
            I => \N__10670\
        );

    \I__2610\ : SRMux
    port map (
            O => \N__10803\,
            I => \N__10670\
        );

    \I__2609\ : SRMux
    port map (
            O => \N__10802\,
            I => \N__10670\
        );

    \I__2608\ : SRMux
    port map (
            O => \N__10801\,
            I => \N__10670\
        );

    \I__2607\ : SRMux
    port map (
            O => \N__10800\,
            I => \N__10670\
        );

    \I__2606\ : Glb2LocalMux
    port map (
            O => \N__10797\,
            I => \N__10670\
        );

    \I__2605\ : SRMux
    port map (
            O => \N__10796\,
            I => \N__10670\
        );

    \I__2604\ : SRMux
    port map (
            O => \N__10795\,
            I => \N__10670\
        );

    \I__2603\ : SRMux
    port map (
            O => \N__10794\,
            I => \N__10670\
        );

    \I__2602\ : SRMux
    port map (
            O => \N__10793\,
            I => \N__10670\
        );

    \I__2601\ : Glb2LocalMux
    port map (
            O => \N__10790\,
            I => \N__10670\
        );

    \I__2600\ : SRMux
    port map (
            O => \N__10789\,
            I => \N__10670\
        );

    \I__2599\ : SRMux
    port map (
            O => \N__10788\,
            I => \N__10670\
        );

    \I__2598\ : SRMux
    port map (
            O => \N__10787\,
            I => \N__10670\
        );

    \I__2597\ : SRMux
    port map (
            O => \N__10786\,
            I => \N__10670\
        );

    \I__2596\ : SRMux
    port map (
            O => \N__10785\,
            I => \N__10670\
        );

    \I__2595\ : SRMux
    port map (
            O => \N__10784\,
            I => \N__10670\
        );

    \I__2594\ : SRMux
    port map (
            O => \N__10783\,
            I => \N__10670\
        );

    \I__2593\ : SRMux
    port map (
            O => \N__10782\,
            I => \N__10670\
        );

    \I__2592\ : SRMux
    port map (
            O => \N__10781\,
            I => \N__10670\
        );

    \I__2591\ : SRMux
    port map (
            O => \N__10780\,
            I => \N__10670\
        );

    \I__2590\ : SRMux
    port map (
            O => \N__10779\,
            I => \N__10670\
        );

    \I__2589\ : SRMux
    port map (
            O => \N__10778\,
            I => \N__10670\
        );

    \I__2588\ : SRMux
    port map (
            O => \N__10777\,
            I => \N__10670\
        );

    \I__2587\ : SRMux
    port map (
            O => \N__10776\,
            I => \N__10670\
        );

    \I__2586\ : SRMux
    port map (
            O => \N__10775\,
            I => \N__10670\
        );

    \I__2585\ : Glb2LocalMux
    port map (
            O => \N__10772\,
            I => \N__10670\
        );

    \I__2584\ : SRMux
    port map (
            O => \N__10771\,
            I => \N__10670\
        );

    \I__2583\ : SRMux
    port map (
            O => \N__10770\,
            I => \N__10670\
        );

    \I__2582\ : SRMux
    port map (
            O => \N__10769\,
            I => \N__10670\
        );

    \I__2581\ : SRMux
    port map (
            O => \N__10768\,
            I => \N__10670\
        );

    \I__2580\ : SRMux
    port map (
            O => \N__10767\,
            I => \N__10670\
        );

    \I__2579\ : SRMux
    port map (
            O => \N__10766\,
            I => \N__10670\
        );

    \I__2578\ : Glb2LocalMux
    port map (
            O => \N__10763\,
            I => \N__10670\
        );

    \I__2577\ : SRMux
    port map (
            O => \N__10762\,
            I => \N__10670\
        );

    \I__2576\ : SRMux
    port map (
            O => \N__10761\,
            I => \N__10670\
        );

    \I__2575\ : SRMux
    port map (
            O => \N__10760\,
            I => \N__10670\
        );

    \I__2574\ : SRMux
    port map (
            O => \N__10759\,
            I => \N__10670\
        );

    \I__2573\ : SRMux
    port map (
            O => \N__10758\,
            I => \N__10670\
        );

    \I__2572\ : SRMux
    port map (
            O => \N__10757\,
            I => \N__10670\
        );

    \I__2571\ : GlobalMux
    port map (
            O => \N__10670\,
            I => \N__10667\
        );

    \I__2570\ : gio2CtrlBuf
    port map (
            O => \N__10667\,
            I => \RESETn_c_i_g\
        );

    \I__2569\ : IoInMux
    port map (
            O => \N__10664\,
            I => \N__10661\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__10661\,
            I => \N__10658\
        );

    \I__2567\ : Span4Mux_s0_v
    port map (
            O => \N__10658\,
            I => \N__10655\
        );

    \I__2566\ : Span4Mux_v
    port map (
            O => \N__10655\,
            I => \N__10652\
        );

    \I__2565\ : Odrv4
    port map (
            O => \N__10652\,
            I => \N_357_i\
        );

    \I__2564\ : IoInMux
    port map (
            O => \N__10649\,
            I => \N__10646\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__10646\,
            I => \N__10643\
        );

    \I__2562\ : Span4Mux_s2_v
    port map (
            O => \N__10643\,
            I => \N__10640\
        );

    \I__2561\ : Span4Mux_v
    port map (
            O => \N__10640\,
            I => \N__10637\
        );

    \I__2560\ : Sp12to4
    port map (
            O => \N__10637\,
            I => \N__10634\
        );

    \I__2559\ : Odrv12
    port map (
            O => \N__10634\,
            I => \N_42\
        );

    \I__2558\ : IoInMux
    port map (
            O => \N__10631\,
            I => \N__10628\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__10628\,
            I => \N__10625\
        );

    \I__2556\ : Span4Mux_s2_v
    port map (
            O => \N__10625\,
            I => \N__10622\
        );

    \I__2555\ : Span4Mux_h
    port map (
            O => \N__10622\,
            I => \N__10619\
        );

    \I__2554\ : Span4Mux_v
    port map (
            O => \N__10619\,
            I => \N__10616\
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__10616\,
            I => \N_231\
        );

    \I__2552\ : InMux
    port map (
            O => \N__10613\,
            I => \N__10610\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__10610\,
            I => \N__10604\
        );

    \I__2550\ : InMux
    port map (
            O => \N__10609\,
            I => \N__10599\
        );

    \I__2549\ : InMux
    port map (
            O => \N__10608\,
            I => \N__10599\
        );

    \I__2548\ : InMux
    port map (
            O => \N__10607\,
            I => \N__10596\
        );

    \I__2547\ : Span4Mux_v
    port map (
            O => \N__10604\,
            I => \N__10589\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__10599\,
            I => \N__10589\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__10596\,
            I => \N__10589\
        );

    \I__2544\ : Span4Mux_h
    port map (
            O => \N__10589\,
            I => \N__10586\
        );

    \I__2543\ : Sp12to4
    port map (
            O => \N__10586\,
            I => \N__10583\
        );

    \I__2542\ : Span12Mux_v
    port map (
            O => \N__10583\,
            I => \N__10580\
        );

    \I__2541\ : Odrv12
    port map (
            O => \N__10580\,
            I => \DRA_c_2\
        );

    \I__2540\ : InMux
    port map (
            O => \N__10577\,
            I => \N__10572\
        );

    \I__2539\ : InMux
    port map (
            O => \N__10576\,
            I => \N__10569\
        );

    \I__2538\ : InMux
    port map (
            O => \N__10575\,
            I => \N__10565\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__10572\,
            I => \N__10560\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__10569\,
            I => \N__10560\
        );

    \I__2535\ : InMux
    port map (
            O => \N__10568\,
            I => \N__10557\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__10565\,
            I => \N__10554\
        );

    \I__2533\ : Span4Mux_h
    port map (
            O => \N__10560\,
            I => \N__10551\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__10557\,
            I => \N__10548\
        );

    \I__2531\ : Sp12to4
    port map (
            O => \N__10554\,
            I => \N__10545\
        );

    \I__2530\ : Sp12to4
    port map (
            O => \N__10551\,
            I => \N__10542\
        );

    \I__2529\ : Span12Mux_h
    port map (
            O => \N__10548\,
            I => \N__10539\
        );

    \I__2528\ : Span12Mux_v
    port map (
            O => \N__10545\,
            I => \N__10536\
        );

    \I__2527\ : Span12Mux_v
    port map (
            O => \N__10542\,
            I => \N__10533\
        );

    \I__2526\ : Span12Mux_v
    port map (
            O => \N__10539\,
            I => \N__10530\
        );

    \I__2525\ : Span12Mux_h
    port map (
            O => \N__10536\,
            I => \N__10527\
        );

    \I__2524\ : Odrv12
    port map (
            O => \N__10533\,
            I => \DRA_c_1\
        );

    \I__2523\ : Odrv12
    port map (
            O => \N__10530\,
            I => \DRA_c_1\
        );

    \I__2522\ : Odrv12
    port map (
            O => \N__10527\,
            I => \DRA_c_1\
        );

    \I__2521\ : InMux
    port map (
            O => \N__10520\,
            I => \N__10514\
        );

    \I__2520\ : InMux
    port map (
            O => \N__10519\,
            I => \N__10514\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__10514\,
            I => \N__10511\
        );

    \I__2518\ : Span4Mux_v
    port map (
            O => \N__10511\,
            I => \N__10508\
        );

    \I__2517\ : Odrv4
    port map (
            O => \N__10508\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2516\ : InMux
    port map (
            O => \N__10505\,
            I => \N__10502\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__10502\,
            I => \N__10496\
        );

    \I__2514\ : InMux
    port map (
            O => \N__10501\,
            I => \N__10491\
        );

    \I__2513\ : InMux
    port map (
            O => \N__10500\,
            I => \N__10491\
        );

    \I__2512\ : InMux
    port map (
            O => \N__10499\,
            I => \N__10488\
        );

    \I__2511\ : Span4Mux_v
    port map (
            O => \N__10496\,
            I => \N__10485\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__10491\,
            I => \N__10480\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__10488\,
            I => \N__10480\
        );

    \I__2508\ : Span4Mux_h
    port map (
            O => \N__10485\,
            I => \N__10475\
        );

    \I__2507\ : Span4Mux_h
    port map (
            O => \N__10480\,
            I => \N__10475\
        );

    \I__2506\ : Sp12to4
    port map (
            O => \N__10475\,
            I => \N__10472\
        );

    \I__2505\ : Span12Mux_v
    port map (
            O => \N__10472\,
            I => \N__10469\
        );

    \I__2504\ : Odrv12
    port map (
            O => \N__10469\,
            I => \DRA_c_3\
        );

    \I__2503\ : InMux
    port map (
            O => \N__10466\,
            I => \N__10461\
        );

    \I__2502\ : InMux
    port map (
            O => \N__10465\,
            I => \N__10458\
        );

    \I__2501\ : InMux
    port map (
            O => \N__10464\,
            I => \N__10455\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__10461\,
            I => \N__10449\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__10458\,
            I => \N__10449\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__10455\,
            I => \N__10446\
        );

    \I__2497\ : InMux
    port map (
            O => \N__10454\,
            I => \N__10443\
        );

    \I__2496\ : Span4Mux_v
    port map (
            O => \N__10449\,
            I => \N__10440\
        );

    \I__2495\ : Span4Mux_v
    port map (
            O => \N__10446\,
            I => \N__10437\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__10443\,
            I => \N__10434\
        );

    \I__2493\ : Span4Mux_v
    port map (
            O => \N__10440\,
            I => \N__10431\
        );

    \I__2492\ : Sp12to4
    port map (
            O => \N__10437\,
            I => \N__10428\
        );

    \I__2491\ : Sp12to4
    port map (
            O => \N__10434\,
            I => \N__10425\
        );

    \I__2490\ : Sp12to4
    port map (
            O => \N__10431\,
            I => \N__10422\
        );

    \I__2489\ : Span12Mux_h
    port map (
            O => \N__10428\,
            I => \N__10419\
        );

    \I__2488\ : Span12Mux_v
    port map (
            O => \N__10425\,
            I => \N__10416\
        );

    \I__2487\ : Span12Mux_h
    port map (
            O => \N__10422\,
            I => \N__10413\
        );

    \I__2486\ : Span12Mux_v
    port map (
            O => \N__10419\,
            I => \N__10408\
        );

    \I__2485\ : Span12Mux_h
    port map (
            O => \N__10416\,
            I => \N__10408\
        );

    \I__2484\ : Odrv12
    port map (
            O => \N__10413\,
            I => \DRA_c_4\
        );

    \I__2483\ : Odrv12
    port map (
            O => \N__10408\,
            I => \DRA_c_4\
        );

    \I__2482\ : InMux
    port map (
            O => \N__10403\,
            I => \N__10400\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__10400\,
            I => \N__10397\
        );

    \I__2480\ : Span4Mux_h
    port map (
            O => \N__10397\,
            I => \N__10394\
        );

    \I__2479\ : Odrv4
    port map (
            O => \N__10394\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2478\ : IoInMux
    port map (
            O => \N__10391\,
            I => \N__10388\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__10388\,
            I => \N__10385\
        );

    \I__2476\ : Span4Mux_s0_v
    port map (
            O => \N__10385\,
            I => \N__10382\
        );

    \I__2475\ : Span4Mux_v
    port map (
            O => \N__10382\,
            I => \N__10379\
        );

    \I__2474\ : Odrv4
    port map (
            O => \N__10379\,
            I => \N_358_i\
        );

    \I__2473\ : InMux
    port map (
            O => \N__10376\,
            I => \N__10372\
        );

    \I__2472\ : InMux
    port map (
            O => \N__10375\,
            I => \N__10369\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__10372\,
            I => \N__10366\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__10369\,
            I => \N__10361\
        );

    \I__2469\ : Span4Mux_h
    port map (
            O => \N__10366\,
            I => \N__10361\
        );

    \I__2468\ : Sp12to4
    port map (
            O => \N__10361\,
            I => \N__10358\
        );

    \I__2467\ : Span12Mux_v
    port map (
            O => \N__10358\,
            I => \N__10354\
        );

    \I__2466\ : InMux
    port map (
            O => \N__10357\,
            I => \N__10351\
        );

    \I__2465\ : Odrv12
    port map (
            O => \N__10354\,
            I => \DS_ENm\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__10351\,
            I => \DS_ENm\
        );

    \I__2463\ : IoInMux
    port map (
            O => \N__10346\,
            I => \N__10343\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__10343\,
            I => \N__10340\
        );

    \I__2461\ : Span4Mux_s2_v
    port map (
            O => \N__10340\,
            I => \N__10337\
        );

    \I__2460\ : Span4Mux_v
    port map (
            O => \N__10337\,
            I => \N__10334\
        );

    \I__2459\ : Sp12to4
    port map (
            O => \N__10334\,
            I => \N__10331\
        );

    \I__2458\ : Odrv12
    port map (
            O => \N__10331\,
            I => \N_40\
        );

    \I__2457\ : InMux
    port map (
            O => \N__10328\,
            I => \N__10323\
        );

    \I__2456\ : InMux
    port map (
            O => \N__10327\,
            I => \N__10317\
        );

    \I__2455\ : InMux
    port map (
            O => \N__10326\,
            I => \N__10317\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__10323\,
            I => \N__10314\
        );

    \I__2453\ : InMux
    port map (
            O => \N__10322\,
            I => \N__10311\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__10317\,
            I => \N__10308\
        );

    \I__2451\ : Span4Mux_h
    port map (
            O => \N__10314\,
            I => \N__10301\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__10311\,
            I => \N__10301\
        );

    \I__2449\ : Span4Mux_v
    port map (
            O => \N__10308\,
            I => \N__10298\
        );

    \I__2448\ : InMux
    port map (
            O => \N__10307\,
            I => \N__10295\
        );

    \I__2447\ : InMux
    port map (
            O => \N__10306\,
            I => \N__10292\
        );

    \I__2446\ : Span4Mux_v
    port map (
            O => \N__10301\,
            I => \N__10288\
        );

    \I__2445\ : Span4Mux_v
    port map (
            O => \N__10298\,
            I => \N__10285\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__10295\,
            I => \N__10280\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__10292\,
            I => \N__10280\
        );

    \I__2442\ : InMux
    port map (
            O => \N__10291\,
            I => \N__10277\
        );

    \I__2441\ : Span4Mux_v
    port map (
            O => \N__10288\,
            I => \N__10273\
        );

    \I__2440\ : Span4Mux_v
    port map (
            O => \N__10285\,
            I => \N__10268\
        );

    \I__2439\ : Span4Mux_v
    port map (
            O => \N__10280\,
            I => \N__10268\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__10277\,
            I => \N__10265\
        );

    \I__2437\ : InMux
    port map (
            O => \N__10276\,
            I => \N__10262\
        );

    \I__2436\ : Sp12to4
    port map (
            O => \N__10273\,
            I => \N__10253\
        );

    \I__2435\ : Sp12to4
    port map (
            O => \N__10268\,
            I => \N__10253\
        );

    \I__2434\ : Sp12to4
    port map (
            O => \N__10265\,
            I => \N__10253\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__10262\,
            I => \N__10253\
        );

    \I__2432\ : Span12Mux_h
    port map (
            O => \N__10253\,
            I => \N__10250\
        );

    \I__2431\ : Odrv12
    port map (
            O => \N__10250\,
            I => \A_c_1\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__10247\,
            I => \N__10237\
        );

    \I__2429\ : CascadeMux
    port map (
            O => \N__10246\,
            I => \N__10233\
        );

    \I__2428\ : InMux
    port map (
            O => \N__10245\,
            I => \N__10230\
        );

    \I__2427\ : CascadeMux
    port map (
            O => \N__10244\,
            I => \N__10227\
        );

    \I__2426\ : InMux
    port map (
            O => \N__10243\,
            I => \N__10222\
        );

    \I__2425\ : InMux
    port map (
            O => \N__10242\,
            I => \N__10222\
        );

    \I__2424\ : InMux
    port map (
            O => \N__10241\,
            I => \N__10217\
        );

    \I__2423\ : InMux
    port map (
            O => \N__10240\,
            I => \N__10217\
        );

    \I__2422\ : InMux
    port map (
            O => \N__10237\,
            I => \N__10214\
        );

    \I__2421\ : InMux
    port map (
            O => \N__10236\,
            I => \N__10211\
        );

    \I__2420\ : InMux
    port map (
            O => \N__10233\,
            I => \N__10208\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__10230\,
            I => \N__10205\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10227\,
            I => \N__10202\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__10222\,
            I => \N__10193\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__10217\,
            I => \N__10193\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__10214\,
            I => \N__10193\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__10211\,
            I => \N__10193\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__10208\,
            I => \N__10190\
        );

    \I__2412\ : Span4Mux_v
    port map (
            O => \N__10205\,
            I => \N__10185\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__10202\,
            I => \N__10185\
        );

    \I__2410\ : Span4Mux_v
    port map (
            O => \N__10193\,
            I => \N__10182\
        );

    \I__2409\ : Span4Mux_v
    port map (
            O => \N__10190\,
            I => \N__10179\
        );

    \I__2408\ : Span4Mux_h
    port map (
            O => \N__10185\,
            I => \N__10176\
        );

    \I__2407\ : Sp12to4
    port map (
            O => \N__10182\,
            I => \N__10173\
        );

    \I__2406\ : Span4Mux_v
    port map (
            O => \N__10179\,
            I => \N__10170\
        );

    \I__2405\ : Span4Mux_v
    port map (
            O => \N__10176\,
            I => \N__10167\
        );

    \I__2404\ : Span12Mux_h
    port map (
            O => \N__10173\,
            I => \N__10160\
        );

    \I__2403\ : Sp12to4
    port map (
            O => \N__10170\,
            I => \N__10160\
        );

    \I__2402\ : Sp12to4
    port map (
            O => \N__10167\,
            I => \N__10160\
        );

    \I__2401\ : Odrv12
    port map (
            O => \N__10160\,
            I => \A_c_0\
        );

    \I__2400\ : InMux
    port map (
            O => \N__10157\,
            I => \N__10151\
        );

    \I__2399\ : InMux
    port map (
            O => \N__10156\,
            I => \N__10148\
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__10155\,
            I => \N__10144\
        );

    \I__2397\ : CascadeMux
    port map (
            O => \N__10154\,
            I => \N__10140\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__10151\,
            I => \N__10134\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__10148\,
            I => \N__10134\
        );

    \I__2394\ : InMux
    port map (
            O => \N__10147\,
            I => \N__10131\
        );

    \I__2393\ : InMux
    port map (
            O => \N__10144\,
            I => \N__10128\
        );

    \I__2392\ : InMux
    port map (
            O => \N__10143\,
            I => \N__10123\
        );

    \I__2391\ : InMux
    port map (
            O => \N__10140\,
            I => \N__10123\
        );

    \I__2390\ : InMux
    port map (
            O => \N__10139\,
            I => \N__10118\
        );

    \I__2389\ : Span4Mux_v
    port map (
            O => \N__10134\,
            I => \N__10115\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__10131\,
            I => \N__10110\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__10128\,
            I => \N__10110\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__10123\,
            I => \N__10107\
        );

    \I__2385\ : InMux
    port map (
            O => \N__10122\,
            I => \N__10102\
        );

    \I__2384\ : InMux
    port map (
            O => \N__10121\,
            I => \N__10102\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__10118\,
            I => \N__10099\
        );

    \I__2382\ : Span4Mux_v
    port map (
            O => \N__10115\,
            I => \N__10096\
        );

    \I__2381\ : Span4Mux_v
    port map (
            O => \N__10110\,
            I => \N__10089\
        );

    \I__2380\ : Span4Mux_h
    port map (
            O => \N__10107\,
            I => \N__10089\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__10102\,
            I => \N__10089\
        );

    \I__2378\ : Span4Mux_v
    port map (
            O => \N__10099\,
            I => \N__10086\
        );

    \I__2377\ : Span4Mux_v
    port map (
            O => \N__10096\,
            I => \N__10081\
        );

    \I__2376\ : Span4Mux_h
    port map (
            O => \N__10089\,
            I => \N__10081\
        );

    \I__2375\ : Span4Mux_v
    port map (
            O => \N__10086\,
            I => \N__10078\
        );

    \I__2374\ : Span4Mux_v
    port map (
            O => \N__10081\,
            I => \N__10075\
        );

    \I__2373\ : Span4Mux_v
    port map (
            O => \N__10078\,
            I => \N__10072\
        );

    \I__2372\ : Span4Mux_h
    port map (
            O => \N__10075\,
            I => \N__10069\
        );

    \I__2371\ : Sp12to4
    port map (
            O => \N__10072\,
            I => \N__10064\
        );

    \I__2370\ : Sp12to4
    port map (
            O => \N__10069\,
            I => \N__10064\
        );

    \I__2369\ : Odrv12
    port map (
            O => \N__10064\,
            I => \SIZ_c_0\
        );

    \I__2368\ : InMux
    port map (
            O => \N__10061\,
            I => \N__10056\
        );

    \I__2367\ : InMux
    port map (
            O => \N__10060\,
            I => \N__10052\
        );

    \I__2366\ : InMux
    port map (
            O => \N__10059\,
            I => \N__10049\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__10056\,
            I => \N__10045\
        );

    \I__2364\ : InMux
    port map (
            O => \N__10055\,
            I => \N__10042\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__10052\,
            I => \N__10039\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__10049\,
            I => \N__10036\
        );

    \I__2361\ : CascadeMux
    port map (
            O => \N__10048\,
            I => \N__10032\
        );

    \I__2360\ : Span4Mux_h
    port map (
            O => \N__10045\,
            I => \N__10027\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__10042\,
            I => \N__10027\
        );

    \I__2358\ : Span4Mux_v
    port map (
            O => \N__10039\,
            I => \N__10024\
        );

    \I__2357\ : Span4Mux_h
    port map (
            O => \N__10036\,
            I => \N__10021\
        );

    \I__2356\ : InMux
    port map (
            O => \N__10035\,
            I => \N__10018\
        );

    \I__2355\ : InMux
    port map (
            O => \N__10032\,
            I => \N__10015\
        );

    \I__2354\ : Sp12to4
    port map (
            O => \N__10027\,
            I => \N__10012\
        );

    \I__2353\ : Span4Mux_v
    port map (
            O => \N__10024\,
            I => \N__10009\
        );

    \I__2352\ : Span4Mux_v
    port map (
            O => \N__10021\,
            I => \N__10006\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__10018\,
            I => \N__10001\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__10015\,
            I => \N__10001\
        );

    \I__2349\ : Span12Mux_v
    port map (
            O => \N__10012\,
            I => \N__9998\
        );

    \I__2348\ : Sp12to4
    port map (
            O => \N__10009\,
            I => \N__9991\
        );

    \I__2347\ : Sp12to4
    port map (
            O => \N__10006\,
            I => \N__9991\
        );

    \I__2346\ : Span12Mux_v
    port map (
            O => \N__10001\,
            I => \N__9991\
        );

    \I__2345\ : Span12Mux_h
    port map (
            O => \N__9998\,
            I => \N__9988\
        );

    \I__2344\ : Span12Mux_h
    port map (
            O => \N__9991\,
            I => \N__9985\
        );

    \I__2343\ : Odrv12
    port map (
            O => \N__9988\,
            I => \SIZ_c_1\
        );

    \I__2342\ : Odrv12
    port map (
            O => \N__9985\,
            I => \SIZ_c_1\
        );

    \I__2341\ : IoInMux
    port map (
            O => \N__9980\,
            I => \N__9977\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__9977\,
            I => \N__9974\
        );

    \I__2339\ : Span4Mux_s3_v
    port map (
            O => \N__9974\,
            I => \N__9971\
        );

    \I__2338\ : Odrv4
    port map (
            O => \N__9971\,
            I => \LLBEn_c\
        );

    \I__2337\ : InMux
    port map (
            O => \N__9968\,
            I => \N__9964\
        );

    \I__2336\ : InMux
    port map (
            O => \N__9967\,
            I => \N__9960\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__9964\,
            I => \N__9955\
        );

    \I__2334\ : InMux
    port map (
            O => \N__9963\,
            I => \N__9952\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__9960\,
            I => \N__9949\
        );

    \I__2332\ : InMux
    port map (
            O => \N__9959\,
            I => \N__9944\
        );

    \I__2331\ : InMux
    port map (
            O => \N__9958\,
            I => \N__9944\
        );

    \I__2330\ : Span4Mux_v
    port map (
            O => \N__9955\,
            I => \N__9939\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__9952\,
            I => \N__9939\
        );

    \I__2328\ : Span4Mux_v
    port map (
            O => \N__9949\,
            I => \N__9934\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__9944\,
            I => \N__9934\
        );

    \I__2326\ : Span4Mux_h
    port map (
            O => \N__9939\,
            I => \N__9930\
        );

    \I__2325\ : Span4Mux_h
    port map (
            O => \N__9934\,
            I => \N__9927\
        );

    \I__2324\ : InMux
    port map (
            O => \N__9933\,
            I => \N__9924\
        );

    \I__2323\ : Odrv4
    port map (
            O => \N__9930\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2322\ : Odrv4
    port map (
            O => \N__9927\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__9924\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2320\ : IoInMux
    port map (
            O => \N__9917\,
            I => \N__9914\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__9914\,
            I => \N__9911\
        );

    \I__2318\ : Span4Mux_s3_h
    port map (
            O => \N__9911\,
            I => \N__9908\
        );

    \I__2317\ : Span4Mux_v
    port map (
            O => \N__9908\,
            I => \N__9905\
        );

    \I__2316\ : Span4Mux_v
    port map (
            O => \N__9905\,
            I => \N__9902\
        );

    \I__2315\ : Sp12to4
    port map (
            O => \N__9902\,
            I => \N__9899\
        );

    \I__2314\ : Odrv12
    port map (
            O => \N__9899\,
            I => \WEn_c\
        );

    \I__2313\ : InMux
    port map (
            O => \N__9896\,
            I => \N__9890\
        );

    \I__2312\ : CascadeMux
    port map (
            O => \N__9895\,
            I => \N__9886\
        );

    \I__2311\ : InMux
    port map (
            O => \N__9894\,
            I => \N__9883\
        );

    \I__2310\ : InMux
    port map (
            O => \N__9893\,
            I => \N__9880\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__9890\,
            I => \N__9877\
        );

    \I__2308\ : InMux
    port map (
            O => \N__9889\,
            I => \N__9872\
        );

    \I__2307\ : InMux
    port map (
            O => \N__9886\,
            I => \N__9872\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__9883\,
            I => \N__9869\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__9880\,
            I => \N__9866\
        );

    \I__2304\ : Span4Mux_v
    port map (
            O => \N__9877\,
            I => \N__9861\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__9872\,
            I => \N__9861\
        );

    \I__2302\ : Span4Mux_h
    port map (
            O => \N__9869\,
            I => \N__9855\
        );

    \I__2301\ : Span4Mux_h
    port map (
            O => \N__9866\,
            I => \N__9855\
        );

    \I__2300\ : Span4Mux_h
    port map (
            O => \N__9861\,
            I => \N__9852\
        );

    \I__2299\ : InMux
    port map (
            O => \N__9860\,
            I => \N__9849\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__9855\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2297\ : Odrv4
    port map (
            O => \N__9852\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__9849\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2295\ : IoInMux
    port map (
            O => \N__9842\,
            I => \N__9839\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__9839\,
            I => \N__9836\
        );

    \I__2293\ : Span4Mux_s1_v
    port map (
            O => \N__9836\,
            I => \N__9833\
        );

    \I__2292\ : Span4Mux_v
    port map (
            O => \N__9833\,
            I => \N__9830\
        );

    \I__2291\ : Span4Mux_v
    port map (
            O => \N__9830\,
            I => \N__9827\
        );

    \I__2290\ : Span4Mux_h
    port map (
            O => \N__9827\,
            I => \N__9824\
        );

    \I__2289\ : Odrv4
    port map (
            O => \N__9824\,
            I => \RASn_c\
        );

    \I__2288\ : InMux
    port map (
            O => \N__9821\,
            I => \N__9818\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__9818\,
            I => \N__9797\
        );

    \I__2286\ : ClkMux
    port map (
            O => \N__9817\,
            I => \N__9713\
        );

    \I__2285\ : ClkMux
    port map (
            O => \N__9816\,
            I => \N__9713\
        );

    \I__2284\ : ClkMux
    port map (
            O => \N__9815\,
            I => \N__9713\
        );

    \I__2283\ : ClkMux
    port map (
            O => \N__9814\,
            I => \N__9713\
        );

    \I__2282\ : ClkMux
    port map (
            O => \N__9813\,
            I => \N__9713\
        );

    \I__2281\ : ClkMux
    port map (
            O => \N__9812\,
            I => \N__9713\
        );

    \I__2280\ : ClkMux
    port map (
            O => \N__9811\,
            I => \N__9713\
        );

    \I__2279\ : ClkMux
    port map (
            O => \N__9810\,
            I => \N__9713\
        );

    \I__2278\ : ClkMux
    port map (
            O => \N__9809\,
            I => \N__9713\
        );

    \I__2277\ : ClkMux
    port map (
            O => \N__9808\,
            I => \N__9713\
        );

    \I__2276\ : ClkMux
    port map (
            O => \N__9807\,
            I => \N__9713\
        );

    \I__2275\ : ClkMux
    port map (
            O => \N__9806\,
            I => \N__9713\
        );

    \I__2274\ : ClkMux
    port map (
            O => \N__9805\,
            I => \N__9713\
        );

    \I__2273\ : ClkMux
    port map (
            O => \N__9804\,
            I => \N__9713\
        );

    \I__2272\ : ClkMux
    port map (
            O => \N__9803\,
            I => \N__9713\
        );

    \I__2271\ : ClkMux
    port map (
            O => \N__9802\,
            I => \N__9713\
        );

    \I__2270\ : ClkMux
    port map (
            O => \N__9801\,
            I => \N__9713\
        );

    \I__2269\ : ClkMux
    port map (
            O => \N__9800\,
            I => \N__9713\
        );

    \I__2268\ : Glb2LocalMux
    port map (
            O => \N__9797\,
            I => \N__9713\
        );

    \I__2267\ : ClkMux
    port map (
            O => \N__9796\,
            I => \N__9713\
        );

    \I__2266\ : ClkMux
    port map (
            O => \N__9795\,
            I => \N__9713\
        );

    \I__2265\ : ClkMux
    port map (
            O => \N__9794\,
            I => \N__9713\
        );

    \I__2264\ : ClkMux
    port map (
            O => \N__9793\,
            I => \N__9713\
        );

    \I__2263\ : ClkMux
    port map (
            O => \N__9792\,
            I => \N__9713\
        );

    \I__2262\ : ClkMux
    port map (
            O => \N__9791\,
            I => \N__9713\
        );

    \I__2261\ : ClkMux
    port map (
            O => \N__9790\,
            I => \N__9713\
        );

    \I__2260\ : ClkMux
    port map (
            O => \N__9789\,
            I => \N__9713\
        );

    \I__2259\ : ClkMux
    port map (
            O => \N__9788\,
            I => \N__9713\
        );

    \I__2258\ : ClkMux
    port map (
            O => \N__9787\,
            I => \N__9713\
        );

    \I__2257\ : ClkMux
    port map (
            O => \N__9786\,
            I => \N__9713\
        );

    \I__2256\ : ClkMux
    port map (
            O => \N__9785\,
            I => \N__9713\
        );

    \I__2255\ : ClkMux
    port map (
            O => \N__9784\,
            I => \N__9713\
        );

    \I__2254\ : ClkMux
    port map (
            O => \N__9783\,
            I => \N__9713\
        );

    \I__2253\ : ClkMux
    port map (
            O => \N__9782\,
            I => \N__9713\
        );

    \I__2252\ : GlobalMux
    port map (
            O => \N__9713\,
            I => \CLK80_PLL\
        );

    \I__2251\ : CascadeMux
    port map (
            O => \N__9710\,
            I => \N__9700\
        );

    \I__2250\ : InMux
    port map (
            O => \N__9709\,
            I => \N__9696\
        );

    \I__2249\ : CascadeMux
    port map (
            O => \N__9708\,
            I => \N__9691\
        );

    \I__2248\ : InMux
    port map (
            O => \N__9707\,
            I => \N__9686\
        );

    \I__2247\ : InMux
    port map (
            O => \N__9706\,
            I => \N__9683\
        );

    \I__2246\ : InMux
    port map (
            O => \N__9705\,
            I => \N__9678\
        );

    \I__2245\ : InMux
    port map (
            O => \N__9704\,
            I => \N__9675\
        );

    \I__2244\ : InMux
    port map (
            O => \N__9703\,
            I => \N__9670\
        );

    \I__2243\ : InMux
    port map (
            O => \N__9700\,
            I => \N__9665\
        );

    \I__2242\ : InMux
    port map (
            O => \N__9699\,
            I => \N__9665\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__9696\,
            I => \N__9662\
        );

    \I__2240\ : CascadeMux
    port map (
            O => \N__9695\,
            I => \N__9658\
        );

    \I__2239\ : InMux
    port map (
            O => \N__9694\,
            I => \N__9653\
        );

    \I__2238\ : InMux
    port map (
            O => \N__9691\,
            I => \N__9646\
        );

    \I__2237\ : InMux
    port map (
            O => \N__9690\,
            I => \N__9646\
        );

    \I__2236\ : InMux
    port map (
            O => \N__9689\,
            I => \N__9646\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__9686\,
            I => \N__9639\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__9683\,
            I => \N__9639\
        );

    \I__2233\ : CascadeMux
    port map (
            O => \N__9682\,
            I => \N__9634\
        );

    \I__2232\ : InMux
    port map (
            O => \N__9681\,
            I => \N__9631\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__9678\,
            I => \N__9626\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__9675\,
            I => \N__9626\
        );

    \I__2229\ : InMux
    port map (
            O => \N__9674\,
            I => \N__9621\
        );

    \I__2228\ : InMux
    port map (
            O => \N__9673\,
            I => \N__9621\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__9670\,
            I => \N__9618\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__9665\,
            I => \N__9613\
        );

    \I__2225\ : Span4Mux_v
    port map (
            O => \N__9662\,
            I => \N__9613\
        );

    \I__2224\ : InMux
    port map (
            O => \N__9661\,
            I => \N__9608\
        );

    \I__2223\ : InMux
    port map (
            O => \N__9658\,
            I => \N__9608\
        );

    \I__2222\ : InMux
    port map (
            O => \N__9657\,
            I => \N__9603\
        );

    \I__2221\ : InMux
    port map (
            O => \N__9656\,
            I => \N__9603\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__9653\,
            I => \N__9598\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__9646\,
            I => \N__9598\
        );

    \I__2218\ : InMux
    port map (
            O => \N__9645\,
            I => \N__9595\
        );

    \I__2217\ : InMux
    port map (
            O => \N__9644\,
            I => \N__9592\
        );

    \I__2216\ : Span4Mux_v
    port map (
            O => \N__9639\,
            I => \N__9589\
        );

    \I__2215\ : InMux
    port map (
            O => \N__9638\,
            I => \N__9586\
        );

    \I__2214\ : InMux
    port map (
            O => \N__9637\,
            I => \N__9581\
        );

    \I__2213\ : InMux
    port map (
            O => \N__9634\,
            I => \N__9581\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__9631\,
            I => \N__9578\
        );

    \I__2211\ : Span12Mux_v
    port map (
            O => \N__9626\,
            I => \N__9573\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__9621\,
            I => \N__9573\
        );

    \I__2209\ : Span4Mux_v
    port map (
            O => \N__9618\,
            I => \N__9568\
        );

    \I__2208\ : Span4Mux_h
    port map (
            O => \N__9613\,
            I => \N__9568\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__9608\,
            I => \N__9561\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__9603\,
            I => \N__9561\
        );

    \I__2205\ : Span4Mux_v
    port map (
            O => \N__9598\,
            I => \N__9561\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__9595\,
            I => \N__9556\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__9592\,
            I => \N__9556\
        );

    \I__2202\ : Odrv4
    port map (
            O => \N__9589\,
            I => \CPU_CYCLEm\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__9586\,
            I => \CPU_CYCLEm\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__9581\,
            I => \CPU_CYCLEm\
        );

    \I__2199\ : Odrv4
    port map (
            O => \N__9578\,
            I => \CPU_CYCLEm\
        );

    \I__2198\ : Odrv12
    port map (
            O => \N__9573\,
            I => \CPU_CYCLEm\
        );

    \I__2197\ : Odrv4
    port map (
            O => \N__9568\,
            I => \CPU_CYCLEm\
        );

    \I__2196\ : Odrv4
    port map (
            O => \N__9561\,
            I => \CPU_CYCLEm\
        );

    \I__2195\ : Odrv12
    port map (
            O => \N__9556\,
            I => \CPU_CYCLEm\
        );

    \I__2194\ : InMux
    port map (
            O => \N__9539\,
            I => \N__9536\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__9536\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\
        );

    \I__2192\ : CascadeMux
    port map (
            O => \N__9533\,
            I => \N__9528\
        );

    \I__2191\ : InMux
    port map (
            O => \N__9532\,
            I => \N__9516\
        );

    \I__2190\ : CascadeMux
    port map (
            O => \N__9531\,
            I => \N__9513\
        );

    \I__2189\ : InMux
    port map (
            O => \N__9528\,
            I => \N__9509\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__9527\,
            I => \N__9506\
        );

    \I__2187\ : CascadeMux
    port map (
            O => \N__9526\,
            I => \N__9503\
        );

    \I__2186\ : InMux
    port map (
            O => \N__9525\,
            I => \N__9499\
        );

    \I__2185\ : CascadeMux
    port map (
            O => \N__9524\,
            I => \N__9495\
        );

    \I__2184\ : InMux
    port map (
            O => \N__9523\,
            I => \N__9489\
        );

    \I__2183\ : InMux
    port map (
            O => \N__9522\,
            I => \N__9484\
        );

    \I__2182\ : InMux
    port map (
            O => \N__9521\,
            I => \N__9484\
        );

    \I__2181\ : InMux
    port map (
            O => \N__9520\,
            I => \N__9479\
        );

    \I__2180\ : InMux
    port map (
            O => \N__9519\,
            I => \N__9479\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__9516\,
            I => \N__9476\
        );

    \I__2178\ : InMux
    port map (
            O => \N__9513\,
            I => \N__9471\
        );

    \I__2177\ : InMux
    port map (
            O => \N__9512\,
            I => \N__9471\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__9509\,
            I => \N__9468\
        );

    \I__2175\ : InMux
    port map (
            O => \N__9506\,
            I => \N__9465\
        );

    \I__2174\ : InMux
    port map (
            O => \N__9503\,
            I => \N__9461\
        );

    \I__2173\ : InMux
    port map (
            O => \N__9502\,
            I => \N__9458\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__9499\,
            I => \N__9455\
        );

    \I__2171\ : InMux
    port map (
            O => \N__9498\,
            I => \N__9448\
        );

    \I__2170\ : InMux
    port map (
            O => \N__9495\,
            I => \N__9448\
        );

    \I__2169\ : InMux
    port map (
            O => \N__9494\,
            I => \N__9448\
        );

    \I__2168\ : InMux
    port map (
            O => \N__9493\,
            I => \N__9443\
        );

    \I__2167\ : InMux
    port map (
            O => \N__9492\,
            I => \N__9443\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__9489\,
            I => \N__9437\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__9484\,
            I => \N__9437\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__9479\,
            I => \N__9432\
        );

    \I__2163\ : Span4Mux_v
    port map (
            O => \N__9476\,
            I => \N__9432\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__9471\,
            I => \N__9427\
        );

    \I__2161\ : Span4Mux_h
    port map (
            O => \N__9468\,
            I => \N__9427\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__9465\,
            I => \N__9424\
        );

    \I__2159\ : InMux
    port map (
            O => \N__9464\,
            I => \N__9421\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__9461\,
            I => \N__9406\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__9458\,
            I => \N__9406\
        );

    \I__2156\ : Span4Mux_h
    port map (
            O => \N__9455\,
            I => \N__9406\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__9448\,
            I => \N__9406\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__9443\,
            I => \N__9406\
        );

    \I__2153\ : InMux
    port map (
            O => \N__9442\,
            I => \N__9403\
        );

    \I__2152\ : Span4Mux_v
    port map (
            O => \N__9437\,
            I => \N__9400\
        );

    \I__2151\ : Span4Mux_h
    port map (
            O => \N__9432\,
            I => \N__9397\
        );

    \I__2150\ : Span4Mux_h
    port map (
            O => \N__9427\,
            I => \N__9394\
        );

    \I__2149\ : Span4Mux_h
    port map (
            O => \N__9424\,
            I => \N__9389\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__9421\,
            I => \N__9389\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9420\,
            I => \N__9382\
        );

    \I__2146\ : InMux
    port map (
            O => \N__9419\,
            I => \N__9382\
        );

    \I__2145\ : InMux
    port map (
            O => \N__9418\,
            I => \N__9382\
        );

    \I__2144\ : InMux
    port map (
            O => \N__9417\,
            I => \N__9379\
        );

    \I__2143\ : Span4Mux_v
    port map (
            O => \N__9406\,
            I => \N__9374\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__9403\,
            I => \N__9374\
        );

    \I__2141\ : Odrv4
    port map (
            O => \N__9400\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2140\ : Odrv4
    port map (
            O => \N__9397\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2139\ : Odrv4
    port map (
            O => \N__9394\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2138\ : Odrv4
    port map (
            O => \N__9389\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__9382\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9379\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2135\ : Odrv4
    port map (
            O => \N__9374\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2134\ : InMux
    port map (
            O => \N__9359\,
            I => \N__9356\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__9356\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__2132\ : InMux
    port map (
            O => \N__9353\,
            I => \N__9350\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__9350\,
            I => \N__9347\
        );

    \I__2130\ : Span4Mux_h
    port map (
            O => \N__9347\,
            I => \N__9344\
        );

    \I__2129\ : Odrv4
    port map (
            O => \N__9344\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9341\,
            I => \N__9338\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__9338\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9335\,
            I => \N__9332\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__9332\,
            I => \N__9329\
        );

    \I__2124\ : Span4Mux_h
    port map (
            O => \N__9329\,
            I => \N__9326\
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__9326\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__2122\ : InMux
    port map (
            O => \N__9323\,
            I => \N__9316\
        );

    \I__2121\ : InMux
    port map (
            O => \N__9322\,
            I => \N__9316\
        );

    \I__2120\ : InMux
    port map (
            O => \N__9321\,
            I => \N__9313\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__9316\,
            I => \N__9310\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__9313\,
            I => \N__9307\
        );

    \I__2117\ : Span4Mux_v
    port map (
            O => \N__9310\,
            I => \N__9303\
        );

    \I__2116\ : Span4Mux_h
    port map (
            O => \N__9307\,
            I => \N__9300\
        );

    \I__2115\ : InMux
    port map (
            O => \N__9306\,
            I => \N__9297\
        );

    \I__2114\ : Span4Mux_v
    port map (
            O => \N__9303\,
            I => \N__9294\
        );

    \I__2113\ : Span4Mux_v
    port map (
            O => \N__9300\,
            I => \N__9291\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__9297\,
            I => \N__9288\
        );

    \I__2111\ : Sp12to4
    port map (
            O => \N__9294\,
            I => \N__9281\
        );

    \I__2110\ : Sp12to4
    port map (
            O => \N__9291\,
            I => \N__9281\
        );

    \I__2109\ : Span12Mux_v
    port map (
            O => \N__9288\,
            I => \N__9281\
        );

    \I__2108\ : Span12Mux_h
    port map (
            O => \N__9281\,
            I => \N__9278\
        );

    \I__2107\ : Odrv12
    port map (
            O => \N__9278\,
            I => \DRA_c_6\
        );

    \I__2106\ : InMux
    port map (
            O => \N__9275\,
            I => \N__9271\
        );

    \I__2105\ : InMux
    port map (
            O => \N__9274\,
            I => \N__9268\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__9271\,
            I => \N__9262\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__9268\,
            I => \N__9262\
        );

    \I__2102\ : InMux
    port map (
            O => \N__9267\,
            I => \N__9259\
        );

    \I__2101\ : Span4Mux_v
    port map (
            O => \N__9262\,
            I => \N__9255\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__9259\,
            I => \N__9252\
        );

    \I__2099\ : InMux
    port map (
            O => \N__9258\,
            I => \N__9249\
        );

    \I__2098\ : Span4Mux_v
    port map (
            O => \N__9255\,
            I => \N__9246\
        );

    \I__2097\ : Sp12to4
    port map (
            O => \N__9252\,
            I => \N__9241\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__9249\,
            I => \N__9241\
        );

    \I__2095\ : Sp12to4
    port map (
            O => \N__9246\,
            I => \N__9236\
        );

    \I__2094\ : Span12Mux_v
    port map (
            O => \N__9241\,
            I => \N__9236\
        );

    \I__2093\ : Span12Mux_h
    port map (
            O => \N__9236\,
            I => \N__9233\
        );

    \I__2092\ : Odrv12
    port map (
            O => \N__9233\,
            I => \DRA_c_5\
        );

    \I__2091\ : InMux
    port map (
            O => \N__9230\,
            I => \N__9227\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__9227\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2089\ : InMux
    port map (
            O => \N__9224\,
            I => \N__9220\
        );

    \I__2088\ : InMux
    port map (
            O => \N__9223\,
            I => \N__9217\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__9220\,
            I => \N__9211\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__9217\,
            I => \N__9211\
        );

    \I__2085\ : InMux
    port map (
            O => \N__9216\,
            I => \N__9208\
        );

    \I__2084\ : Span4Mux_v
    port map (
            O => \N__9211\,
            I => \N__9204\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__9208\,
            I => \N__9201\
        );

    \I__2082\ : InMux
    port map (
            O => \N__9207\,
            I => \N__9198\
        );

    \I__2081\ : Sp12to4
    port map (
            O => \N__9204\,
            I => \N__9193\
        );

    \I__2080\ : Span12Mux_v
    port map (
            O => \N__9201\,
            I => \N__9193\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__9198\,
            I => \N__9190\
        );

    \I__2078\ : Span12Mux_h
    port map (
            O => \N__9193\,
            I => \N__9187\
        );

    \I__2077\ : Span12Mux_h
    port map (
            O => \N__9190\,
            I => \N__9184\
        );

    \I__2076\ : Odrv12
    port map (
            O => \N__9187\,
            I => \DRA_c_8\
        );

    \I__2075\ : Odrv12
    port map (
            O => \N__9184\,
            I => \DRA_c_8\
        );

    \I__2074\ : InMux
    port map (
            O => \N__9179\,
            I => \N__9176\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__9176\,
            I => \N__9173\
        );

    \I__2072\ : Odrv4
    port map (
            O => \N__9173\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2071\ : InMux
    port map (
            O => \N__9170\,
            I => \N__9167\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__9167\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__2069\ : CascadeMux
    port map (
            O => \N__9164\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_\
        );

    \I__2068\ : InMux
    port map (
            O => \N__9161\,
            I => \N__9158\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__9158\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__2066\ : IoInMux
    port map (
            O => \N__9155\,
            I => \N__9152\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__9152\,
            I => \N__9149\
        );

    \I__2064\ : IoSpan4Mux
    port map (
            O => \N__9149\,
            I => \N__9146\
        );

    \I__2063\ : Span4Mux_s3_v
    port map (
            O => \N__9146\,
            I => \N__9143\
        );

    \I__2062\ : Span4Mux_v
    port map (
            O => \N__9143\,
            I => \N__9140\
        );

    \I__2061\ : Odrv4
    port map (
            O => \N__9140\,
            I => \CMA_c_1\
        );

    \I__2060\ : CEMux
    port map (
            O => \N__9137\,
            I => \N__9134\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__9134\,
            I => \N__9131\
        );

    \I__2058\ : Span4Mux_h
    port map (
            O => \N__9131\,
            I => \N__9124\
        );

    \I__2057\ : CEMux
    port map (
            O => \N__9130\,
            I => \N__9121\
        );

    \I__2056\ : CEMux
    port map (
            O => \N__9129\,
            I => \N__9118\
        );

    \I__2055\ : CEMux
    port map (
            O => \N__9128\,
            I => \N__9115\
        );

    \I__2054\ : CEMux
    port map (
            O => \N__9127\,
            I => \N__9112\
        );

    \I__2053\ : Odrv4
    port map (
            O => \N__9124\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__9121\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__9118\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__9115\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__9112\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2048\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9098\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__9098\,
            I => \N__9095\
        );

    \I__2046\ : Span4Mux_v
    port map (
            O => \N__9095\,
            I => \N__9092\
        );

    \I__2045\ : Sp12to4
    port map (
            O => \N__9092\,
            I => \N__9089\
        );

    \I__2044\ : Span12Mux_h
    port map (
            O => \N__9089\,
            I => \N__9086\
        );

    \I__2043\ : Odrv12
    port map (
            O => \N__9086\,
            I => \A_c_13\
        );

    \I__2042\ : InMux
    port map (
            O => \N__9083\,
            I => \N__9080\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__9080\,
            I => \N__9077\
        );

    \I__2040\ : Sp12to4
    port map (
            O => \N__9077\,
            I => \N__9074\
        );

    \I__2039\ : Span12Mux_v
    port map (
            O => \N__9074\,
            I => \N__9071\
        );

    \I__2038\ : Span12Mux_h
    port map (
            O => \N__9071\,
            I => \N__9068\
        );

    \I__2037\ : Odrv12
    port map (
            O => \N__9068\,
            I => \A_c_6\
        );

    \I__2036\ : InMux
    port map (
            O => \N__9065\,
            I => \N__9062\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__9062\,
            I => \N__9059\
        );

    \I__2034\ : Span4Mux_h
    port map (
            O => \N__9059\,
            I => \N__9056\
        );

    \I__2033\ : Odrv4
    port map (
            O => \N__9056\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__2032\ : CascadeMux
    port map (
            O => \N__9053\,
            I => \N__9050\
        );

    \I__2031\ : InMux
    port map (
            O => \N__9050\,
            I => \N__9047\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__9047\,
            I => \N__9044\
        );

    \I__2029\ : Odrv4
    port map (
            O => \N__9044\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2028\ : InMux
    port map (
            O => \N__9041\,
            I => \N__9036\
        );

    \I__2027\ : InMux
    port map (
            O => \N__9040\,
            I => \N__9033\
        );

    \I__2026\ : InMux
    port map (
            O => \N__9039\,
            I => \N__9030\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__9036\,
            I => \N__9027\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__9033\,
            I => \N__9019\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__9030\,
            I => \N__9019\
        );

    \I__2022\ : Span4Mux_h
    port map (
            O => \N__9027\,
            I => \N__9019\
        );

    \I__2021\ : InMux
    port map (
            O => \N__9026\,
            I => \N__9016\
        );

    \I__2020\ : Sp12to4
    port map (
            O => \N__9019\,
            I => \N__9011\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__9016\,
            I => \N__9011\
        );

    \I__2018\ : Span12Mux_v
    port map (
            O => \N__9011\,
            I => \N__9008\
        );

    \I__2017\ : Span12Mux_h
    port map (
            O => \N__9008\,
            I => \N__9005\
        );

    \I__2016\ : Odrv12
    port map (
            O => \N__9005\,
            I => \DRA_c_7\
        );

    \I__2015\ : InMux
    port map (
            O => \N__9002\,
            I => \N__8999\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__8999\,
            I => \N__8996\
        );

    \I__2013\ : Span4Mux_h
    port map (
            O => \N__8996\,
            I => \N__8993\
        );

    \I__2012\ : Odrv4
    port map (
            O => \N__8993\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2011\ : InMux
    port map (
            O => \N__8990\,
            I => \N__8987\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__8987\,
            I => \N__8984\
        );

    \I__2009\ : Span4Mux_v
    port map (
            O => \N__8984\,
            I => \N__8981\
        );

    \I__2008\ : Span4Mux_h
    port map (
            O => \N__8981\,
            I => \N__8978\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__8978\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2006\ : InMux
    port map (
            O => \N__8975\,
            I => \N__8972\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__8972\,
            I => \N__8969\
        );

    \I__2004\ : Span4Mux_h
    port map (
            O => \N__8969\,
            I => \N__8966\
        );

    \I__2003\ : Span4Mux_v
    port map (
            O => \N__8966\,
            I => \N__8963\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__8963\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__2001\ : InMux
    port map (
            O => \N__8960\,
            I => \N__8957\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__8957\,
            I => \N__8953\
        );

    \I__1999\ : InMux
    port map (
            O => \N__8956\,
            I => \N__8950\
        );

    \I__1998\ : Span4Mux_v
    port map (
            O => \N__8953\,
            I => \N__8945\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__8950\,
            I => \N__8945\
        );

    \I__1996\ : Span4Mux_h
    port map (
            O => \N__8945\,
            I => \N__8942\
        );

    \I__1995\ : Sp12to4
    port map (
            O => \N__8942\,
            I => \N__8939\
        );

    \I__1994\ : Span12Mux_h
    port map (
            O => \N__8939\,
            I => \N__8936\
        );

    \I__1993\ : Span12Mux_v
    port map (
            O => \N__8936\,
            I => \N__8933\
        );

    \I__1992\ : Odrv12
    port map (
            O => \N__8933\,
            I => \DRA_c_0\
        );

    \I__1991\ : InMux
    port map (
            O => \N__8930\,
            I => \N__8927\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__8927\,
            I => \N__8924\
        );

    \I__1989\ : Odrv12
    port map (
            O => \N__8924\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__1988\ : IoInMux
    port map (
            O => \N__8921\,
            I => \N__8918\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__8918\,
            I => \N__8915\
        );

    \I__1986\ : Span4Mux_s3_v
    port map (
            O => \N__8915\,
            I => \N__8912\
        );

    \I__1985\ : Span4Mux_v
    port map (
            O => \N__8912\,
            I => \N__8909\
        );

    \I__1984\ : Sp12to4
    port map (
            O => \N__8909\,
            I => \N__8906\
        );

    \I__1983\ : Span12Mux_h
    port map (
            O => \N__8906\,
            I => \N__8903\
        );

    \I__1982\ : Odrv12
    port map (
            O => \N__8903\,
            I => \CASn_c\
        );

    \I__1981\ : InMux
    port map (
            O => \N__8900\,
            I => \N__8897\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__8897\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__1979\ : IoInMux
    port map (
            O => \N__8894\,
            I => \N__8891\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__8891\,
            I => \N__8888\
        );

    \I__1977\ : Span4Mux_s2_v
    port map (
            O => \N__8888\,
            I => \N__8885\
        );

    \I__1976\ : Span4Mux_v
    port map (
            O => \N__8885\,
            I => \N__8882\
        );

    \I__1975\ : Span4Mux_h
    port map (
            O => \N__8882\,
            I => \N__8879\
        );

    \I__1974\ : Odrv4
    port map (
            O => \N__8879\,
            I => \CMA_c_0\
        );

    \I__1973\ : InMux
    port map (
            O => \N__8876\,
            I => \N__8872\
        );

    \I__1972\ : InMux
    port map (
            O => \N__8875\,
            I => \N__8868\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__8872\,
            I => \N__8865\
        );

    \I__1970\ : InMux
    port map (
            O => \N__8871\,
            I => \N__8862\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__8868\,
            I => \N__8856\
        );

    \I__1968\ : Span4Mux_v
    port map (
            O => \N__8865\,
            I => \N__8856\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__8862\,
            I => \N__8853\
        );

    \I__1966\ : CascadeMux
    port map (
            O => \N__8861\,
            I => \N__8850\
        );

    \I__1965\ : Span4Mux_v
    port map (
            O => \N__8856\,
            I => \N__8847\
        );

    \I__1964\ : Span12Mux_h
    port map (
            O => \N__8853\,
            I => \N__8844\
        );

    \I__1963\ : InMux
    port map (
            O => \N__8850\,
            I => \N__8841\
        );

    \I__1962\ : Odrv4
    port map (
            O => \N__8847\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1961\ : Odrv12
    port map (
            O => \N__8844\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__8841\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1959\ : IoInMux
    port map (
            O => \N__8834\,
            I => \N__8831\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__8831\,
            I => \N__8828\
        );

    \I__1957\ : Span12Mux_s10_v
    port map (
            O => \N__8828\,
            I => \N__8825\
        );

    \I__1956\ : Odrv12
    port map (
            O => \N__8825\,
            I => \CMA_c_10\
        );

    \I__1955\ : InMux
    port map (
            O => \N__8822\,
            I => \N__8819\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__8819\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\
        );

    \I__1953\ : InMux
    port map (
            O => \N__8816\,
            I => \N__8813\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__8813\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\
        );

    \I__1951\ : InMux
    port map (
            O => \N__8810\,
            I => \N__8807\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__8807\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\
        );

    \I__1949\ : IoInMux
    port map (
            O => \N__8804\,
            I => \N__8801\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__8801\,
            I => \N__8798\
        );

    \I__1947\ : IoSpan4Mux
    port map (
            O => \N__8798\,
            I => \N__8795\
        );

    \I__1946\ : Span4Mux_s2_h
    port map (
            O => \N__8795\,
            I => \N__8792\
        );

    \I__1945\ : Sp12to4
    port map (
            O => \N__8792\,
            I => \N__8789\
        );

    \I__1944\ : Span12Mux_h
    port map (
            O => \N__8789\,
            I => \N__8786\
        );

    \I__1943\ : Odrv12
    port map (
            O => \N__8786\,
            I => \CMA_c_5\
        );

    \I__1942\ : CascadeMux
    port map (
            O => \N__8783\,
            I => \N__8778\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__8782\,
            I => \N__8775\
        );

    \I__1940\ : CascadeMux
    port map (
            O => \N__8781\,
            I => \N__8772\
        );

    \I__1939\ : InMux
    port map (
            O => \N__8778\,
            I => \N__8767\
        );

    \I__1938\ : InMux
    port map (
            O => \N__8775\,
            I => \N__8763\
        );

    \I__1937\ : InMux
    port map (
            O => \N__8772\,
            I => \N__8760\
        );

    \I__1936\ : InMux
    port map (
            O => \N__8771\,
            I => \N__8752\
        );

    \I__1935\ : InMux
    port map (
            O => \N__8770\,
            I => \N__8752\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__8767\,
            I => \N__8749\
        );

    \I__1933\ : InMux
    port map (
            O => \N__8766\,
            I => \N__8746\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__8763\,
            I => \N__8743\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__8760\,
            I => \N__8740\
        );

    \I__1930\ : InMux
    port map (
            O => \N__8759\,
            I => \N__8733\
        );

    \I__1929\ : InMux
    port map (
            O => \N__8758\,
            I => \N__8733\
        );

    \I__1928\ : InMux
    port map (
            O => \N__8757\,
            I => \N__8733\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__8752\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1926\ : Odrv4
    port map (
            O => \N__8749\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__8746\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1924\ : Odrv4
    port map (
            O => \N__8743\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1923\ : Odrv4
    port map (
            O => \N__8740\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__8733\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1921\ : InMux
    port map (
            O => \N__8720\,
            I => \N__8712\
        );

    \I__1920\ : InMux
    port map (
            O => \N__8719\,
            I => \N__8707\
        );

    \I__1919\ : InMux
    port map (
            O => \N__8718\,
            I => \N__8707\
        );

    \I__1918\ : InMux
    port map (
            O => \N__8717\,
            I => \N__8704\
        );

    \I__1917\ : InMux
    port map (
            O => \N__8716\,
            I => \N__8699\
        );

    \I__1916\ : InMux
    port map (
            O => \N__8715\,
            I => \N__8699\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__8712\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__8707\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__8704\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__8699\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__1911\ : IoInMux
    port map (
            O => \N__8690\,
            I => \N__8687\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__8687\,
            I => \N__8684\
        );

    \I__1909\ : Span4Mux_s3_h
    port map (
            O => \N__8684\,
            I => \N__8681\
        );

    \I__1908\ : Sp12to4
    port map (
            O => \N__8681\,
            I => \N__8678\
        );

    \I__1907\ : Span12Mux_s9_v
    port map (
            O => \N__8678\,
            I => \N__8675\
        );

    \I__1906\ : Span12Mux_h
    port map (
            O => \N__8675\,
            I => \N__8672\
        );

    \I__1905\ : Odrv12
    port map (
            O => \N__8672\,
            I => \CMA_c_4\
        );

    \I__1904\ : InMux
    port map (
            O => \N__8669\,
            I => \N__8666\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__8666\,
            I => \N__8663\
        );

    \I__1902\ : Span4Mux_v
    port map (
            O => \N__8663\,
            I => \N__8660\
        );

    \I__1901\ : Span4Mux_v
    port map (
            O => \N__8660\,
            I => \N__8657\
        );

    \I__1900\ : Sp12to4
    port map (
            O => \N__8657\,
            I => \N__8654\
        );

    \I__1899\ : Span12Mux_h
    port map (
            O => \N__8654\,
            I => \N__8651\
        );

    \I__1898\ : Odrv12
    port map (
            O => \N__8651\,
            I => \A_c_19\
        );

    \I__1897\ : IoInMux
    port map (
            O => \N__8648\,
            I => \N__8645\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__8645\,
            I => \N__8642\
        );

    \I__1895\ : IoSpan4Mux
    port map (
            O => \N__8642\,
            I => \N__8639\
        );

    \I__1894\ : Span4Mux_s2_h
    port map (
            O => \N__8639\,
            I => \N__8636\
        );

    \I__1893\ : Sp12to4
    port map (
            O => \N__8636\,
            I => \N__8633\
        );

    \I__1892\ : Span12Mux_h
    port map (
            O => \N__8633\,
            I => \N__8630\
        );

    \I__1891\ : Odrv12
    port map (
            O => \N__8630\,
            I => \CMA_c_9\
        );

    \I__1890\ : CascadeMux
    port map (
            O => \N__8627\,
            I => \N__8624\
        );

    \I__1889\ : InMux
    port map (
            O => \N__8624\,
            I => \N__8621\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__8621\,
            I => \N__8618\
        );

    \I__1887\ : Span4Mux_h
    port map (
            O => \N__8618\,
            I => \N__8615\
        );

    \I__1886\ : Sp12to4
    port map (
            O => \N__8615\,
            I => \N__8612\
        );

    \I__1885\ : Span12Mux_v
    port map (
            O => \N__8612\,
            I => \N__8609\
        );

    \I__1884\ : Span12Mux_h
    port map (
            O => \N__8609\,
            I => \N__8606\
        );

    \I__1883\ : Odrv12
    port map (
            O => \N__8606\,
            I => \A_c_17\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__8603\,
            I => \N__8598\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__8602\,
            I => \N__8595\
        );

    \I__1880\ : InMux
    port map (
            O => \N__8601\,
            I => \N__8590\
        );

    \I__1879\ : InMux
    port map (
            O => \N__8598\,
            I => \N__8590\
        );

    \I__1878\ : InMux
    port map (
            O => \N__8595\,
            I => \N__8587\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8590\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__8587\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1875\ : IoInMux
    port map (
            O => \N__8582\,
            I => \N__8579\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__8579\,
            I => \N__8576\
        );

    \I__1873\ : Span4Mux_s3_h
    port map (
            O => \N__8576\,
            I => \N__8573\
        );

    \I__1872\ : Sp12to4
    port map (
            O => \N__8573\,
            I => \N__8570\
        );

    \I__1871\ : Span12Mux_v
    port map (
            O => \N__8570\,
            I => \N__8567\
        );

    \I__1870\ : Span12Mux_h
    port map (
            O => \N__8567\,
            I => \N__8564\
        );

    \I__1869\ : Odrv12
    port map (
            O => \N__8564\,
            I => \CMA_c_8\
        );

    \I__1868\ : InMux
    port map (
            O => \N__8561\,
            I => \N__8558\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__8558\,
            I => \N__8555\
        );

    \I__1866\ : Span4Mux_v
    port map (
            O => \N__8555\,
            I => \N__8552\
        );

    \I__1865\ : Sp12to4
    port map (
            O => \N__8552\,
            I => \N__8549\
        );

    \I__1864\ : Span12Mux_h
    port map (
            O => \N__8549\,
            I => \N__8546\
        );

    \I__1863\ : Span12Mux_v
    port map (
            O => \N__8546\,
            I => \N__8543\
        );

    \I__1862\ : Odrv12
    port map (
            O => \N__8543\,
            I => \A_c_3\
        );

    \I__1861\ : InMux
    port map (
            O => \N__8540\,
            I => \N__8537\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__8537\,
            I => \N__8534\
        );

    \I__1859\ : Span12Mux_h
    port map (
            O => \N__8534\,
            I => \N__8531\
        );

    \I__1858\ : Odrv12
    port map (
            O => \N__8531\,
            I => \A_c_10\
        );

    \I__1857\ : CascadeMux
    port map (
            O => \N__8528\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\
        );

    \I__1856\ : InMux
    port map (
            O => \N__8525\,
            I => \N__8519\
        );

    \I__1855\ : InMux
    port map (
            O => \N__8524\,
            I => \N__8519\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__8519\,
            I => \N__8516\
        );

    \I__1853\ : Odrv4
    port map (
            O => \N__8516\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__1852\ : InMux
    port map (
            O => \N__8513\,
            I => \N__8510\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__8510\,
            I => \N__8507\
        );

    \I__1850\ : Span4Mux_h
    port map (
            O => \N__8507\,
            I => \N__8504\
        );

    \I__1849\ : Odrv4
    port map (
            O => \N__8504\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__1848\ : InMux
    port map (
            O => \N__8501\,
            I => \N__8498\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__8498\,
            I => \N__8495\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__8495\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1845\ : InMux
    port map (
            O => \N__8492\,
            I => \N__8489\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__8489\,
            I => \N__8486\
        );

    \I__1843\ : Odrv4
    port map (
            O => \N__8486\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__8483\,
            I => \N__8478\
        );

    \I__1841\ : CascadeMux
    port map (
            O => \N__8482\,
            I => \N__8475\
        );

    \I__1840\ : InMux
    port map (
            O => \N__8481\,
            I => \N__8467\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8478\,
            I => \N__8467\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8475\,
            I => \N__8467\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8474\,
            I => \N__8464\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__8467\,
            I => \N__8461\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__8464\,
            I => \N__8458\
        );

    \I__1834\ : Span4Mux_v
    port map (
            O => \N__8461\,
            I => \N__8455\
        );

    \I__1833\ : Span4Mux_v
    port map (
            O => \N__8458\,
            I => \N__8450\
        );

    \I__1832\ : Span4Mux_h
    port map (
            O => \N__8455\,
            I => \N__8450\
        );

    \I__1831\ : Span4Mux_v
    port map (
            O => \N__8450\,
            I => \N__8447\
        );

    \I__1830\ : Span4Mux_v
    port map (
            O => \N__8447\,
            I => \N__8444\
        );

    \I__1829\ : Odrv4
    port map (
            O => \N__8444\,
            I => \CLK40_PLL_i\
        );

    \I__1828\ : IoInMux
    port map (
            O => \N__8441\,
            I => \N__8437\
        );

    \I__1827\ : IoInMux
    port map (
            O => \N__8440\,
            I => \N__8434\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__8437\,
            I => \N__8431\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__8434\,
            I => \N__8428\
        );

    \I__1824\ : Span4Mux_s0_v
    port map (
            O => \N__8431\,
            I => \N__8425\
        );

    \I__1823\ : Span4Mux_s0_v
    port map (
            O => \N__8428\,
            I => \N__8422\
        );

    \I__1822\ : Span4Mux_v
    port map (
            O => \N__8425\,
            I => \N__8419\
        );

    \I__1821\ : Span4Mux_v
    port map (
            O => \N__8422\,
            I => \N__8416\
        );

    \I__1820\ : Sp12to4
    port map (
            O => \N__8419\,
            I => \N__8410\
        );

    \I__1819\ : Sp12to4
    port map (
            O => \N__8416\,
            I => \N__8410\
        );

    \I__1818\ : IoInMux
    port map (
            O => \N__8415\,
            I => \N__8407\
        );

    \I__1817\ : Span12Mux_h
    port map (
            O => \N__8410\,
            I => \N__8404\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__8407\,
            I => \N__8401\
        );

    \I__1815\ : Span12Mux_v
    port map (
            O => \N__8404\,
            I => \N__8396\
        );

    \I__1814\ : Span12Mux_s5_h
    port map (
            O => \N__8401\,
            I => \N__8396\
        );

    \I__1813\ : Odrv12
    port map (
            O => \N__8396\,
            I => \CLK40_PLL_i_i\
        );

    \I__1812\ : InMux
    port map (
            O => \N__8393\,
            I => \N__8383\
        );

    \I__1811\ : InMux
    port map (
            O => \N__8392\,
            I => \N__8376\
        );

    \I__1810\ : InMux
    port map (
            O => \N__8391\,
            I => \N__8376\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8390\,
            I => \N__8376\
        );

    \I__1808\ : InMux
    port map (
            O => \N__8389\,
            I => \N__8365\
        );

    \I__1807\ : InMux
    port map (
            O => \N__8388\,
            I => \N__8365\
        );

    \I__1806\ : InMux
    port map (
            O => \N__8387\,
            I => \N__8365\
        );

    \I__1805\ : InMux
    port map (
            O => \N__8386\,
            I => \N__8356\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__8383\,
            I => \N__8353\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__8376\,
            I => \N__8350\
        );

    \I__1802\ : InMux
    port map (
            O => \N__8375\,
            I => \N__8345\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8374\,
            I => \N__8345\
        );

    \I__1800\ : InMux
    port map (
            O => \N__8373\,
            I => \N__8342\
        );

    \I__1799\ : InMux
    port map (
            O => \N__8372\,
            I => \N__8339\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__8365\,
            I => \N__8336\
        );

    \I__1797\ : InMux
    port map (
            O => \N__8364\,
            I => \N__8329\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8363\,
            I => \N__8329\
        );

    \I__1795\ : InMux
    port map (
            O => \N__8362\,
            I => \N__8329\
        );

    \I__1794\ : InMux
    port map (
            O => \N__8361\,
            I => \N__8326\
        );

    \I__1793\ : InMux
    port map (
            O => \N__8360\,
            I => \N__8321\
        );

    \I__1792\ : InMux
    port map (
            O => \N__8359\,
            I => \N__8321\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__8356\,
            I => \N__8318\
        );

    \I__1790\ : Span4Mux_v
    port map (
            O => \N__8353\,
            I => \N__8315\
        );

    \I__1789\ : Span4Mux_v
    port map (
            O => \N__8350\,
            I => \N__8308\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__8345\,
            I => \N__8308\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__8342\,
            I => \N__8308\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__8339\,
            I => \N__8305\
        );

    \I__1785\ : Span4Mux_h
    port map (
            O => \N__8336\,
            I => \N__8296\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__8329\,
            I => \N__8296\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__8326\,
            I => \N__8296\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__8321\,
            I => \N__8296\
        );

    \I__1781\ : Sp12to4
    port map (
            O => \N__8318\,
            I => \N__8292\
        );

    \I__1780\ : Span4Mux_v
    port map (
            O => \N__8315\,
            I => \N__8287\
        );

    \I__1779\ : Span4Mux_v
    port map (
            O => \N__8308\,
            I => \N__8287\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__8305\,
            I => \N__8282\
        );

    \I__1777\ : Span4Mux_v
    port map (
            O => \N__8296\,
            I => \N__8282\
        );

    \I__1776\ : InMux
    port map (
            O => \N__8295\,
            I => \N__8279\
        );

    \I__1775\ : Span12Mux_v
    port map (
            O => \N__8292\,
            I => \N__8270\
        );

    \I__1774\ : Sp12to4
    port map (
            O => \N__8287\,
            I => \N__8270\
        );

    \I__1773\ : Sp12to4
    port map (
            O => \N__8282\,
            I => \N__8270\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__8279\,
            I => \N__8270\
        );

    \I__1771\ : Span12Mux_h
    port map (
            O => \N__8270\,
            I => \N__8267\
        );

    \I__1770\ : Odrv12
    port map (
            O => \N__8267\,
            I => \RESETn_c\
        );

    \I__1769\ : IoInMux
    port map (
            O => \N__8264\,
            I => \N__8261\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__8261\,
            I => \N__8258\
        );

    \I__1767\ : Span12Mux_s1_v
    port map (
            O => \N__8258\,
            I => \N__8255\
        );

    \I__1766\ : Odrv12
    port map (
            O => \N__8255\,
            I => \RESETn_c_i\
        );

    \I__1765\ : InMux
    port map (
            O => \N__8252\,
            I => \N__8245\
        );

    \I__1764\ : InMux
    port map (
            O => \N__8251\,
            I => \N__8245\
        );

    \I__1763\ : InMux
    port map (
            O => \N__8250\,
            I => \N__8242\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__8245\,
            I => \N__8236\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__8242\,
            I => \N__8236\
        );

    \I__1760\ : CascadeMux
    port map (
            O => \N__8241\,
            I => \N__8233\
        );

    \I__1759\ : Span4Mux_v
    port map (
            O => \N__8236\,
            I => \N__8229\
        );

    \I__1758\ : InMux
    port map (
            O => \N__8233\,
            I => \N__8226\
        );

    \I__1757\ : InMux
    port map (
            O => \N__8232\,
            I => \N__8223\
        );

    \I__1756\ : Span4Mux_v
    port map (
            O => \N__8229\,
            I => \N__8216\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__8226\,
            I => \N__8216\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__8223\,
            I => \N__8216\
        );

    \I__1753\ : Span4Mux_v
    port map (
            O => \N__8216\,
            I => \N__8212\
        );

    \I__1752\ : InMux
    port map (
            O => \N__8215\,
            I => \N__8209\
        );

    \I__1751\ : Span4Mux_v
    port map (
            O => \N__8212\,
            I => \N__8206\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__8209\,
            I => \N__8203\
        );

    \I__1749\ : Sp12to4
    port map (
            O => \N__8206\,
            I => \N__8198\
        );

    \I__1748\ : Span12Mux_v
    port map (
            O => \N__8203\,
            I => \N__8198\
        );

    \I__1747\ : Span12Mux_h
    port map (
            O => \N__8198\,
            I => \N__8195\
        );

    \I__1746\ : Odrv12
    port map (
            O => \N__8195\,
            I => \CASLn_c\
        );

    \I__1745\ : InMux
    port map (
            O => \N__8192\,
            I => \N__8184\
        );

    \I__1744\ : InMux
    port map (
            O => \N__8191\,
            I => \N__8184\
        );

    \I__1743\ : InMux
    port map (
            O => \N__8190\,
            I => \N__8181\
        );

    \I__1742\ : InMux
    port map (
            O => \N__8189\,
            I => \N__8178\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__8184\,
            I => \N__8173\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__8181\,
            I => \N__8173\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__8178\,
            I => \N__8168\
        );

    \I__1738\ : Span4Mux_v
    port map (
            O => \N__8173\,
            I => \N__8165\
        );

    \I__1737\ : InMux
    port map (
            O => \N__8172\,
            I => \N__8160\
        );

    \I__1736\ : InMux
    port map (
            O => \N__8171\,
            I => \N__8160\
        );

    \I__1735\ : Span4Mux_v
    port map (
            O => \N__8168\,
            I => \N__8157\
        );

    \I__1734\ : Sp12to4
    port map (
            O => \N__8165\,
            I => \N__8154\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__8160\,
            I => \N__8151\
        );

    \I__1732\ : Span4Mux_v
    port map (
            O => \N__8157\,
            I => \N__8148\
        );

    \I__1731\ : Span12Mux_h
    port map (
            O => \N__8154\,
            I => \N__8145\
        );

    \I__1730\ : Span12Mux_v
    port map (
            O => \N__8151\,
            I => \N__8142\
        );

    \I__1729\ : Sp12to4
    port map (
            O => \N__8148\,
            I => \N__8139\
        );

    \I__1728\ : Span12Mux_v
    port map (
            O => \N__8145\,
            I => \N__8134\
        );

    \I__1727\ : Span12Mux_h
    port map (
            O => \N__8142\,
            I => \N__8134\
        );

    \I__1726\ : Span12Mux_h
    port map (
            O => \N__8139\,
            I => \N__8131\
        );

    \I__1725\ : Odrv12
    port map (
            O => \N__8134\,
            I => \CASUn_c\
        );

    \I__1724\ : Odrv12
    port map (
            O => \N__8131\,
            I => \CASUn_c\
        );

    \I__1723\ : InMux
    port map (
            O => \N__8126\,
            I => \N__8121\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8125\,
            I => \N__8118\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8124\,
            I => \N__8115\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__8121\,
            I => \N__8112\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__8118\,
            I => \N__8109\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__8115\,
            I => \N__8106\
        );

    \I__1717\ : Span4Mux_h
    port map (
            O => \N__8112\,
            I => \N__8103\
        );

    \I__1716\ : Span12Mux_h
    port map (
            O => \N__8109\,
            I => \N__8100\
        );

    \I__1715\ : Span4Mux_v
    port map (
            O => \N__8106\,
            I => \N__8097\
        );

    \I__1714\ : Span4Mux_v
    port map (
            O => \N__8103\,
            I => \N__8094\
        );

    \I__1713\ : Span12Mux_v
    port map (
            O => \N__8100\,
            I => \N__8091\
        );

    \I__1712\ : Span4Mux_h
    port map (
            O => \N__8097\,
            I => \N__8088\
        );

    \I__1711\ : Span4Mux_v
    port map (
            O => \N__8094\,
            I => \N__8085\
        );

    \I__1710\ : Odrv12
    port map (
            O => \N__8091\,
            I => \REG_CYCLEm\
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__8088\,
            I => \REG_CYCLEm\
        );

    \I__1708\ : Odrv4
    port map (
            O => \N__8085\,
            I => \REG_CYCLEm\
        );

    \I__1707\ : IoInMux
    port map (
            O => \N__8078\,
            I => \N__8075\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__8075\,
            I => \N__8072\
        );

    \I__1705\ : Span4Mux_s1_v
    port map (
            O => \N__8072\,
            I => \N__8069\
        );

    \I__1704\ : Span4Mux_h
    port map (
            O => \N__8069\,
            I => \N__8066\
        );

    \I__1703\ : Sp12to4
    port map (
            O => \N__8066\,
            I => \N__8063\
        );

    \I__1702\ : Span12Mux_h
    port map (
            O => \N__8063\,
            I => \N__8060\
        );

    \I__1701\ : Odrv12
    port map (
            O => \N__8060\,
            I => \DRDENn_c\
        );

    \I__1700\ : IoInMux
    port map (
            O => \N__8057\,
            I => \N__8054\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__8054\,
            I => \N__8051\
        );

    \I__1698\ : Span4Mux_s3_v
    port map (
            O => \N__8051\,
            I => \N__8048\
        );

    \I__1697\ : Span4Mux_v
    port map (
            O => \N__8048\,
            I => \N__8045\
        );

    \I__1696\ : Span4Mux_h
    port map (
            O => \N__8045\,
            I => \N__8042\
        );

    \I__1695\ : Odrv4
    port map (
            O => \N__8042\,
            I => \CRCSn_c\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8039\,
            I => \N__8036\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__8036\,
            I => \N__8033\
        );

    \I__1692\ : Span4Mux_v
    port map (
            O => \N__8033\,
            I => \N__8030\
        );

    \I__1691\ : Span4Mux_h
    port map (
            O => \N__8030\,
            I => \N__8027\
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__8027\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1689\ : IoInMux
    port map (
            O => \N__8024\,
            I => \N__8021\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__8021\,
            I => \N__8018\
        );

    \I__1687\ : IoSpan4Mux
    port map (
            O => \N__8018\,
            I => \N__8015\
        );

    \I__1686\ : Span4Mux_s1_h
    port map (
            O => \N__8015\,
            I => \N__8012\
        );

    \I__1685\ : Sp12to4
    port map (
            O => \N__8012\,
            I => \N__8009\
        );

    \I__1684\ : Span12Mux_h
    port map (
            O => \N__8009\,
            I => \N__8006\
        );

    \I__1683\ : Odrv12
    port map (
            O => \N__8006\,
            I => \CMA_c_3\
        );

    \I__1682\ : InMux
    port map (
            O => \N__8003\,
            I => \N__8000\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__8000\,
            I => \N__7997\
        );

    \I__1680\ : Span4Mux_v
    port map (
            O => \N__7997\,
            I => \N__7994\
        );

    \I__1679\ : Span4Mux_v
    port map (
            O => \N__7994\,
            I => \N__7991\
        );

    \I__1678\ : Sp12to4
    port map (
            O => \N__7991\,
            I => \N__7988\
        );

    \I__1677\ : Span12Mux_h
    port map (
            O => \N__7988\,
            I => \N__7985\
        );

    \I__1676\ : Odrv12
    port map (
            O => \N__7985\,
            I => \A_c_7\
        );

    \I__1675\ : CascadeMux
    port map (
            O => \N__7982\,
            I => \U712_CHIP_RAM.N_463_cascade_\
        );

    \I__1674\ : InMux
    port map (
            O => \N__7979\,
            I => \N__7976\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__7976\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i\
        );

    \I__1672\ : InMux
    port map (
            O => \N__7973\,
            I => \N__7958\
        );

    \I__1671\ : InMux
    port map (
            O => \N__7972\,
            I => \N__7958\
        );

    \I__1670\ : InMux
    port map (
            O => \N__7971\,
            I => \N__7958\
        );

    \I__1669\ : InMux
    port map (
            O => \N__7970\,
            I => \N__7955\
        );

    \I__1668\ : InMux
    port map (
            O => \N__7969\,
            I => \N__7952\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__7968\,
            I => \N__7946\
        );

    \I__1666\ : CascadeMux
    port map (
            O => \N__7967\,
            I => \N__7942\
        );

    \I__1665\ : InMux
    port map (
            O => \N__7966\,
            I => \N__7937\
        );

    \I__1664\ : InMux
    port map (
            O => \N__7965\,
            I => \N__7937\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__7958\,
            I => \N__7934\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__7955\,
            I => \N__7929\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__7952\,
            I => \N__7929\
        );

    \I__1660\ : InMux
    port map (
            O => \N__7951\,
            I => \N__7924\
        );

    \I__1659\ : InMux
    port map (
            O => \N__7950\,
            I => \N__7924\
        );

    \I__1658\ : InMux
    port map (
            O => \N__7949\,
            I => \N__7918\
        );

    \I__1657\ : InMux
    port map (
            O => \N__7946\,
            I => \N__7915\
        );

    \I__1656\ : InMux
    port map (
            O => \N__7945\,
            I => \N__7910\
        );

    \I__1655\ : InMux
    port map (
            O => \N__7942\,
            I => \N__7910\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__7937\,
            I => \N__7907\
        );

    \I__1653\ : Span4Mux_h
    port map (
            O => \N__7934\,
            I => \N__7904\
        );

    \I__1652\ : Span4Mux_v
    port map (
            O => \N__7929\,
            I => \N__7899\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__7924\,
            I => \N__7899\
        );

    \I__1650\ : InMux
    port map (
            O => \N__7923\,
            I => \N__7896\
        );

    \I__1649\ : InMux
    port map (
            O => \N__7922\,
            I => \N__7893\
        );

    \I__1648\ : InMux
    port map (
            O => \N__7921\,
            I => \N__7890\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__7918\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__7915\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__7910\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1644\ : Odrv4
    port map (
            O => \N__7907\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1643\ : Odrv4
    port map (
            O => \N__7904\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1642\ : Odrv4
    port map (
            O => \N__7899\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__7896\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__7893\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__7890\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1638\ : InMux
    port map (
            O => \N__7871\,
            I => \N__7864\
        );

    \I__1637\ : InMux
    port map (
            O => \N__7870\,
            I => \N__7861\
        );

    \I__1636\ : InMux
    port map (
            O => \N__7869\,
            I => \N__7858\
        );

    \I__1635\ : InMux
    port map (
            O => \N__7868\,
            I => \N__7855\
        );

    \I__1634\ : CascadeMux
    port map (
            O => \N__7867\,
            I => \N__7852\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__7864\,
            I => \N__7841\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__7861\,
            I => \N__7841\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__7858\,
            I => \N__7836\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__7855\,
            I => \N__7836\
        );

    \I__1629\ : InMux
    port map (
            O => \N__7852\,
            I => \N__7833\
        );

    \I__1628\ : InMux
    port map (
            O => \N__7851\,
            I => \N__7829\
        );

    \I__1627\ : InMux
    port map (
            O => \N__7850\,
            I => \N__7826\
        );

    \I__1626\ : InMux
    port map (
            O => \N__7849\,
            I => \N__7823\
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__7848\,
            I => \N__7820\
        );

    \I__1624\ : CascadeMux
    port map (
            O => \N__7847\,
            I => \N__7816\
        );

    \I__1623\ : InMux
    port map (
            O => \N__7846\,
            I => \N__7805\
        );

    \I__1622\ : Span4Mux_v
    port map (
            O => \N__7841\,
            I => \N__7802\
        );

    \I__1621\ : Span4Mux_v
    port map (
            O => \N__7836\,
            I => \N__7797\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__7833\,
            I => \N__7797\
        );

    \I__1619\ : InMux
    port map (
            O => \N__7832\,
            I => \N__7794\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__7829\,
            I => \N__7787\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__7826\,
            I => \N__7787\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__7823\,
            I => \N__7787\
        );

    \I__1615\ : InMux
    port map (
            O => \N__7820\,
            I => \N__7778\
        );

    \I__1614\ : InMux
    port map (
            O => \N__7819\,
            I => \N__7778\
        );

    \I__1613\ : InMux
    port map (
            O => \N__7816\,
            I => \N__7778\
        );

    \I__1612\ : InMux
    port map (
            O => \N__7815\,
            I => \N__7778\
        );

    \I__1611\ : InMux
    port map (
            O => \N__7814\,
            I => \N__7775\
        );

    \I__1610\ : InMux
    port map (
            O => \N__7813\,
            I => \N__7762\
        );

    \I__1609\ : InMux
    port map (
            O => \N__7812\,
            I => \N__7762\
        );

    \I__1608\ : InMux
    port map (
            O => \N__7811\,
            I => \N__7762\
        );

    \I__1607\ : InMux
    port map (
            O => \N__7810\,
            I => \N__7762\
        );

    \I__1606\ : InMux
    port map (
            O => \N__7809\,
            I => \N__7762\
        );

    \I__1605\ : InMux
    port map (
            O => \N__7808\,
            I => \N__7762\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__7805\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1603\ : Odrv4
    port map (
            O => \N__7802\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1602\ : Odrv4
    port map (
            O => \N__7797\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__7794\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1600\ : Odrv4
    port map (
            O => \N__7787\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__7778\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__7775\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__7762\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1596\ : InMux
    port map (
            O => \N__7745\,
            I => \N__7742\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__7742\,
            I => \N__7737\
        );

    \I__1594\ : InMux
    port map (
            O => \N__7741\,
            I => \N__7734\
        );

    \I__1593\ : InMux
    port map (
            O => \N__7740\,
            I => \N__7731\
        );

    \I__1592\ : Span4Mux_v
    port map (
            O => \N__7737\,
            I => \N__7726\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__7734\,
            I => \N__7726\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__7731\,
            I => \N__7723\
        );

    \I__1589\ : Span4Mux_h
    port map (
            O => \N__7726\,
            I => \N__7720\
        );

    \I__1588\ : Odrv12
    port map (
            O => \N__7723\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRTZ0Z_2\
        );

    \I__1587\ : Odrv4
    port map (
            O => \N__7720\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRTZ0Z_2\
        );

    \I__1586\ : InMux
    port map (
            O => \N__7715\,
            I => \N__7712\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__7712\,
            I => \N__7709\
        );

    \I__1584\ : Odrv4
    port map (
            O => \N__7709\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__1583\ : InMux
    port map (
            O => \N__7706\,
            I => \N__7703\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__7703\,
            I => \N__7700\
        );

    \I__1581\ : Odrv12
    port map (
            O => \N__7700\,
            I => \U712_CHIP_RAM.un3_DMA_CYCLE_START\
        );

    \I__1580\ : InMux
    port map (
            O => \N__7697\,
            I => \N__7691\
        );

    \I__1579\ : InMux
    port map (
            O => \N__7696\,
            I => \N__7691\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__7691\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1577\ : InMux
    port map (
            O => \N__7688\,
            I => \N__7685\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__7685\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1575\ : InMux
    port map (
            O => \N__7682\,
            I => \N__7679\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__7679\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__1573\ : IoInMux
    port map (
            O => \N__7676\,
            I => \N__7673\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__7673\,
            I => \N__7670\
        );

    \I__1571\ : Span4Mux_s1_v
    port map (
            O => \N__7670\,
            I => \N__7667\
        );

    \I__1570\ : Span4Mux_v
    port map (
            O => \N__7667\,
            I => \N__7664\
        );

    \I__1569\ : Span4Mux_v
    port map (
            O => \N__7664\,
            I => \N__7661\
        );

    \I__1568\ : Odrv4
    port map (
            O => \N__7661\,
            I => \CMA_c_2\
        );

    \I__1567\ : InMux
    port map (
            O => \N__7658\,
            I => \N__7655\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__7655\,
            I => \N__7652\
        );

    \I__1565\ : Span4Mux_h
    port map (
            O => \N__7652\,
            I => \N__7649\
        );

    \I__1564\ : Span4Mux_v
    port map (
            O => \N__7649\,
            I => \N__7646\
        );

    \I__1563\ : Odrv4
    port map (
            O => \N__7646\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__7643\,
            I => \U712_CHIP_RAM.CMA_5_0_8_cascade_\
        );

    \I__1561\ : InMux
    port map (
            O => \N__7640\,
            I => \N__7634\
        );

    \I__1560\ : InMux
    port map (
            O => \N__7639\,
            I => \N__7634\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__7634\,
            I => \N__7631\
        );

    \I__1558\ : Span4Mux_v
    port map (
            O => \N__7631\,
            I => \N__7628\
        );

    \I__1557\ : Span4Mux_v
    port map (
            O => \N__7628\,
            I => \N__7625\
        );

    \I__1556\ : Sp12to4
    port map (
            O => \N__7625\,
            I => \N__7622\
        );

    \I__1555\ : Span12Mux_h
    port map (
            O => \N__7622\,
            I => \N__7619\
        );

    \I__1554\ : Odrv12
    port map (
            O => \N__7619\,
            I => \A_c_14\
        );

    \I__1553\ : CascadeMux
    port map (
            O => \N__7616\,
            I => \N__7613\
        );

    \I__1552\ : InMux
    port map (
            O => \N__7613\,
            I => \N__7606\
        );

    \I__1551\ : InMux
    port map (
            O => \N__7612\,
            I => \N__7596\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7611\,
            I => \N__7596\
        );

    \I__1549\ : InMux
    port map (
            O => \N__7610\,
            I => \N__7596\
        );

    \I__1548\ : InMux
    port map (
            O => \N__7609\,
            I => \N__7596\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__7606\,
            I => \N__7593\
        );

    \I__1546\ : InMux
    port map (
            O => \N__7605\,
            I => \N__7590\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__7596\,
            I => \N__7585\
        );

    \I__1544\ : Span4Mux_v
    port map (
            O => \N__7593\,
            I => \N__7580\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__7590\,
            I => \N__7580\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7589\,
            I => \N__7575\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7588\,
            I => \N__7575\
        );

    \I__1540\ : Odrv12
    port map (
            O => \N__7585\,
            I => \DMA_CYCLEm\
        );

    \I__1539\ : Odrv4
    port map (
            O => \N__7580\,
            I => \DMA_CYCLEm\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7575\,
            I => \DMA_CYCLEm\
        );

    \I__1537\ : InMux
    port map (
            O => \N__7568\,
            I => \N__7563\
        );

    \I__1536\ : CascadeMux
    port map (
            O => \N__7567\,
            I => \N__7559\
        );

    \I__1535\ : CascadeMux
    port map (
            O => \N__7566\,
            I => \N__7556\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__7563\,
            I => \N__7553\
        );

    \I__1533\ : InMux
    port map (
            O => \N__7562\,
            I => \N__7550\
        );

    \I__1532\ : InMux
    port map (
            O => \N__7559\,
            I => \N__7547\
        );

    \I__1531\ : InMux
    port map (
            O => \N__7556\,
            I => \N__7542\
        );

    \I__1530\ : Span4Mux_v
    port map (
            O => \N__7553\,
            I => \N__7537\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__7550\,
            I => \N__7537\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__7547\,
            I => \N__7534\
        );

    \I__1527\ : InMux
    port map (
            O => \N__7546\,
            I => \N__7531\
        );

    \I__1526\ : InMux
    port map (
            O => \N__7545\,
            I => \N__7528\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__7542\,
            I => \N__7525\
        );

    \I__1524\ : Span4Mux_v
    port map (
            O => \N__7537\,
            I => \N__7522\
        );

    \I__1523\ : Span4Mux_h
    port map (
            O => \N__7534\,
            I => \N__7518\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7531\,
            I => \N__7513\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__7528\,
            I => \N__7513\
        );

    \I__1520\ : Span4Mux_h
    port map (
            O => \N__7525\,
            I => \N__7507\
        );

    \I__1519\ : Span4Mux_h
    port map (
            O => \N__7522\,
            I => \N__7504\
        );

    \I__1518\ : InMux
    port map (
            O => \N__7521\,
            I => \N__7501\
        );

    \I__1517\ : Span4Mux_h
    port map (
            O => \N__7518\,
            I => \N__7496\
        );

    \I__1516\ : Span4Mux_h
    port map (
            O => \N__7513\,
            I => \N__7496\
        );

    \I__1515\ : InMux
    port map (
            O => \N__7512\,
            I => \N__7491\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7511\,
            I => \N__7491\
        );

    \I__1513\ : InMux
    port map (
            O => \N__7510\,
            I => \N__7488\
        );

    \I__1512\ : Odrv4
    port map (
            O => \N__7507\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1511\ : Odrv4
    port map (
            O => \N__7504\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__7501\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1509\ : Odrv4
    port map (
            O => \N__7496\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7491\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__7488\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7475\,
            I => \N__7472\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__7472\,
            I => \N__7469\
        );

    \I__1504\ : Span4Mux_v
    port map (
            O => \N__7469\,
            I => \N__7465\
        );

    \I__1503\ : InMux
    port map (
            O => \N__7468\,
            I => \N__7462\
        );

    \I__1502\ : Odrv4
    port map (
            O => \N__7465\,
            I => \U712_CHIP_RAM.N_201_i_i_a2_3_1\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__7462\,
            I => \U712_CHIP_RAM.N_201_i_i_a2_3_1\
        );

    \I__1500\ : SRMux
    port map (
            O => \N__7457\,
            I => \N__7454\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__7454\,
            I => \N__7451\
        );

    \I__1498\ : Span4Mux_h
    port map (
            O => \N__7451\,
            I => \N__7448\
        );

    \I__1497\ : Odrv4
    port map (
            O => \N__7448\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1496\ : CascadeMux
    port map (
            O => \N__7445\,
            I => \N__7440\
        );

    \I__1495\ : InMux
    port map (
            O => \N__7444\,
            I => \N__7429\
        );

    \I__1494\ : CascadeMux
    port map (
            O => \N__7443\,
            I => \N__7423\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7440\,
            I => \N__7420\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7439\,
            I => \N__7417\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7438\,
            I => \N__7410\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7437\,
            I => \N__7403\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7436\,
            I => \N__7403\
        );

    \I__1488\ : InMux
    port map (
            O => \N__7435\,
            I => \N__7403\
        );

    \I__1487\ : InMux
    port map (
            O => \N__7434\,
            I => \N__7396\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7433\,
            I => \N__7396\
        );

    \I__1485\ : InMux
    port map (
            O => \N__7432\,
            I => \N__7396\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__7429\,
            I => \N__7392\
        );

    \I__1483\ : InMux
    port map (
            O => \N__7428\,
            I => \N__7387\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7427\,
            I => \N__7387\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7426\,
            I => \N__7382\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7423\,
            I => \N__7375\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7420\,
            I => \N__7372\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__7417\,
            I => \N__7369\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7416\,
            I => \N__7360\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7415\,
            I => \N__7360\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7414\,
            I => \N__7360\
        );

    \I__1474\ : InMux
    port map (
            O => \N__7413\,
            I => \N__7360\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__7410\,
            I => \N__7353\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__7403\,
            I => \N__7353\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__7396\,
            I => \N__7353\
        );

    \I__1470\ : InMux
    port map (
            O => \N__7395\,
            I => \N__7350\
        );

    \I__1469\ : Span4Mux_v
    port map (
            O => \N__7392\,
            I => \N__7345\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__7387\,
            I => \N__7345\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7340\
        );

    \I__1466\ : InMux
    port map (
            O => \N__7385\,
            I => \N__7340\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__7382\,
            I => \N__7337\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7381\,
            I => \N__7334\
        );

    \I__1463\ : InMux
    port map (
            O => \N__7380\,
            I => \N__7327\
        );

    \I__1462\ : InMux
    port map (
            O => \N__7379\,
            I => \N__7327\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7378\,
            I => \N__7327\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__7375\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1459\ : Odrv12
    port map (
            O => \N__7372\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1458\ : Odrv4
    port map (
            O => \N__7369\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__7360\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1456\ : Odrv4
    port map (
            O => \N__7353\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__7350\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1454\ : Odrv4
    port map (
            O => \N__7345\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__7340\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1452\ : Odrv4
    port map (
            O => \N__7337\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__7334\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__7327\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1449\ : InMux
    port map (
            O => \N__7304\,
            I => \N__7298\
        );

    \I__1448\ : InMux
    port map (
            O => \N__7303\,
            I => \N__7298\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__7298\,
            I => \N__7295\
        );

    \I__1446\ : Span4Mux_v
    port map (
            O => \N__7295\,
            I => \N__7291\
        );

    \I__1445\ : InMux
    port map (
            O => \N__7294\,
            I => \N__7288\
        );

    \I__1444\ : Span4Mux_v
    port map (
            O => \N__7291\,
            I => \N__7279\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__7288\,
            I => \N__7279\
        );

    \I__1442\ : InMux
    port map (
            O => \N__7287\,
            I => \N__7276\
        );

    \I__1441\ : InMux
    port map (
            O => \N__7286\,
            I => \N__7273\
        );

    \I__1440\ : InMux
    port map (
            O => \N__7285\,
            I => \N__7270\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7284\,
            I => \N__7265\
        );

    \I__1438\ : Span4Mux_v
    port map (
            O => \N__7279\,
            I => \N__7256\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__7276\,
            I => \N__7256\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__7273\,
            I => \N__7256\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__7270\,
            I => \N__7256\
        );

    \I__1434\ : InMux
    port map (
            O => \N__7269\,
            I => \N__7251\
        );

    \I__1433\ : InMux
    port map (
            O => \N__7268\,
            I => \N__7251\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__7265\,
            I => \N__7248\
        );

    \I__1431\ : Span4Mux_v
    port map (
            O => \N__7256\,
            I => \N__7242\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__7251\,
            I => \N__7239\
        );

    \I__1429\ : Span4Mux_v
    port map (
            O => \N__7248\,
            I => \N__7236\
        );

    \I__1428\ : InMux
    port map (
            O => \N__7247\,
            I => \N__7229\
        );

    \I__1427\ : InMux
    port map (
            O => \N__7246\,
            I => \N__7229\
        );

    \I__1426\ : InMux
    port map (
            O => \N__7245\,
            I => \N__7229\
        );

    \I__1425\ : Odrv4
    port map (
            O => \N__7242\,
            I => \WRITE_CYCLEm\
        );

    \I__1424\ : Odrv4
    port map (
            O => \N__7239\,
            I => \WRITE_CYCLEm\
        );

    \I__1423\ : Odrv4
    port map (
            O => \N__7236\,
            I => \WRITE_CYCLEm\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__7229\,
            I => \WRITE_CYCLEm\
        );

    \I__1421\ : InMux
    port map (
            O => \N__7220\,
            I => \N__7214\
        );

    \I__1420\ : InMux
    port map (
            O => \N__7219\,
            I => \N__7211\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7218\,
            I => \N__7206\
        );

    \I__1418\ : InMux
    port map (
            O => \N__7217\,
            I => \N__7203\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__7214\,
            I => \N__7199\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__7211\,
            I => \N__7196\
        );

    \I__1415\ : InMux
    port map (
            O => \N__7210\,
            I => \N__7188\
        );

    \I__1414\ : InMux
    port map (
            O => \N__7209\,
            I => \N__7188\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__7206\,
            I => \N__7183\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__7203\,
            I => \N__7183\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7202\,
            I => \N__7180\
        );

    \I__1410\ : Span4Mux_h
    port map (
            O => \N__7199\,
            I => \N__7175\
        );

    \I__1409\ : Span4Mux_h
    port map (
            O => \N__7196\,
            I => \N__7175\
        );

    \I__1408\ : InMux
    port map (
            O => \N__7195\,
            I => \N__7168\
        );

    \I__1407\ : InMux
    port map (
            O => \N__7194\,
            I => \N__7168\
        );

    \I__1406\ : InMux
    port map (
            O => \N__7193\,
            I => \N__7168\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__7188\,
            I => \N__7161\
        );

    \I__1404\ : Span4Mux_v
    port map (
            O => \N__7183\,
            I => \N__7161\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__7180\,
            I => \N__7161\
        );

    \I__1402\ : Odrv4
    port map (
            O => \N__7175\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__7168\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1400\ : Odrv4
    port map (
            O => \N__7161\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__7154\,
            I => \U712_CHIP_RAM.N_306_cascade_\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7151\,
            I => \N__7147\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__7150\,
            I => \N__7139\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__7147\,
            I => \N__7135\
        );

    \I__1395\ : InMux
    port map (
            O => \N__7146\,
            I => \N__7132\
        );

    \I__1394\ : InMux
    port map (
            O => \N__7145\,
            I => \N__7127\
        );

    \I__1393\ : InMux
    port map (
            O => \N__7144\,
            I => \N__7127\
        );

    \I__1392\ : InMux
    port map (
            O => \N__7143\,
            I => \N__7122\
        );

    \I__1391\ : CascadeMux
    port map (
            O => \N__7142\,
            I => \N__7118\
        );

    \I__1390\ : InMux
    port map (
            O => \N__7139\,
            I => \N__7115\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__7138\,
            I => \N__7109\
        );

    \I__1388\ : Span4Mux_h
    port map (
            O => \N__7135\,
            I => \N__7102\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__7132\,
            I => \N__7102\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__7127\,
            I => \N__7102\
        );

    \I__1385\ : InMux
    port map (
            O => \N__7126\,
            I => \N__7099\
        );

    \I__1384\ : InMux
    port map (
            O => \N__7125\,
            I => \N__7094\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__7122\,
            I => \N__7091\
        );

    \I__1382\ : InMux
    port map (
            O => \N__7121\,
            I => \N__7086\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7118\,
            I => \N__7086\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7115\,
            I => \N__7083\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7114\,
            I => \N__7080\
        );

    \I__1378\ : CascadeMux
    port map (
            O => \N__7113\,
            I => \N__7076\
        );

    \I__1377\ : CascadeMux
    port map (
            O => \N__7112\,
            I => \N__7073\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7109\,
            I => \N__7066\
        );

    \I__1375\ : Span4Mux_v
    port map (
            O => \N__7102\,
            I => \N__7063\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__7099\,
            I => \N__7060\
        );

    \I__1373\ : InMux
    port map (
            O => \N__7098\,
            I => \N__7055\
        );

    \I__1372\ : InMux
    port map (
            O => \N__7097\,
            I => \N__7055\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__7094\,
            I => \N__7044\
        );

    \I__1370\ : Span4Mux_v
    port map (
            O => \N__7091\,
            I => \N__7044\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__7086\,
            I => \N__7044\
        );

    \I__1368\ : Span4Mux_v
    port map (
            O => \N__7083\,
            I => \N__7044\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__7080\,
            I => \N__7044\
        );

    \I__1366\ : InMux
    port map (
            O => \N__7079\,
            I => \N__7037\
        );

    \I__1365\ : InMux
    port map (
            O => \N__7076\,
            I => \N__7037\
        );

    \I__1364\ : InMux
    port map (
            O => \N__7073\,
            I => \N__7037\
        );

    \I__1363\ : InMux
    port map (
            O => \N__7072\,
            I => \N__7034\
        );

    \I__1362\ : InMux
    port map (
            O => \N__7071\,
            I => \N__7031\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7070\,
            I => \N__7026\
        );

    \I__1360\ : InMux
    port map (
            O => \N__7069\,
            I => \N__7026\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__7066\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1358\ : Odrv4
    port map (
            O => \N__7063\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1357\ : Odrv12
    port map (
            O => \N__7060\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__7055\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1355\ : Odrv4
    port map (
            O => \N__7044\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__7037\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__7034\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__7031\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__7026\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1350\ : InMux
    port map (
            O => \N__7007\,
            I => \N__7004\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__7004\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_i_0\
        );

    \I__1348\ : InMux
    port map (
            O => \N__7001\,
            I => \N__6997\
        );

    \I__1347\ : InMux
    port map (
            O => \N__7000\,
            I => \N__6994\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__6997\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__6994\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__1344\ : InMux
    port map (
            O => \N__6989\,
            I => \N__6985\
        );

    \I__1343\ : InMux
    port map (
            O => \N__6988\,
            I => \N__6982\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__6985\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__6982\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1340\ : CascadeMux
    port map (
            O => \N__6977\,
            I => \N__6973\
        );

    \I__1339\ : InMux
    port map (
            O => \N__6976\,
            I => \N__6970\
        );

    \I__1338\ : InMux
    port map (
            O => \N__6973\,
            I => \N__6967\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__6970\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__6967\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__1335\ : InMux
    port map (
            O => \N__6962\,
            I => \N__6958\
        );

    \I__1334\ : InMux
    port map (
            O => \N__6961\,
            I => \N__6955\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__6958\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__6955\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__1331\ : InMux
    port map (
            O => \N__6950\,
            I => \N__6946\
        );

    \I__1330\ : InMux
    port map (
            O => \N__6949\,
            I => \N__6943\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__6946\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__6943\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1327\ : InMux
    port map (
            O => \N__6938\,
            I => \N__6934\
        );

    \I__1326\ : InMux
    port map (
            O => \N__6937\,
            I => \N__6931\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__6934\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__6931\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1323\ : InMux
    port map (
            O => \N__6926\,
            I => \N__6922\
        );

    \I__1322\ : InMux
    port map (
            O => \N__6925\,
            I => \N__6919\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__6922\,
            I => \N__6916\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__6919\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1319\ : Odrv4
    port map (
            O => \N__6916\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1318\ : InMux
    port map (
            O => \N__6911\,
            I => \N__6908\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__6908\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__6905\,
            I => \N__6902\
        );

    \I__1315\ : InMux
    port map (
            O => \N__6902\,
            I => \N__6898\
        );

    \I__1314\ : InMux
    port map (
            O => \N__6901\,
            I => \N__6895\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__6898\,
            I => \N__6892\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__6895\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1311\ : Odrv12
    port map (
            O => \N__6892\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1310\ : InMux
    port map (
            O => \N__6887\,
            I => \N__6884\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__6884\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__1308\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6877\
        );

    \I__1307\ : InMux
    port map (
            O => \N__6880\,
            I => \N__6874\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__6877\,
            I => \N__6871\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__6874\,
            I => \N__6866\
        );

    \I__1304\ : Span4Mux_h
    port map (
            O => \N__6871\,
            I => \N__6863\
        );

    \I__1303\ : InMux
    port map (
            O => \N__6870\,
            I => \N__6860\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6869\,
            I => \N__6857\
        );

    \I__1301\ : Odrv4
    port map (
            O => \N__6866\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1300\ : Odrv4
    port map (
            O => \N__6863\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__6860\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__6857\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1297\ : InMux
    port map (
            O => \N__6848\,
            I => \N__6835\
        );

    \I__1296\ : InMux
    port map (
            O => \N__6847\,
            I => \N__6835\
        );

    \I__1295\ : InMux
    port map (
            O => \N__6846\,
            I => \N__6835\
        );

    \I__1294\ : InMux
    port map (
            O => \N__6845\,
            I => \N__6828\
        );

    \I__1293\ : InMux
    port map (
            O => \N__6844\,
            I => \N__6828\
        );

    \I__1292\ : InMux
    port map (
            O => \N__6843\,
            I => \N__6828\
        );

    \I__1291\ : InMux
    port map (
            O => \N__6842\,
            I => \N__6825\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__6835\,
            I => \N__6820\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__6828\,
            I => \N__6820\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__6825\,
            I => \U712_CHIP_RAM.N_62\
        );

    \I__1287\ : Odrv4
    port map (
            O => \N__6820\,
            I => \U712_CHIP_RAM.N_62\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6815\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__6812\,
            I => \N__6808\
        );

    \I__1284\ : InMux
    port map (
            O => \N__6811\,
            I => \N__6805\
        );

    \I__1283\ : InMux
    port map (
            O => \N__6808\,
            I => \N__6802\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__6805\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__6802\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1280\ : CEMux
    port map (
            O => \N__6797\,
            I => \N__6793\
        );

    \I__1279\ : CEMux
    port map (
            O => \N__6796\,
            I => \N__6790\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__6793\,
            I => \N__6787\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6790\,
            I => \N__6784\
        );

    \I__1276\ : Odrv4
    port map (
            O => \N__6787\,
            I => \U712_CHIP_RAM.N_434_i\
        );

    \I__1275\ : Odrv4
    port map (
            O => \N__6784\,
            I => \U712_CHIP_RAM.N_434_i\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6779\,
            I => \bfn_11_7_0_\
        );

    \I__1273\ : InMux
    port map (
            O => \N__6776\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__1272\ : InMux
    port map (
            O => \N__6773\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__1271\ : InMux
    port map (
            O => \N__6770\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__1270\ : InMux
    port map (
            O => \N__6767\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__1269\ : InMux
    port map (
            O => \N__6764\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__1268\ : InMux
    port map (
            O => \N__6761\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__1267\ : InMux
    port map (
            O => \N__6758\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__1266\ : CascadeMux
    port map (
            O => \N__6755\,
            I => \N__6751\
        );

    \I__1265\ : CascadeMux
    port map (
            O => \N__6754\,
            I => \N__6748\
        );

    \I__1264\ : InMux
    port map (
            O => \N__6751\,
            I => \N__6744\
        );

    \I__1263\ : InMux
    port map (
            O => \N__6748\,
            I => \N__6741\
        );

    \I__1262\ : InMux
    port map (
            O => \N__6747\,
            I => \N__6738\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__6744\,
            I => \N__6735\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__6741\,
            I => \N__6726\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__6738\,
            I => \N__6723\
        );

    \I__1258\ : Glb2LocalMux
    port map (
            O => \N__6735\,
            I => \N__6704\
        );

    \I__1257\ : ClkMux
    port map (
            O => \N__6734\,
            I => \N__6704\
        );

    \I__1256\ : ClkMux
    port map (
            O => \N__6733\,
            I => \N__6704\
        );

    \I__1255\ : ClkMux
    port map (
            O => \N__6732\,
            I => \N__6704\
        );

    \I__1254\ : ClkMux
    port map (
            O => \N__6731\,
            I => \N__6704\
        );

    \I__1253\ : ClkMux
    port map (
            O => \N__6730\,
            I => \N__6704\
        );

    \I__1252\ : ClkMux
    port map (
            O => \N__6729\,
            I => \N__6704\
        );

    \I__1251\ : Glb2LocalMux
    port map (
            O => \N__6726\,
            I => \N__6704\
        );

    \I__1250\ : Glb2LocalMux
    port map (
            O => \N__6723\,
            I => \N__6704\
        );

    \I__1249\ : GlobalMux
    port map (
            O => \N__6704\,
            I => \N__6701\
        );

    \I__1248\ : gio2CtrlBuf
    port map (
            O => \N__6701\,
            I => \C1_c_g\
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__6698\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\
        );

    \I__1246\ : CascadeMux
    port map (
            O => \N__6695\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_\
        );

    \I__1245\ : IoInMux
    port map (
            O => \N__6692\,
            I => \N__6689\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__6689\,
            I => \N__6686\
        );

    \I__1243\ : IoSpan4Mux
    port map (
            O => \N__6686\,
            I => \N__6683\
        );

    \I__1242\ : Span4Mux_s3_h
    port map (
            O => \N__6683\,
            I => \N__6680\
        );

    \I__1241\ : Sp12to4
    port map (
            O => \N__6680\,
            I => \N__6677\
        );

    \I__1240\ : Span12Mux_h
    port map (
            O => \N__6677\,
            I => \N__6674\
        );

    \I__1239\ : Odrv12
    port map (
            O => \N__6674\,
            I => \CMA_c_6\
        );

    \I__1238\ : InMux
    port map (
            O => \N__6671\,
            I => \N__6668\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__6668\,
            I => \N__6665\
        );

    \I__1236\ : Span4Mux_h
    port map (
            O => \N__6665\,
            I => \N__6662\
        );

    \I__1235\ : Odrv4
    port map (
            O => \N__6662\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_1\
        );

    \I__1234\ : InMux
    port map (
            O => \N__6659\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__1233\ : InMux
    port map (
            O => \N__6656\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__1232\ : InMux
    port map (
            O => \N__6653\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__1231\ : InMux
    port map (
            O => \N__6650\,
            I => \N__6646\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6649\,
            I => \N__6643\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__6646\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__6643\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1227\ : InMux
    port map (
            O => \N__6638\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__1226\ : InMux
    port map (
            O => \N__6635\,
            I => \N__6631\
        );

    \I__1225\ : InMux
    port map (
            O => \N__6634\,
            I => \N__6628\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__6631\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__6628\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1222\ : InMux
    port map (
            O => \N__6623\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6620\,
            I => \N__6616\
        );

    \I__1220\ : InMux
    port map (
            O => \N__6619\,
            I => \N__6613\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__6616\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__6613\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1217\ : InMux
    port map (
            O => \N__6608\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__1216\ : InMux
    port map (
            O => \N__6605\,
            I => \N__6602\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__6602\,
            I => \N__6599\
        );

    \I__1214\ : Odrv12
    port map (
            O => \N__6599\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2Z0Z_0\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6596\,
            I => \N__6593\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__6593\,
            I => \U712_BYTE_ENABLE.N_431\
        );

    \I__1211\ : CascadeMux
    port map (
            O => \N__6590\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2Z0Z_0_cascade_\
        );

    \I__1210\ : IoInMux
    port map (
            O => \N__6587\,
            I => \N__6584\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__6584\,
            I => \N__6581\
        );

    \I__1208\ : Span12Mux_s3_v
    port map (
            O => \N__6581\,
            I => \N__6578\
        );

    \I__1207\ : Span12Mux_v
    port map (
            O => \N__6578\,
            I => \N__6575\
        );

    \I__1206\ : Odrv12
    port map (
            O => \N__6575\,
            I => \N_45_i\
        );

    \I__1205\ : InMux
    port map (
            O => \N__6572\,
            I => \N__6566\
        );

    \I__1204\ : InMux
    port map (
            O => \N__6571\,
            I => \N__6566\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__6566\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2Z0Z_0\
        );

    \I__1202\ : InMux
    port map (
            O => \N__6563\,
            I => \N__6559\
        );

    \I__1201\ : InMux
    port map (
            O => \N__6562\,
            I => \N__6556\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__6559\,
            I => \N__6551\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__6556\,
            I => \N__6548\
        );

    \I__1198\ : InMux
    port map (
            O => \N__6555\,
            I => \N__6545\
        );

    \I__1197\ : InMux
    port map (
            O => \N__6554\,
            I => \N__6542\
        );

    \I__1196\ : Span4Mux_v
    port map (
            O => \N__6551\,
            I => \N__6539\
        );

    \I__1195\ : Span4Mux_v
    port map (
            O => \N__6548\,
            I => \N__6536\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__6545\,
            I => \N__6533\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__6542\,
            I => \N__6530\
        );

    \I__1192\ : Sp12to4
    port map (
            O => \N__6539\,
            I => \N__6525\
        );

    \I__1191\ : Sp12to4
    port map (
            O => \N__6536\,
            I => \N__6525\
        );

    \I__1190\ : Span4Mux_v
    port map (
            O => \N__6533\,
            I => \N__6522\
        );

    \I__1189\ : Span12Mux_h
    port map (
            O => \N__6530\,
            I => \N__6519\
        );

    \I__1188\ : Span12Mux_h
    port map (
            O => \N__6525\,
            I => \N__6516\
        );

    \I__1187\ : Sp12to4
    port map (
            O => \N__6522\,
            I => \N__6513\
        );

    \I__1186\ : Span12Mux_v
    port map (
            O => \N__6519\,
            I => \N__6510\
        );

    \I__1185\ : Span12Mux_v
    port map (
            O => \N__6516\,
            I => \N__6505\
        );

    \I__1184\ : Span12Mux_h
    port map (
            O => \N__6513\,
            I => \N__6505\
        );

    \I__1183\ : Odrv12
    port map (
            O => \N__6510\,
            I => \RnW_c\
        );

    \I__1182\ : Odrv12
    port map (
            O => \N__6505\,
            I => \RnW_c\
        );

    \I__1181\ : IoInMux
    port map (
            O => \N__6500\,
            I => \N__6497\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6497\,
            I => \N__6494\
        );

    \I__1179\ : IoSpan4Mux
    port map (
            O => \N__6494\,
            I => \N__6491\
        );

    \I__1178\ : Span4Mux_s1_h
    port map (
            O => \N__6491\,
            I => \N__6488\
        );

    \I__1177\ : Span4Mux_v
    port map (
            O => \N__6488\,
            I => \N__6485\
        );

    \I__1176\ : Sp12to4
    port map (
            O => \N__6485\,
            I => \N__6482\
        );

    \I__1175\ : Span12Mux_s10_h
    port map (
            O => \N__6482\,
            I => \N__6479\
        );

    \I__1174\ : Odrv12
    port map (
            O => \N__6479\,
            I => \N_344\
        );

    \I__1173\ : IoInMux
    port map (
            O => \N__6476\,
            I => \N__6473\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__6473\,
            I => \N__6470\
        );

    \I__1171\ : Span12Mux_s8_v
    port map (
            O => \N__6470\,
            I => \N__6467\
        );

    \I__1170\ : Odrv12
    port map (
            O => \N__6467\,
            I => \DMA_LATCH_EN_c\
        );

    \I__1169\ : InMux
    port map (
            O => \N__6464\,
            I => \N__6461\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__6461\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\
        );

    \I__1167\ : InMux
    port map (
            O => \N__6458\,
            I => \N__6455\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6455\,
            I => \N__6452\
        );

    \I__1165\ : Odrv4
    port map (
            O => \N__6452\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__1164\ : CascadeMux
    port map (
            O => \N__6449\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_\
        );

    \I__1163\ : IoInMux
    port map (
            O => \N__6446\,
            I => \N__6443\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__6443\,
            I => \N__6440\
        );

    \I__1161\ : Span4Mux_s1_h
    port map (
            O => \N__6440\,
            I => \N__6437\
        );

    \I__1160\ : Sp12to4
    port map (
            O => \N__6437\,
            I => \N__6434\
        );

    \I__1159\ : Span12Mux_s10_v
    port map (
            O => \N__6434\,
            I => \N__6431\
        );

    \I__1158\ : Span12Mux_h
    port map (
            O => \N__6431\,
            I => \N__6428\
        );

    \I__1157\ : Odrv12
    port map (
            O => \N__6428\,
            I => \CMA_c_7\
        );

    \I__1156\ : InMux
    port map (
            O => \N__6425\,
            I => \N__6422\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__6422\,
            I => \N__6419\
        );

    \I__1154\ : Span4Mux_v
    port map (
            O => \N__6419\,
            I => \N__6416\
        );

    \I__1153\ : Span4Mux_v
    port map (
            O => \N__6416\,
            I => \N__6413\
        );

    \I__1152\ : Sp12to4
    port map (
            O => \N__6413\,
            I => \N__6410\
        );

    \I__1151\ : Span12Mux_h
    port map (
            O => \N__6410\,
            I => \N__6407\
        );

    \I__1150\ : Odrv12
    port map (
            O => \N__6407\,
            I => \A_c_8\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6404\,
            I => \N__6401\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__6401\,
            I => \N__6398\
        );

    \I__1147\ : Sp12to4
    port map (
            O => \N__6398\,
            I => \N__6395\
        );

    \I__1146\ : Span12Mux_v
    port map (
            O => \N__6395\,
            I => \N__6392\
        );

    \I__1145\ : Span12Mux_h
    port map (
            O => \N__6392\,
            I => \N__6389\
        );

    \I__1144\ : Odrv12
    port map (
            O => \N__6389\,
            I => \A_c_15\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__6386\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNO_6Z0Z_1_cascade_\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6383\,
            I => \N__6380\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__6380\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6377\,
            I => \N__6371\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__6376\,
            I => \N__6368\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6375\,
            I => \N__6365\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6374\,
            I => \N__6361\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6371\,
            I => \N__6358\
        );

    \I__1135\ : InMux
    port map (
            O => \N__6368\,
            I => \N__6351\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__6365\,
            I => \N__6348\
        );

    \I__1133\ : InMux
    port map (
            O => \N__6364\,
            I => \N__6345\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__6361\,
            I => \N__6340\
        );

    \I__1131\ : Span4Mux_h
    port map (
            O => \N__6358\,
            I => \N__6340\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6357\,
            I => \N__6337\
        );

    \I__1129\ : InMux
    port map (
            O => \N__6356\,
            I => \N__6330\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6355\,
            I => \N__6330\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6354\,
            I => \N__6330\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__6351\,
            I => \U712_CHIP_RAM.N_287\
        );

    \I__1125\ : Odrv4
    port map (
            O => \N__6348\,
            I => \U712_CHIP_RAM.N_287\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__6345\,
            I => \U712_CHIP_RAM.N_287\
        );

    \I__1123\ : Odrv4
    port map (
            O => \N__6340\,
            I => \U712_CHIP_RAM.N_287\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__6337\,
            I => \U712_CHIP_RAM.N_287\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__6330\,
            I => \U712_CHIP_RAM.N_287\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6317\,
            I => \N__6314\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__6314\,
            I => \N__6311\
        );

    \I__1118\ : Span4Mux_v
    port map (
            O => \N__6311\,
            I => \N__6308\
        );

    \I__1117\ : Odrv4
    port map (
            O => \N__6308\,
            I => \U712_CHIP_RAM.N_388\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6305\,
            I => \N__6302\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__6302\,
            I => \U712_CHIP_RAM.N_370\
        );

    \I__1114\ : InMux
    port map (
            O => \N__6299\,
            I => \N__6296\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__6296\,
            I => \U712_BYTE_ENABLE.un1_CUUBEn_i_0_aZ0Z2\
        );

    \I__1112\ : IoInMux
    port map (
            O => \N__6293\,
            I => \N__6290\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__6290\,
            I => \N__6287\
        );

    \I__1110\ : IoSpan4Mux
    port map (
            O => \N__6287\,
            I => \N__6284\
        );

    \I__1109\ : Span4Mux_s1_h
    port map (
            O => \N__6284\,
            I => \N__6281\
        );

    \I__1108\ : Span4Mux_v
    port map (
            O => \N__6281\,
            I => \N__6278\
        );

    \I__1107\ : Sp12to4
    port map (
            O => \N__6278\,
            I => \N__6275\
        );

    \I__1106\ : Span12Mux_s10_h
    port map (
            O => \N__6275\,
            I => \N__6272\
        );

    \I__1105\ : Odrv12
    port map (
            O => \N__6272\,
            I => \N_38_i\
        );

    \I__1104\ : CascadeMux
    port map (
            O => \N__6269\,
            I => \U712_BYTE_ENABLE.N_426_cascade_\
        );

    \I__1103\ : IoInMux
    port map (
            O => \N__6266\,
            I => \N__6263\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__6263\,
            I => \N__6260\
        );

    \I__1101\ : IoSpan4Mux
    port map (
            O => \N__6260\,
            I => \N__6257\
        );

    \I__1100\ : Span4Mux_s1_h
    port map (
            O => \N__6257\,
            I => \N__6254\
        );

    \I__1099\ : Sp12to4
    port map (
            O => \N__6254\,
            I => \N__6251\
        );

    \I__1098\ : Span12Mux_h
    port map (
            O => \N__6251\,
            I => \N__6248\
        );

    \I__1097\ : Span12Mux_v
    port map (
            O => \N__6248\,
            I => \N__6245\
        );

    \I__1096\ : Odrv12
    port map (
            O => \N__6245\,
            I => \N_47_i\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6242\,
            I => \N__6239\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6239\,
            I => \N__6236\
        );

    \I__1093\ : Odrv4
    port map (
            O => \N__6236\,
            I => \U712_BYTE_ENABLE.un1_CLMBEn_i_0_aZ0Z2\
        );

    \I__1092\ : IoInMux
    port map (
            O => \N__6233\,
            I => \N__6230\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__6230\,
            I => \N__6225\
        );

    \I__1090\ : CascadeMux
    port map (
            O => \N__6229\,
            I => \N__6220\
        );

    \I__1089\ : CascadeMux
    port map (
            O => \N__6228\,
            I => \N__6217\
        );

    \I__1088\ : IoSpan4Mux
    port map (
            O => \N__6225\,
            I => \N__6214\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6224\,
            I => \N__6205\
        );

    \I__1086\ : InMux
    port map (
            O => \N__6223\,
            I => \N__6205\
        );

    \I__1085\ : InMux
    port map (
            O => \N__6220\,
            I => \N__6205\
        );

    \I__1084\ : InMux
    port map (
            O => \N__6217\,
            I => \N__6205\
        );

    \I__1083\ : Span4Mux_s3_v
    port map (
            O => \N__6214\,
            I => \N__6202\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__6205\,
            I => \N__6199\
        );

    \I__1081\ : Span4Mux_v
    port map (
            O => \N__6202\,
            I => \N__6195\
        );

    \I__1080\ : Span4Mux_v
    port map (
            O => \N__6199\,
            I => \N__6192\
        );

    \I__1079\ : InMux
    port map (
            O => \N__6198\,
            I => \N__6189\
        );

    \I__1078\ : Odrv4
    port map (
            O => \N__6195\,
            I => \DBENn_c\
        );

    \I__1077\ : Odrv4
    port map (
            O => \N__6192\,
            I => \DBENn_c\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__6189\,
            I => \DBENn_c\
        );

    \I__1075\ : IoInMux
    port map (
            O => \N__6182\,
            I => \N__6179\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__6179\,
            I => \N__6176\
        );

    \I__1073\ : Span4Mux_s2_h
    port map (
            O => \N__6176\,
            I => \N__6173\
        );

    \I__1072\ : Span4Mux_h
    port map (
            O => \N__6173\,
            I => \N__6170\
        );

    \I__1071\ : Sp12to4
    port map (
            O => \N__6170\,
            I => \N__6167\
        );

    \I__1070\ : Span12Mux_v
    port map (
            O => \N__6167\,
            I => \N__6164\
        );

    \I__1069\ : Odrv12
    port map (
            O => \N__6164\,
            I => \N_46_i\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__6161\,
            I => \U712_CHIP_RAM.N_287_cascade_\
        );

    \I__1067\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6155\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__6155\,
            I => \U712_CHIP_RAM.N_436\
        );

    \I__1065\ : CascadeMux
    port map (
            O => \N__6152\,
            I => \N__6148\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6151\,
            I => \N__6141\
        );

    \I__1063\ : InMux
    port map (
            O => \N__6148\,
            I => \N__6141\
        );

    \I__1062\ : InMux
    port map (
            O => \N__6147\,
            I => \N__6136\
        );

    \I__1061\ : InMux
    port map (
            O => \N__6146\,
            I => \N__6136\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__6141\,
            I => \N__6133\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__6136\,
            I => \N__6130\
        );

    \I__1058\ : Span4Mux_h
    port map (
            O => \N__6133\,
            I => \N__6127\
        );

    \I__1057\ : Odrv4
    port map (
            O => \N__6130\,
            I => \U712_CHIP_RAM.N_283\
        );

    \I__1056\ : Odrv4
    port map (
            O => \N__6127\,
            I => \U712_CHIP_RAM.N_283\
        );

    \I__1055\ : CascadeMux
    port map (
            O => \N__6122\,
            I => \N__6119\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6119\,
            I => \N__6116\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__6116\,
            I => \N__6113\
        );

    \I__1052\ : Odrv12
    port map (
            O => \N__6113\,
            I => \U712_CHIP_RAM.N_347\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6110\,
            I => \N__6107\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__6107\,
            I => \N__6104\
        );

    \I__1049\ : Odrv4
    port map (
            O => \N__6104\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_i_0_2\
        );

    \I__1048\ : CascadeMux
    port map (
            O => \N__6101\,
            I => \N__6098\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6098\,
            I => \N__6095\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__6095\,
            I => \N__6092\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__6092\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_129_i_0_0\
        );

    \I__1044\ : CascadeMux
    port map (
            O => \N__6089\,
            I => \N__6084\
        );

    \I__1043\ : InMux
    port map (
            O => \N__6088\,
            I => \N__6078\
        );

    \I__1042\ : InMux
    port map (
            O => \N__6087\,
            I => \N__6075\
        );

    \I__1041\ : InMux
    port map (
            O => \N__6084\,
            I => \N__6070\
        );

    \I__1040\ : InMux
    port map (
            O => \N__6083\,
            I => \N__6059\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6082\,
            I => \N__6059\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6059\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__6078\,
            I => \N__6056\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__6075\,
            I => \N__6053\
        );

    \I__1035\ : InMux
    port map (
            O => \N__6074\,
            I => \N__6050\
        );

    \I__1034\ : InMux
    port map (
            O => \N__6073\,
            I => \N__6047\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__6070\,
            I => \N__6044\
        );

    \I__1032\ : InMux
    port map (
            O => \N__6069\,
            I => \N__6039\
        );

    \I__1031\ : InMux
    port map (
            O => \N__6068\,
            I => \N__6039\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6067\,
            I => \N__6034\
        );

    \I__1029\ : InMux
    port map (
            O => \N__6066\,
            I => \N__6034\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__6059\,
            I => \U712_CHIP_RAM.N_286\
        );

    \I__1027\ : Odrv4
    port map (
            O => \N__6056\,
            I => \U712_CHIP_RAM.N_286\
        );

    \I__1026\ : Odrv4
    port map (
            O => \N__6053\,
            I => \U712_CHIP_RAM.N_286\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__6050\,
            I => \U712_CHIP_RAM.N_286\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__6047\,
            I => \U712_CHIP_RAM.N_286\
        );

    \I__1023\ : Odrv12
    port map (
            O => \N__6044\,
            I => \U712_CHIP_RAM.N_286\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__6039\,
            I => \U712_CHIP_RAM.N_286\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__6034\,
            I => \U712_CHIP_RAM.N_286\
        );

    \I__1020\ : CEMux
    port map (
            O => \N__6017\,
            I => \N__6014\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__6014\,
            I => \N__6011\
        );

    \I__1018\ : Odrv4
    port map (
            O => \N__6011\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__6008\,
            I => \N__6005\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6005\,
            I => \N__6000\
        );

    \I__1015\ : InMux
    port map (
            O => \N__6004\,
            I => \N__5997\
        );

    \I__1014\ : InMux
    port map (
            O => \N__6003\,
            I => \N__5994\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__6000\,
            I => \N__5988\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__5997\,
            I => \N__5983\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__5994\,
            I => \N__5983\
        );

    \I__1010\ : InMux
    port map (
            O => \N__5993\,
            I => \N__5980\
        );

    \I__1009\ : InMux
    port map (
            O => \N__5992\,
            I => \N__5977\
        );

    \I__1008\ : InMux
    port map (
            O => \N__5991\,
            I => \N__5974\
        );

    \I__1007\ : Span4Mux_h
    port map (
            O => \N__5988\,
            I => \N__5971\
        );

    \I__1006\ : Span4Mux_h
    port map (
            O => \N__5983\,
            I => \N__5966\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__5980\,
            I => \N__5966\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__5977\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5974\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1002\ : Odrv4
    port map (
            O => \N__5971\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1001\ : Odrv4
    port map (
            O => \N__5966\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1000\ : CascadeMux
    port map (
            O => \N__5957\,
            I => \N__5954\
        );

    \I__999\ : InMux
    port map (
            O => \N__5954\,
            I => \N__5950\
        );

    \I__998\ : InMux
    port map (
            O => \N__5953\,
            I => \N__5945\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__5950\,
            I => \N__5942\
        );

    \I__996\ : InMux
    port map (
            O => \N__5949\,
            I => \N__5939\
        );

    \I__995\ : InMux
    port map (
            O => \N__5948\,
            I => \N__5936\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5945\,
            I => \N__5929\
        );

    \I__993\ : Span4Mux_h
    port map (
            O => \N__5942\,
            I => \N__5929\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__5939\,
            I => \N__5929\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__5936\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__990\ : Odrv4
    port map (
            O => \N__5929\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__989\ : CascadeMux
    port map (
            O => \N__5924\,
            I => \N__5921\
        );

    \I__988\ : InMux
    port map (
            O => \N__5921\,
            I => \N__5916\
        );

    \I__987\ : InMux
    port map (
            O => \N__5920\,
            I => \N__5911\
        );

    \I__986\ : InMux
    port map (
            O => \N__5919\,
            I => \N__5908\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__5916\,
            I => \N__5905\
        );

    \I__984\ : InMux
    port map (
            O => \N__5915\,
            I => \N__5902\
        );

    \I__983\ : InMux
    port map (
            O => \N__5914\,
            I => \N__5899\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__5911\,
            I => \N__5892\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__5908\,
            I => \N__5892\
        );

    \I__980\ : Span4Mux_h
    port map (
            O => \N__5905\,
            I => \N__5892\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__5902\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__5899\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__977\ : Odrv4
    port map (
            O => \N__5892\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__976\ : InMux
    port map (
            O => \N__5885\,
            I => \N__5880\
        );

    \I__975\ : InMux
    port map (
            O => \N__5884\,
            I => \N__5877\
        );

    \I__974\ : InMux
    port map (
            O => \N__5883\,
            I => \N__5874\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__5880\,
            I => \N__5866\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__5877\,
            I => \N__5863\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__5874\,
            I => \N__5860\
        );

    \I__970\ : InMux
    port map (
            O => \N__5873\,
            I => \N__5857\
        );

    \I__969\ : InMux
    port map (
            O => \N__5872\,
            I => \N__5854\
        );

    \I__968\ : InMux
    port map (
            O => \N__5871\,
            I => \N__5851\
        );

    \I__967\ : InMux
    port map (
            O => \N__5870\,
            I => \N__5846\
        );

    \I__966\ : InMux
    port map (
            O => \N__5869\,
            I => \N__5846\
        );

    \I__965\ : Span4Mux_h
    port map (
            O => \N__5866\,
            I => \N__5843\
        );

    \I__964\ : Span4Mux_h
    port map (
            O => \N__5863\,
            I => \N__5836\
        );

    \I__963\ : Span4Mux_h
    port map (
            O => \N__5860\,
            I => \N__5836\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__5857\,
            I => \N__5836\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__5854\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__5851\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__5846\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__958\ : Odrv4
    port map (
            O => \N__5843\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__957\ : Odrv4
    port map (
            O => \N__5836\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__956\ : CascadeMux
    port map (
            O => \N__5825\,
            I => \U712_REG_SM.C1_SYNC_RNIAS4F1_0Z0Z_1_cascade_\
        );

    \I__955\ : InMux
    port map (
            O => \N__5822\,
            I => \N__5819\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__5819\,
            I => \N__5816\
        );

    \I__953\ : Span4Mux_v
    port map (
            O => \N__5816\,
            I => \N__5812\
        );

    \I__952\ : InMux
    port map (
            O => \N__5815\,
            I => \N__5809\
        );

    \I__951\ : Sp12to4
    port map (
            O => \N__5812\,
            I => \N__5804\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__5809\,
            I => \N__5804\
        );

    \I__949\ : Odrv12
    port map (
            O => \N__5804\,
            I => \U712_REG_SM.ASn_0_sqmuxa_1\
        );

    \I__948\ : InMux
    port map (
            O => \N__5801\,
            I => \N__5798\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__5798\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a2_0_1\
        );

    \I__946\ : CascadeMux
    port map (
            O => \N__5795\,
            I => \N__5787\
        );

    \I__945\ : InMux
    port map (
            O => \N__5794\,
            I => \N__5782\
        );

    \I__944\ : InMux
    port map (
            O => \N__5793\,
            I => \N__5782\
        );

    \I__943\ : InMux
    port map (
            O => \N__5792\,
            I => \N__5777\
        );

    \I__942\ : InMux
    port map (
            O => \N__5791\,
            I => \N__5777\
        );

    \I__941\ : InMux
    port map (
            O => \N__5790\,
            I => \N__5774\
        );

    \I__940\ : InMux
    port map (
            O => \N__5787\,
            I => \N__5771\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__5782\,
            I => \N__5766\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__5777\,
            I => \N__5766\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__5774\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__5771\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__935\ : Odrv12
    port map (
            O => \N__5766\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__934\ : CascadeMux
    port map (
            O => \N__5759\,
            I => \N__5756\
        );

    \I__933\ : InMux
    port map (
            O => \N__5756\,
            I => \N__5752\
        );

    \I__932\ : CascadeMux
    port map (
            O => \N__5755\,
            I => \N__5749\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__5752\,
            I => \N__5744\
        );

    \I__930\ : InMux
    port map (
            O => \N__5749\,
            I => \N__5741\
        );

    \I__929\ : InMux
    port map (
            O => \N__5748\,
            I => \N__5738\
        );

    \I__928\ : InMux
    port map (
            O => \N__5747\,
            I => \N__5735\
        );

    \I__927\ : Span4Mux_h
    port map (
            O => \N__5744\,
            I => \N__5732\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__5741\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__5738\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__5735\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__923\ : Odrv4
    port map (
            O => \N__5732\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__5723\,
            I => \N__5719\
        );

    \I__921\ : InMux
    port map (
            O => \N__5722\,
            I => \N__5716\
        );

    \I__920\ : InMux
    port map (
            O => \N__5719\,
            I => \N__5713\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__5716\,
            I => \N__5707\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5713\,
            I => \N__5707\
        );

    \I__917\ : InMux
    port map (
            O => \N__5712\,
            I => \N__5704\
        );

    \I__916\ : Odrv12
    port map (
            O => \N__5707\,
            I => \U712_REG_SM.C1_SYNC_RNIAS4F1_0Z0Z_1\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__5704\,
            I => \U712_REG_SM.C1_SYNC_RNIAS4F1_0Z0Z_1\
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__5699\,
            I => \N__5696\
        );

    \I__913\ : InMux
    port map (
            O => \N__5696\,
            I => \N__5693\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__5693\,
            I => \N__5690\
        );

    \I__911\ : Odrv4
    port map (
            O => \N__5690\,
            I => \U712_REG_SM.N_104\
        );

    \I__910\ : CascadeMux
    port map (
            O => \N__5687\,
            I => \U712_CHIP_RAM.N_414_cascade_\
        );

    \I__909\ : InMux
    port map (
            O => \N__5684\,
            I => \N__5681\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__5681\,
            I => \N__5678\
        );

    \I__907\ : Span4Mux_h
    port map (
            O => \N__5678\,
            I => \N__5675\
        );

    \I__906\ : Odrv4
    port map (
            O => \N__5675\,
            I => \U712_CHIP_RAM.N_86\
        );

    \I__905\ : InMux
    port map (
            O => \N__5672\,
            I => \N__5666\
        );

    \I__904\ : InMux
    port map (
            O => \N__5671\,
            I => \N__5663\
        );

    \I__903\ : InMux
    port map (
            O => \N__5670\,
            I => \N__5660\
        );

    \I__902\ : CascadeMux
    port map (
            O => \N__5669\,
            I => \N__5657\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__5666\,
            I => \N__5654\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__5663\,
            I => \N__5651\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__5660\,
            I => \N__5648\
        );

    \I__898\ : InMux
    port map (
            O => \N__5657\,
            I => \N__5644\
        );

    \I__897\ : Span4Mux_v
    port map (
            O => \N__5654\,
            I => \N__5641\
        );

    \I__896\ : Span4Mux_v
    port map (
            O => \N__5651\,
            I => \N__5636\
        );

    \I__895\ : Span4Mux_h
    port map (
            O => \N__5648\,
            I => \N__5636\
        );

    \I__894\ : InMux
    port map (
            O => \N__5647\,
            I => \N__5633\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__5644\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__892\ : Odrv4
    port map (
            O => \N__5641\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__891\ : Odrv4
    port map (
            O => \N__5636\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__5633\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__5624\,
            I => \N__5621\
        );

    \I__888\ : InMux
    port map (
            O => \N__5621\,
            I => \N__5614\
        );

    \I__887\ : InMux
    port map (
            O => \N__5620\,
            I => \N__5611\
        );

    \I__886\ : InMux
    port map (
            O => \N__5619\,
            I => \N__5608\
        );

    \I__885\ : InMux
    port map (
            O => \N__5618\,
            I => \N__5605\
        );

    \I__884\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5602\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__5614\,
            I => \N__5599\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__5611\,
            I => \N__5596\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__5608\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__5605\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__5602\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__878\ : Odrv4
    port map (
            O => \N__5599\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__877\ : Odrv12
    port map (
            O => \N__5596\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__876\ : InMux
    port map (
            O => \N__5585\,
            I => \N__5579\
        );

    \I__875\ : InMux
    port map (
            O => \N__5584\,
            I => \N__5579\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__5579\,
            I => \N__5576\
        );

    \I__873\ : Odrv4
    port map (
            O => \N__5576\,
            I => \U712_CHIP_RAM.N_373\
        );

    \I__872\ : InMux
    port map (
            O => \N__5573\,
            I => \N__5569\
        );

    \I__871\ : InMux
    port map (
            O => \N__5572\,
            I => \N__5564\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__5569\,
            I => \N__5560\
        );

    \I__869\ : InMux
    port map (
            O => \N__5568\,
            I => \N__5555\
        );

    \I__868\ : InMux
    port map (
            O => \N__5567\,
            I => \N__5555\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__5564\,
            I => \N__5552\
        );

    \I__866\ : InMux
    port map (
            O => \N__5563\,
            I => \N__5549\
        );

    \I__865\ : Span4Mux_v
    port map (
            O => \N__5560\,
            I => \N__5544\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__5555\,
            I => \N__5544\
        );

    \I__863\ : Odrv4
    port map (
            O => \N__5552\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__5549\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__861\ : Odrv4
    port map (
            O => \N__5544\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__5537\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_\
        );

    \I__859\ : InMux
    port map (
            O => \N__5534\,
            I => \N__5531\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5531\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_1\
        );

    \I__857\ : CascadeMux
    port map (
            O => \N__5528\,
            I => \U712_CHIP_RAM.N_286_cascade_\
        );

    \I__856\ : InMux
    port map (
            O => \N__5525\,
            I => \N__5522\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__5522\,
            I => \N__5517\
        );

    \I__854\ : InMux
    port map (
            O => \N__5521\,
            I => \N__5512\
        );

    \I__853\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5512\
        );

    \I__852\ : Odrv4
    port map (
            O => \N__5517\,
            I => \U712_CHIP_RAM.N_486\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__5512\,
            I => \U712_CHIP_RAM.N_486\
        );

    \I__850\ : InMux
    port map (
            O => \N__5507\,
            I => \N__5504\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__5504\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a2_1\
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__5501\,
            I => \U712_CHIP_RAM.N_371_1_cascade_\
        );

    \I__847\ : InMux
    port map (
            O => \N__5498\,
            I => \N__5495\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__5495\,
            I => \N__5492\
        );

    \I__845\ : Span4Mux_v
    port map (
            O => \N__5492\,
            I => \N__5489\
        );

    \I__844\ : Span4Mux_h
    port map (
            O => \N__5489\,
            I => \N__5486\
        );

    \I__843\ : Odrv4
    port map (
            O => \N__5486\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_a2_0\
        );

    \I__842\ : CascadeMux
    port map (
            O => \N__5483\,
            I => \N__5480\
        );

    \I__841\ : InMux
    port map (
            O => \N__5480\,
            I => \N__5477\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__5477\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_0_0_0\
        );

    \I__839\ : InMux
    port map (
            O => \N__5474\,
            I => \N__5471\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__5471\,
            I => \U712_CHIP_RAM.N_371_1\
        );

    \I__837\ : InMux
    port map (
            O => \N__5468\,
            I => \N__5465\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__5465\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__835\ : CascadeMux
    port map (
            O => \N__5462\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\
        );

    \I__834\ : CascadeMux
    port map (
            O => \N__5459\,
            I => \N__5456\
        );

    \I__833\ : InMux
    port map (
            O => \N__5456\,
            I => \N__5449\
        );

    \I__832\ : InMux
    port map (
            O => \N__5455\,
            I => \N__5449\
        );

    \I__831\ : InMux
    port map (
            O => \N__5454\,
            I => \N__5439\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__5449\,
            I => \N__5436\
        );

    \I__829\ : InMux
    port map (
            O => \N__5448\,
            I => \N__5433\
        );

    \I__828\ : InMux
    port map (
            O => \N__5447\,
            I => \N__5430\
        );

    \I__827\ : InMux
    port map (
            O => \N__5446\,
            I => \N__5427\
        );

    \I__826\ : InMux
    port map (
            O => \N__5445\,
            I => \N__5424\
        );

    \I__825\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5417\
        );

    \I__824\ : InMux
    port map (
            O => \N__5443\,
            I => \N__5417\
        );

    \I__823\ : InMux
    port map (
            O => \N__5442\,
            I => \N__5417\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5439\,
            I => \N__5414\
        );

    \I__821\ : Span4Mux_h
    port map (
            O => \N__5436\,
            I => \N__5411\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__5433\,
            I => \U712_CHIP_RAM.N_288\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__5430\,
            I => \U712_CHIP_RAM.N_288\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__5427\,
            I => \U712_CHIP_RAM.N_288\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__5424\,
            I => \U712_CHIP_RAM.N_288\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__5417\,
            I => \U712_CHIP_RAM.N_288\
        );

    \I__815\ : Odrv4
    port map (
            O => \N__5414\,
            I => \U712_CHIP_RAM.N_288\
        );

    \I__814\ : Odrv4
    port map (
            O => \N__5411\,
            I => \U712_CHIP_RAM.N_288\
        );

    \I__813\ : CEMux
    port map (
            O => \N__5396\,
            I => \N__5393\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5393\,
            I => \N__5390\
        );

    \I__811\ : Span4Mux_v
    port map (
            O => \N__5390\,
            I => \N__5387\
        );

    \I__810\ : Odrv4
    port map (
            O => \N__5387\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0\
        );

    \I__809\ : InMux
    port map (
            O => \N__5384\,
            I => \N__5381\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__5381\,
            I => \U712_CHIP_RAM.N_329\
        );

    \I__807\ : InMux
    port map (
            O => \N__5378\,
            I => \N__5375\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__5375\,
            I => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\
        );

    \I__805\ : CascadeMux
    port map (
            O => \N__5372\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_i_0_cascade_\
        );

    \I__804\ : InMux
    port map (
            O => \N__5369\,
            I => \N__5366\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5366\,
            I => \N__5362\
        );

    \I__802\ : InMux
    port map (
            O => \N__5365\,
            I => \N__5359\
        );

    \I__801\ : Odrv4
    port map (
            O => \N__5362\,
            I => \U712_CHIP_RAM.N_11_2\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__5359\,
            I => \U712_CHIP_RAM.N_11_2\
        );

    \I__799\ : InMux
    port map (
            O => \N__5354\,
            I => \N__5350\
        );

    \I__798\ : InMux
    port map (
            O => \N__5353\,
            I => \N__5347\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5350\,
            I => \N__5344\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__5347\,
            I => \REG_TACK\
        );

    \I__795\ : Odrv4
    port map (
            O => \N__5344\,
            I => \REG_TACK\
        );

    \I__794\ : InMux
    port map (
            O => \N__5339\,
            I => \N__5333\
        );

    \I__793\ : InMux
    port map (
            O => \N__5338\,
            I => \N__5333\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__5333\,
            I => \CPU_TACKm\
        );

    \I__791\ : CascadeMux
    port map (
            O => \N__5330\,
            I => \N__5327\
        );

    \I__790\ : InMux
    port map (
            O => \N__5327\,
            I => \N__5322\
        );

    \I__789\ : InMux
    port map (
            O => \N__5326\,
            I => \N__5319\
        );

    \I__788\ : InMux
    port map (
            O => \N__5325\,
            I => \N__5316\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5322\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__5319\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__5316\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__784\ : CascadeMux
    port map (
            O => \N__5309\,
            I => \N__5306\
        );

    \I__783\ : InMux
    port map (
            O => \N__5306\,
            I => \N__5302\
        );

    \I__782\ : InMux
    port map (
            O => \N__5305\,
            I => \N__5299\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__5302\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__5299\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__779\ : CascadeMux
    port map (
            O => \N__5294\,
            I => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\
        );

    \I__778\ : InMux
    port map (
            O => \N__5291\,
            I => \N__5286\
        );

    \I__777\ : InMux
    port map (
            O => \N__5290\,
            I => \N__5283\
        );

    \I__776\ : InMux
    port map (
            O => \N__5289\,
            I => \N__5280\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5286\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__5283\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__5280\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__772\ : InMux
    port map (
            O => \N__5273\,
            I => \N__5270\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__5270\,
            I => \U712_CYCLE_TERM.N_316_i_0_en\
        );

    \I__770\ : CEMux
    port map (
            O => \N__5267\,
            I => \N__5264\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__5264\,
            I => \U712_CYCLE_TERM.N_316_i_0_en_0\
        );

    \I__768\ : InMux
    port map (
            O => \N__5261\,
            I => \N__5258\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__5258\,
            I => \N__5254\
        );

    \I__766\ : InMux
    port map (
            O => \N__5257\,
            I => \N__5251\
        );

    \I__765\ : Odrv4
    port map (
            O => \N__5254\,
            I => \U712_BYTE_ENABLE.N_282_i\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5251\,
            I => \U712_BYTE_ENABLE.N_282_i\
        );

    \I__763\ : InMux
    port map (
            O => \N__5246\,
            I => \N__5243\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__5243\,
            I => \N__5240\
        );

    \I__761\ : Span12Mux_v
    port map (
            O => \N__5240\,
            I => \N__5237\
        );

    \I__760\ : Span12Mux_h
    port map (
            O => \N__5237\,
            I => \N__5234\
        );

    \I__759\ : Odrv12
    port map (
            O => \N__5234\,
            I => \A_c_4\
        );

    \I__758\ : InMux
    port map (
            O => \N__5231\,
            I => \N__5228\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__5228\,
            I => \N__5225\
        );

    \I__756\ : Span4Mux_v
    port map (
            O => \N__5225\,
            I => \N__5222\
        );

    \I__755\ : Sp12to4
    port map (
            O => \N__5222\,
            I => \N__5219\
        );

    \I__754\ : Span12Mux_h
    port map (
            O => \N__5219\,
            I => \N__5216\
        );

    \I__753\ : Odrv12
    port map (
            O => \N__5216\,
            I => \A_c_11\
        );

    \I__752\ : InMux
    port map (
            O => \N__5213\,
            I => \N__5210\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__5210\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\
        );

    \I__750\ : CascadeMux
    port map (
            O => \N__5207\,
            I => \U712_CHIP_RAM.N_15_cascade_\
        );

    \I__749\ : InMux
    port map (
            O => \N__5204\,
            I => \N__5201\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__5201\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_0_0\
        );

    \I__747\ : InMux
    port map (
            O => \N__5198\,
            I => \N__5195\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__5195\,
            I => \N__5192\
        );

    \I__745\ : Span4Mux_v
    port map (
            O => \N__5192\,
            I => \N__5189\
        );

    \I__744\ : Span4Mux_v
    port map (
            O => \N__5189\,
            I => \N__5186\
        );

    \I__743\ : Sp12to4
    port map (
            O => \N__5186\,
            I => \N__5183\
        );

    \I__742\ : Odrv12
    port map (
            O => \N__5183\,
            I => \A_c_5\
        );

    \I__741\ : InMux
    port map (
            O => \N__5180\,
            I => \N__5177\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__5177\,
            I => \N__5174\
        );

    \I__739\ : Span4Mux_v
    port map (
            O => \N__5174\,
            I => \N__5171\
        );

    \I__738\ : Span4Mux_h
    port map (
            O => \N__5171\,
            I => \N__5168\
        );

    \I__737\ : Sp12to4
    port map (
            O => \N__5168\,
            I => \N__5165\
        );

    \I__736\ : Odrv12
    port map (
            O => \N__5165\,
            I => \A_c_12\
        );

    \I__735\ : CascadeMux
    port map (
            O => \N__5162\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\
        );

    \I__734\ : InMux
    port map (
            O => \N__5159\,
            I => \N__5156\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__5156\,
            I => \N__5153\
        );

    \I__732\ : Odrv4
    port map (
            O => \N__5153\,
            I => \U712_CHIP_RAM.N_448\
        );

    \I__731\ : CascadeMux
    port map (
            O => \N__5150\,
            I => \U712_CHIP_RAM.N_345_cascade_\
        );

    \I__730\ : InMux
    port map (
            O => \N__5147\,
            I => \N__5144\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__5144\,
            I => \N__5141\
        );

    \I__728\ : Span12Mux_h
    port map (
            O => \N__5141\,
            I => \N__5138\
        );

    \I__727\ : Span12Mux_v
    port map (
            O => \N__5138\,
            I => \N__5135\
        );

    \I__726\ : Odrv12
    port map (
            O => \N__5135\,
            I => \A_c_2\
        );

    \I__725\ : InMux
    port map (
            O => \N__5132\,
            I => \N__5129\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__5129\,
            I => \N__5126\
        );

    \I__723\ : Span4Mux_v
    port map (
            O => \N__5126\,
            I => \N__5123\
        );

    \I__722\ : Sp12to4
    port map (
            O => \N__5123\,
            I => \N__5120\
        );

    \I__721\ : Odrv12
    port map (
            O => \N__5120\,
            I => \A_c_9\
        );

    \I__720\ : CascadeMux
    port map (
            O => \N__5117\,
            I => \U712_CHIP_RAM.N_288_cascade_\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__5114\,
            I => \U712_CHIP_RAM.N_372_cascade_\
        );

    \I__718\ : InMux
    port map (
            O => \N__5111\,
            I => \N__5108\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__5108\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0\
        );

    \I__716\ : CascadeMux
    port map (
            O => \N__5105\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_\
        );

    \I__715\ : CascadeMux
    port map (
            O => \N__5102\,
            I => \N__5099\
        );

    \I__714\ : InMux
    port map (
            O => \N__5099\,
            I => \N__5096\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__5096\,
            I => \N__5087\
        );

    \I__712\ : InMux
    port map (
            O => \N__5095\,
            I => \N__5084\
        );

    \I__711\ : InMux
    port map (
            O => \N__5094\,
            I => \N__5081\
        );

    \I__710\ : InMux
    port map (
            O => \N__5093\,
            I => \N__5076\
        );

    \I__709\ : InMux
    port map (
            O => \N__5092\,
            I => \N__5076\
        );

    \I__708\ : InMux
    port map (
            O => \N__5091\,
            I => \N__5071\
        );

    \I__707\ : InMux
    port map (
            O => \N__5090\,
            I => \N__5071\
        );

    \I__706\ : Odrv4
    port map (
            O => \N__5087\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__5084\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__5081\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__5076\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5071\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3\
        );

    \I__701\ : CascadeMux
    port map (
            O => \N__5060\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1_1_cascade_\
        );

    \I__700\ : CascadeMux
    port map (
            O => \N__5057\,
            I => \U712_CHIP_RAM.N_366_cascade_\
        );

    \I__699\ : CascadeMux
    port map (
            O => \N__5054\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_0_cascade_\
        );

    \I__698\ : IoInMux
    port map (
            O => \N__5051\,
            I => \N__5048\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__5048\,
            I => \N__5045\
        );

    \I__696\ : Span4Mux_s0_v
    port map (
            O => \N__5045\,
            I => \N__5042\
        );

    \I__695\ : Sp12to4
    port map (
            O => \N__5042\,
            I => \N__5038\
        );

    \I__694\ : InMux
    port map (
            O => \N__5041\,
            I => \N__5035\
        );

    \I__693\ : Span12Mux_h
    port map (
            O => \N__5038\,
            I => \N__5032\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__5035\,
            I => \N__5029\
        );

    \I__691\ : Odrv12
    port map (
            O => \N__5032\,
            I => \CONSTANT_ONE_NET\
        );

    \I__690\ : Odrv4
    port map (
            O => \N__5029\,
            I => \CONSTANT_ONE_NET\
        );

    \I__689\ : CascadeMux
    port map (
            O => \N__5024\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_cascade_\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__5021\,
            I => \N__5017\
        );

    \I__687\ : InMux
    port map (
            O => \N__5020\,
            I => \N__5012\
        );

    \I__686\ : InMux
    port map (
            O => \N__5017\,
            I => \N__5012\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__5012\,
            I => \N__5009\
        );

    \I__684\ : Odrv4
    port map (
            O => \N__5009\,
            I => \U712_CHIP_RAM.N_304\
        );

    \I__683\ : CascadeMux
    port map (
            O => \N__5006\,
            I => \U712_CHIP_RAM.N_62_cascade_\
        );

    \I__682\ : CascadeMux
    port map (
            O => \N__5003\,
            I => \N__4999\
        );

    \I__681\ : InMux
    port map (
            O => \N__5002\,
            I => \N__4995\
        );

    \I__680\ : InMux
    port map (
            O => \N__4999\,
            I => \N__4992\
        );

    \I__679\ : InMux
    port map (
            O => \N__4998\,
            I => \N__4989\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__4995\,
            I => \U712_CHIP_RAM.N_452\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__4992\,
            I => \U712_CHIP_RAM.N_452\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__4989\,
            I => \U712_CHIP_RAM.N_452\
        );

    \I__675\ : CascadeMux
    port map (
            O => \N__4982\,
            I => \U712_CHIP_RAM.N_452_cascade_\
        );

    \I__674\ : InMux
    port map (
            O => \N__4979\,
            I => \N__4974\
        );

    \I__673\ : InMux
    port map (
            O => \N__4978\,
            I => \N__4971\
        );

    \I__672\ : InMux
    port map (
            O => \N__4977\,
            I => \N__4968\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__4974\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__4971\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__4968\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__668\ : CascadeMux
    port map (
            O => \N__4961\,
            I => \U712_CHIP_RAM.N_11_cascade_\
        );

    \I__667\ : IoInMux
    port map (
            O => \N__4958\,
            I => \N__4955\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__4955\,
            I => \N__4952\
        );

    \I__665\ : Span4Mux_s0_h
    port map (
            O => \N__4952\,
            I => \N__4949\
        );

    \I__664\ : Sp12to4
    port map (
            O => \N__4949\,
            I => \N__4946\
        );

    \I__663\ : Span12Mux_v
    port map (
            O => \N__4946\,
            I => \N__4943\
        );

    \I__662\ : Span12Mux_h
    port map (
            O => \N__4943\,
            I => \N__4939\
        );

    \I__661\ : InMux
    port map (
            O => \N__4942\,
            I => \N__4936\
        );

    \I__660\ : Odrv12
    port map (
            O => \N__4939\,
            I => \CLK_EN_c\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__4936\,
            I => \CLK_EN_c\
        );

    \I__658\ : InMux
    port map (
            O => \N__4931\,
            I => \N__4927\
        );

    \I__657\ : InMux
    port map (
            O => \N__4930\,
            I => \N__4924\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__4927\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__4924\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__654\ : InMux
    port map (
            O => \N__4919\,
            I => \N__4907\
        );

    \I__653\ : InMux
    port map (
            O => \N__4918\,
            I => \N__4907\
        );

    \I__652\ : InMux
    port map (
            O => \N__4917\,
            I => \N__4907\
        );

    \I__651\ : InMux
    port map (
            O => \N__4916\,
            I => \N__4907\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__4907\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__649\ : InMux
    port map (
            O => \N__4904\,
            I => \N__4897\
        );

    \I__648\ : InMux
    port map (
            O => \N__4903\,
            I => \N__4897\
        );

    \I__647\ : InMux
    port map (
            O => \N__4902\,
            I => \N__4894\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__4897\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__4894\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__644\ : IoInMux
    port map (
            O => \N__4889\,
            I => \N__4886\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__4886\,
            I => \N__4883\
        );

    \I__642\ : Span4Mux_s0_h
    port map (
            O => \N__4883\,
            I => \N__4880\
        );

    \I__641\ : Sp12to4
    port map (
            O => \N__4880\,
            I => \N__4877\
        );

    \I__640\ : Span12Mux_v
    port map (
            O => \N__4877\,
            I => \N__4873\
        );

    \I__639\ : InMux
    port map (
            O => \N__4876\,
            I => \N__4870\
        );

    \I__638\ : Odrv12
    port map (
            O => \N__4873\,
            I => \TACK_OUTn\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__4870\,
            I => \TACK_OUTn\
        );

    \I__636\ : InMux
    port map (
            O => \N__4865\,
            I => \N__4862\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__4862\,
            I => \N__4859\
        );

    \I__634\ : Span4Mux_h
    port map (
            O => \N__4859\,
            I => \N__4856\
        );

    \I__633\ : Span4Mux_v
    port map (
            O => \N__4856\,
            I => \N__4853\
        );

    \I__632\ : Odrv4
    port map (
            O => \N__4853\,
            I => \TACK_EN_i_ess\
        );

    \I__631\ : InMux
    port map (
            O => \N__4850\,
            I => \N__4847\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4847\,
            I => \N__4844\
        );

    \I__629\ : Sp12to4
    port map (
            O => \N__4844\,
            I => \N__4841\
        );

    \I__628\ : Span12Mux_v
    port map (
            O => \N__4841\,
            I => \N__4838\
        );

    \I__627\ : Span12Mux_h
    port map (
            O => \N__4838\,
            I => \N__4835\
        );

    \I__626\ : Odrv12
    port map (
            O => \N__4835\,
            I => \A_c_18\
        );

    \I__625\ : InMux
    port map (
            O => \N__4832\,
            I => \N__4829\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__4829\,
            I => \N__4826\
        );

    \I__623\ : Sp12to4
    port map (
            O => \N__4826\,
            I => \N__4823\
        );

    \I__622\ : Span12Mux_v
    port map (
            O => \N__4823\,
            I => \N__4820\
        );

    \I__621\ : Span12Mux_h
    port map (
            O => \N__4820\,
            I => \N__4817\
        );

    \I__620\ : Odrv12
    port map (
            O => \N__4817\,
            I => \A_c_16\
        );

    \I__619\ : InMux
    port map (
            O => \N__4814\,
            I => \N__4810\
        );

    \I__618\ : InMux
    port map (
            O => \N__4813\,
            I => \N__4807\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__4810\,
            I => \U712_CHIP_RAM.N_489\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__4807\,
            I => \U712_CHIP_RAM.N_489\
        );

    \I__615\ : InMux
    port map (
            O => \N__4802\,
            I => \N__4799\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__4799\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\
        );

    \I__613\ : InMux
    port map (
            O => \N__4796\,
            I => \N__4793\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__4793\,
            I => \N__4789\
        );

    \I__611\ : InMux
    port map (
            O => \N__4792\,
            I => \N__4786\
        );

    \I__610\ : Span4Mux_h
    port map (
            O => \N__4789\,
            I => \N__4781\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__4786\,
            I => \N__4781\
        );

    \I__608\ : Span4Mux_v
    port map (
            O => \N__4781\,
            I => \N__4778\
        );

    \I__607\ : Sp12to4
    port map (
            O => \N__4778\,
            I => \N__4775\
        );

    \I__606\ : Span12Mux_h
    port map (
            O => \N__4775\,
            I => \N__4772\
        );

    \I__605\ : Span12Mux_v
    port map (
            O => \N__4772\,
            I => \N__4769\
        );

    \I__604\ : Odrv12
    port map (
            O => \N__4769\,
            I => \TSn_c\
        );

    \I__603\ : CascadeMux
    port map (
            O => \N__4766\,
            I => \N__4763\
        );

    \I__602\ : InMux
    port map (
            O => \N__4763\,
            I => \N__4760\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__4760\,
            I => \N__4757\
        );

    \I__600\ : Span12Mux_h
    port map (
            O => \N__4757\,
            I => \N__4754\
        );

    \I__599\ : Span12Mux_v
    port map (
            O => \N__4754\,
            I => \N__4751\
        );

    \I__598\ : Odrv12
    port map (
            O => \N__4751\,
            I => \RAMSPACEn_c\
        );

    \I__597\ : InMux
    port map (
            O => \N__4748\,
            I => \N__4744\
        );

    \I__596\ : InMux
    port map (
            O => \N__4747\,
            I => \N__4741\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__4744\,
            I => \N__4738\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__4741\,
            I => \N__4735\
        );

    \I__593\ : Span4Mux_v
    port map (
            O => \N__4738\,
            I => \N__4732\
        );

    \I__592\ : Span4Mux_v
    port map (
            O => \N__4735\,
            I => \N__4729\
        );

    \I__591\ : Sp12to4
    port map (
            O => \N__4732\,
            I => \N__4726\
        );

    \I__590\ : Span4Mux_h
    port map (
            O => \N__4729\,
            I => \N__4723\
        );

    \I__589\ : Span12Mux_h
    port map (
            O => \N__4726\,
            I => \N__4718\
        );

    \I__588\ : Sp12to4
    port map (
            O => \N__4723\,
            I => \N__4718\
        );

    \I__587\ : Span12Mux_v
    port map (
            O => \N__4718\,
            I => \N__4715\
        );

    \I__586\ : Odrv12
    port map (
            O => \N__4715\,
            I => \AWEn_c\
        );

    \I__585\ : IoInMux
    port map (
            O => \N__4712\,
            I => \N__4709\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__4709\,
            I => \N__4706\
        );

    \I__583\ : Span4Mux_s2_v
    port map (
            O => \N__4706\,
            I => \N__4703\
        );

    \I__582\ : Span4Mux_v
    port map (
            O => \N__4703\,
            I => \N__4700\
        );

    \I__581\ : Span4Mux_v
    port map (
            O => \N__4700\,
            I => \N__4696\
        );

    \I__580\ : InMux
    port map (
            O => \N__4699\,
            I => \N__4693\
        );

    \I__579\ : Odrv4
    port map (
            O => \N__4696\,
            I => \DBDIR_c\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__4693\,
            I => \DBDIR_c\
        );

    \I__577\ : InMux
    port map (
            O => \N__4688\,
            I => \N__4684\
        );

    \I__576\ : InMux
    port map (
            O => \N__4687\,
            I => \N__4681\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__4684\,
            I => \U712_REG_SM.STATE_COUNT_RNI4BRHZ0Z_3\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__4681\,
            I => \U712_REG_SM.STATE_COUNT_RNI4BRHZ0Z_3\
        );

    \I__573\ : InMux
    port map (
            O => \N__4676\,
            I => \N__4673\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__4673\,
            I => \U712_REG_SM.N_400\
        );

    \I__571\ : InMux
    port map (
            O => \N__4670\,
            I => \N__4667\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__4667\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_12_0\
        );

    \I__569\ : IoInMux
    port map (
            O => \N__4664\,
            I => \N__4661\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__4661\,
            I => \N__4658\
        );

    \I__567\ : IoSpan4Mux
    port map (
            O => \N__4658\,
            I => \N__4655\
        );

    \I__566\ : Sp12to4
    port map (
            O => \N__4655\,
            I => \N__4652\
        );

    \I__565\ : Span12Mux_s6_v
    port map (
            O => \N__4652\,
            I => \N__4649\
        );

    \I__564\ : Span12Mux_v
    port map (
            O => \N__4649\,
            I => \N__4645\
        );

    \I__563\ : InMux
    port map (
            O => \N__4648\,
            I => \N__4642\
        );

    \I__562\ : Odrv12
    port map (
            O => \N__4645\,
            I => \LATCH_CLK_c\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__4642\,
            I => \LATCH_CLK_c\
        );

    \I__560\ : InMux
    port map (
            O => \N__4637\,
            I => \N__4633\
        );

    \I__559\ : InMux
    port map (
            O => \N__4636\,
            I => \N__4630\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__4633\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__4630\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__556\ : InMux
    port map (
            O => \N__4625\,
            I => \N__4622\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__4622\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\
        );

    \I__554\ : CascadeMux
    port map (
            O => \N__4619\,
            I => \U712_CHIP_RAM.N_361_cascade_\
        );

    \I__553\ : CascadeMux
    port map (
            O => \N__4616\,
            I => \N__4613\
        );

    \I__552\ : InMux
    port map (
            O => \N__4613\,
            I => \N__4610\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__4610\,
            I => \N__4607\
        );

    \I__550\ : Span4Mux_v
    port map (
            O => \N__4607\,
            I => \N__4604\
        );

    \I__549\ : Sp12to4
    port map (
            O => \N__4604\,
            I => \N__4601\
        );

    \I__548\ : Span12Mux_h
    port map (
            O => \N__4601\,
            I => \N__4598\
        );

    \I__547\ : Span12Mux_v
    port map (
            O => \N__4598\,
            I => \N__4595\
        );

    \I__546\ : Odrv12
    port map (
            O => \N__4595\,
            I => \A_c_20\
        );

    \I__545\ : InMux
    port map (
            O => \N__4592\,
            I => \N__4588\
        );

    \I__544\ : InMux
    port map (
            O => \N__4591\,
            I => \N__4585\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4588\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__4585\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__541\ : CascadeMux
    port map (
            O => \N__4580\,
            I => \U712_CHIP_RAM.N_416_cascade_\
        );

    \I__540\ : CascadeMux
    port map (
            O => \N__4577\,
            I => \U712_CHIP_RAM.BANK0_RNOZ0Z_0_cascade_\
        );

    \I__539\ : InMux
    port map (
            O => \N__4574\,
            I => \N__4571\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__4571\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_i_i_0\
        );

    \I__537\ : IoInMux
    port map (
            O => \N__4568\,
            I => \N__4565\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4565\,
            I => \N__4562\
        );

    \I__535\ : Span4Mux_s3_v
    port map (
            O => \N__4562\,
            I => \N__4559\
        );

    \I__534\ : Span4Mux_v
    port map (
            O => \N__4559\,
            I => \N__4556\
        );

    \I__533\ : Span4Mux_v
    port map (
            O => \N__4556\,
            I => \N__4553\
        );

    \I__532\ : Span4Mux_h
    port map (
            O => \N__4553\,
            I => \N__4549\
        );

    \I__531\ : InMux
    port map (
            O => \N__4552\,
            I => \N__4546\
        );

    \I__530\ : Odrv4
    port map (
            O => \N__4549\,
            I => \BANK0_c\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__4546\,
            I => \BANK0_c\
        );

    \I__528\ : CascadeMux
    port map (
            O => \N__4541\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3_cascade_\
        );

    \I__527\ : CascadeMux
    port map (
            O => \N__4538\,
            I => \U712_CHIP_RAM.N_410_cascade_\
        );

    \I__526\ : IoInMux
    port map (
            O => \N__4535\,
            I => \N__4532\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__4532\,
            I => \N__4529\
        );

    \I__524\ : IoSpan4Mux
    port map (
            O => \N__4529\,
            I => \N__4526\
        );

    \I__523\ : Span4Mux_s3_h
    port map (
            O => \N__4526\,
            I => \N__4522\
        );

    \I__522\ : InMux
    port map (
            O => \N__4525\,
            I => \N__4519\
        );

    \I__521\ : Span4Mux_h
    port map (
            O => \N__4522\,
            I => \N__4516\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__4519\,
            I => \N__4513\
        );

    \I__519\ : Sp12to4
    port map (
            O => \N__4516\,
            I => \N__4510\
        );

    \I__518\ : Span4Mux_v
    port map (
            O => \N__4513\,
            I => \N__4507\
        );

    \I__517\ : Span12Mux_h
    port map (
            O => \N__4510\,
            I => \N__4502\
        );

    \I__516\ : Sp12to4
    port map (
            O => \N__4507\,
            I => \N__4502\
        );

    \I__515\ : Span12Mux_h
    port map (
            O => \N__4502\,
            I => \N__4499\
        );

    \I__514\ : Span12Mux_v
    port map (
            O => \N__4499\,
            I => \N__4496\
        );

    \I__513\ : Odrv12
    port map (
            O => \N__4496\,
            I => \C3_c\
        );

    \I__512\ : CEMux
    port map (
            O => \N__4493\,
            I => \N__4490\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__4490\,
            I => \N__4487\
        );

    \I__510\ : Odrv12
    port map (
            O => \N__4487\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0\
        );

    \I__509\ : InMux
    port map (
            O => \N__4484\,
            I => \N__4481\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__4481\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0\
        );

    \I__507\ : InMux
    port map (
            O => \N__4478\,
            I => \N__4475\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__4475\,
            I => \U712_CHIP_RAM.N_409\
        );

    \I__505\ : InMux
    port map (
            O => \N__4472\,
            I => \N__4468\
        );

    \I__504\ : InMux
    port map (
            O => \N__4471\,
            I => \N__4465\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4468\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0_1\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__4465\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0_1\
        );

    \I__501\ : CascadeMux
    port map (
            O => \N__4460\,
            I => \U712_CHIP_RAM.N_489_cascade_\
        );

    \I__500\ : CascadeMux
    port map (
            O => \N__4457\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_0_cascade_\
        );

    \I__499\ : CascadeMux
    port map (
            O => \N__4454\,
            I => \U712_REG_SM.N_346_cascade_\
        );

    \I__498\ : InMux
    port map (
            O => \N__4451\,
            I => \N__4447\
        );

    \I__497\ : InMux
    port map (
            O => \N__4450\,
            I => \N__4443\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__4447\,
            I => \N__4437\
        );

    \I__495\ : InMux
    port map (
            O => \N__4446\,
            I => \N__4434\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4443\,
            I => \N__4431\
        );

    \I__493\ : InMux
    port map (
            O => \N__4442\,
            I => \N__4424\
        );

    \I__492\ : InMux
    port map (
            O => \N__4441\,
            I => \N__4424\
        );

    \I__491\ : InMux
    port map (
            O => \N__4440\,
            I => \N__4424\
        );

    \I__490\ : Odrv4
    port map (
            O => \N__4437\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4434\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__488\ : Odrv4
    port map (
            O => \N__4431\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__4424\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__486\ : InMux
    port map (
            O => \N__4415\,
            I => \N__4409\
        );

    \I__485\ : InMux
    port map (
            O => \N__4414\,
            I => \N__4400\
        );

    \I__484\ : InMux
    port map (
            O => \N__4413\,
            I => \N__4400\
        );

    \I__483\ : InMux
    port map (
            O => \N__4412\,
            I => \N__4400\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__4409\,
            I => \N__4397\
        );

    \I__481\ : InMux
    port map (
            O => \N__4408\,
            I => \N__4394\
        );

    \I__480\ : InMux
    port map (
            O => \N__4407\,
            I => \N__4391\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4400\,
            I => \N__4388\
        );

    \I__478\ : Span4Mux_h
    port map (
            O => \N__4397\,
            I => \N__4385\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__4394\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__4391\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__475\ : Odrv4
    port map (
            O => \N__4388\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__474\ : Odrv4
    port map (
            O => \N__4385\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__473\ : CascadeMux
    port map (
            O => \N__4376\,
            I => \U712_REG_SM.STATE_COUNT_srsts_i_i_0_o2_0_1_3_cascade_\
        );

    \I__472\ : InMux
    port map (
            O => \N__4373\,
            I => \N__4370\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__4370\,
            I => \N__4366\
        );

    \I__470\ : InMux
    port map (
            O => \N__4369\,
            I => \N__4363\
        );

    \I__469\ : Odrv4
    port map (
            O => \N__4366\,
            I => \U712_REG_SM.N_342\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__4363\,
            I => \U712_REG_SM.N_342\
        );

    \I__467\ : InMux
    port map (
            O => \N__4358\,
            I => \N__4355\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__4355\,
            I => \U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0_0\
        );

    \I__465\ : CascadeMux
    port map (
            O => \N__4352\,
            I => \N__4349\
        );

    \I__464\ : InMux
    port map (
            O => \N__4349\,
            I => \N__4346\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__4346\,
            I => \U712_REG_SM.N_106\
        );

    \I__462\ : InMux
    port map (
            O => \N__4343\,
            I => \N__4340\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__4340\,
            I => \U712_REG_SM.N_379\
        );

    \I__460\ : InMux
    port map (
            O => \N__4337\,
            I => \N__4333\
        );

    \I__459\ : InMux
    port map (
            O => \N__4336\,
            I => \N__4330\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__4333\,
            I => \N__4326\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__4330\,
            I => \N__4323\
        );

    \I__456\ : InMux
    port map (
            O => \N__4329\,
            I => \N__4320\
        );

    \I__455\ : Span4Mux_v
    port map (
            O => \N__4326\,
            I => \N__4317\
        );

    \I__454\ : Span4Mux_v
    port map (
            O => \N__4323\,
            I => \N__4312\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__4320\,
            I => \N__4312\
        );

    \I__452\ : Span4Mux_v
    port map (
            O => \N__4317\,
            I => \N__4309\
        );

    \I__451\ : Span4Mux_v
    port map (
            O => \N__4312\,
            I => \N__4306\
        );

    \I__450\ : Sp12to4
    port map (
            O => \N__4309\,
            I => \N__4301\
        );

    \I__449\ : Sp12to4
    port map (
            O => \N__4306\,
            I => \N__4301\
        );

    \I__448\ : Span12Mux_h
    port map (
            O => \N__4301\,
            I => \N__4298\
        );

    \I__447\ : Odrv12
    port map (
            O => \N__4298\,
            I => \DBRn_c\
        );

    \I__446\ : IoInMux
    port map (
            O => \N__4295\,
            I => \N__4292\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__4292\,
            I => \N__4289\
        );

    \I__444\ : Span4Mux_s2_v
    port map (
            O => \N__4289\,
            I => \N__4285\
        );

    \I__443\ : InMux
    port map (
            O => \N__4288\,
            I => \N__4282\
        );

    \I__442\ : Sp12to4
    port map (
            O => \N__4285\,
            I => \N__4279\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__4282\,
            I => \N__4275\
        );

    \I__440\ : Span12Mux_s9_h
    port map (
            O => \N__4279\,
            I => \N__4272\
        );

    \I__439\ : CascadeMux
    port map (
            O => \N__4278\,
            I => \N__4269\
        );

    \I__438\ : Span4Mux_v
    port map (
            O => \N__4275\,
            I => \N__4266\
        );

    \I__437\ : Span12Mux_v
    port map (
            O => \N__4272\,
            I => \N__4263\
        );

    \I__436\ : InMux
    port map (
            O => \N__4269\,
            I => \N__4260\
        );

    \I__435\ : Span4Mux_v
    port map (
            O => \N__4266\,
            I => \N__4257\
        );

    \I__434\ : Odrv12
    port map (
            O => \N__4263\,
            I => \REGENn_c\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__4260\,
            I => \REGENn_c\
        );

    \I__432\ : Odrv4
    port map (
            O => \N__4257\,
            I => \REGENn_c\
        );

    \I__431\ : IoInMux
    port map (
            O => \N__4250\,
            I => \N__4247\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__4247\,
            I => \N__4244\
        );

    \I__429\ : Odrv12
    port map (
            O => \N__4244\,
            I => \VBENn_c\
        );

    \I__428\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4235\
        );

    \I__427\ : InMux
    port map (
            O => \N__4240\,
            I => \N__4235\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__4235\,
            I => \U712_REG_SM.N_319\
        );

    \I__425\ : IoInMux
    port map (
            O => \N__4232\,
            I => \N__4229\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__4229\,
            I => \N__4226\
        );

    \I__423\ : Span4Mux_s1_v
    port map (
            O => \N__4226\,
            I => \N__4223\
        );

    \I__422\ : Span4Mux_v
    port map (
            O => \N__4223\,
            I => \N__4220\
        );

    \I__421\ : Sp12to4
    port map (
            O => \N__4220\,
            I => \N__4217\
        );

    \I__420\ : Span12Mux_h
    port map (
            O => \N__4217\,
            I => \N__4214\
        );

    \I__419\ : Span12Mux_v
    port map (
            O => \N__4214\,
            I => \N__4210\
        );

    \I__418\ : InMux
    port map (
            O => \N__4213\,
            I => \N__4207\
        );

    \I__417\ : Odrv12
    port map (
            O => \N__4210\,
            I => \ASn_c\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__4207\,
            I => \ASn_c\
        );

    \I__415\ : CascadeMux
    port map (
            O => \N__4202\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_cascade_\
        );

    \I__414\ : InMux
    port map (
            O => \N__4199\,
            I => \N__4196\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__4196\,
            I => \N__4193\
        );

    \I__412\ : Span4Mux_v
    port map (
            O => \N__4193\,
            I => \N__4190\
        );

    \I__411\ : Odrv4
    port map (
            O => \N__4190\,
            I => \DBRn_c_i\
        );

    \I__410\ : CascadeMux
    port map (
            O => \N__4187\,
            I => \N__4181\
        );

    \I__409\ : InMux
    port map (
            O => \N__4186\,
            I => \N__4177\
        );

    \I__408\ : InMux
    port map (
            O => \N__4185\,
            I => \N__4174\
        );

    \I__407\ : InMux
    port map (
            O => \N__4184\,
            I => \N__4171\
        );

    \I__406\ : InMux
    port map (
            O => \N__4181\,
            I => \N__4166\
        );

    \I__405\ : InMux
    port map (
            O => \N__4180\,
            I => \N__4166\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__4177\,
            I => \U712_REG_SM.C1_SYNC_RNIAS4F1Z0Z_1\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__4174\,
            I => \U712_REG_SM.C1_SYNC_RNIAS4F1Z0Z_1\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__4171\,
            I => \U712_REG_SM.C1_SYNC_RNIAS4F1Z0Z_1\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__4166\,
            I => \U712_REG_SM.C1_SYNC_RNIAS4F1Z0Z_1\
        );

    \I__400\ : InMux
    port map (
            O => \N__4157\,
            I => \N__4154\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__4154\,
            I => \N__4151\
        );

    \I__398\ : Odrv4
    port map (
            O => \N__4151\,
            I => \U712_REG_SM.N_348\
        );

    \I__397\ : CascadeMux
    port map (
            O => \N__4148\,
            I => \DBRn_c_i_cascade_\
        );

    \I__396\ : IoInMux
    port map (
            O => \N__4145\,
            I => \N__4142\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__4142\,
            I => \N__4139\
        );

    \I__394\ : IoSpan4Mux
    port map (
            O => \N__4139\,
            I => \N__4136\
        );

    \I__393\ : Span4Mux_s3_h
    port map (
            O => \N__4136\,
            I => \N__4133\
        );

    \I__392\ : Span4Mux_h
    port map (
            O => \N__4133\,
            I => \N__4130\
        );

    \I__391\ : Odrv4
    port map (
            O => \N__4130\,
            I => \DBRn_c_i_0\
        );

    \I__390\ : InMux
    port map (
            O => \N__4127\,
            I => \N__4124\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__4124\,
            I => \N__4120\
        );

    \I__388\ : IoInMux
    port map (
            O => \N__4123\,
            I => \N__4117\
        );

    \I__387\ : Span4Mux_v
    port map (
            O => \N__4120\,
            I => \N__4114\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__4117\,
            I => \N__4111\
        );

    \I__385\ : Sp12to4
    port map (
            O => \N__4114\,
            I => \N__4108\
        );

    \I__384\ : IoSpan4Mux
    port map (
            O => \N__4111\,
            I => \N__4105\
        );

    \I__383\ : Span12Mux_h
    port map (
            O => \N__4108\,
            I => \N__4102\
        );

    \I__382\ : IoSpan4Mux
    port map (
            O => \N__4105\,
            I => \N__4099\
        );

    \I__381\ : Span12Mux_v
    port map (
            O => \N__4102\,
            I => \N__4096\
        );

    \I__380\ : IoSpan4Mux
    port map (
            O => \N__4099\,
            I => \N__4093\
        );

    \I__379\ : Odrv12
    port map (
            O => \N__4096\,
            I => \C1_c\
        );

    \I__378\ : Odrv4
    port map (
            O => \N__4093\,
            I => \C1_c\
        );

    \I__377\ : InMux
    port map (
            O => \N__4088\,
            I => \N__4082\
        );

    \I__376\ : InMux
    port map (
            O => \N__4087\,
            I => \N__4082\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__4082\,
            I => \U712_REG_SM.REG_CYCLE_START_RNITO6SZ0Z1\
        );

    \I__374\ : InMux
    port map (
            O => \N__4079\,
            I => \N__4075\
        );

    \I__373\ : InMux
    port map (
            O => \N__4078\,
            I => \N__4072\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__4075\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__4072\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__370\ : IoInMux
    port map (
            O => \N__4067\,
            I => \N__4064\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__4064\,
            I => \N__4061\
        );

    \I__368\ : Span12Mux_s5_h
    port map (
            O => \N__4061\,
            I => \N__4058\
        );

    \I__367\ : Odrv12
    port map (
            O => \N__4058\,
            I => \N_1062_i\
        );

    \I__366\ : IoInMux
    port map (
            O => \N__4055\,
            I => \N__4052\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__4052\,
            I => \N__4049\
        );

    \I__364\ : Span4Mux_s3_v
    port map (
            O => \N__4049\,
            I => \N__4046\
        );

    \I__363\ : Span4Mux_h
    port map (
            O => \N__4046\,
            I => \N__4043\
        );

    \I__362\ : Odrv4
    port map (
            O => \N__4043\,
            I => \CLK80_PLL_i_i\
        );

    \I__361\ : CascadeMux
    port map (
            O => \N__4040\,
            I => \N__4037\
        );

    \I__360\ : InMux
    port map (
            O => \N__4037\,
            I => \N__4034\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__4034\,
            I => \N__4031\
        );

    \I__358\ : Span4Mux_h
    port map (
            O => \N__4031\,
            I => \N__4028\
        );

    \I__357\ : Span4Mux_v
    port map (
            O => \N__4028\,
            I => \N__4025\
        );

    \I__356\ : Span4Mux_v
    port map (
            O => \N__4025\,
            I => \N__4022\
        );

    \I__355\ : Odrv4
    port map (
            O => \N__4022\,
            I => \REGSPACEn_c\
        );

    \I__354\ : InMux
    port map (
            O => \N__4019\,
            I => \N__4014\
        );

    \I__353\ : InMux
    port map (
            O => \N__4018\,
            I => \N__4009\
        );

    \I__352\ : InMux
    port map (
            O => \N__4017\,
            I => \N__4009\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__4014\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__4009\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__349\ : IoInMux
    port map (
            O => \N__4004\,
            I => \N__4001\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__4001\,
            I => \N__3998\
        );

    \I__347\ : IoSpan4Mux
    port map (
            O => \N__3998\,
            I => \N__3995\
        );

    \I__346\ : Span4Mux_s2_v
    port map (
            O => \N__3995\,
            I => \N__3992\
        );

    \I__345\ : Sp12to4
    port map (
            O => \N__3992\,
            I => \N__3989\
        );

    \I__344\ : Span12Mux_v
    port map (
            O => \N__3989\,
            I => \N__3986\
        );

    \I__343\ : Odrv12
    port map (
            O => \N__3986\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__6732\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__6729\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            I => \N__6730\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            I => \N__6731\
        );

    \INVU712_CHIP_RAM.DMA_A20C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A20C_net\,
            I => \N__6734\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_7_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8264\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4123\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4145\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4535\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \TACKn_obuft_RNO_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4865\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_1062_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_3_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9821\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001101"
        )
    port map (
            in0 => \N__4792\,
            in1 => \N__4019\,
            in2 => \N__4040\,
            in3 => \N__8126\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9810\,
            ce => 'H',
            sr => \N__10806\
        );

    \U712_REG_SM.REG_CYCLE_START_RNITO6S1_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4017\,
            in2 => \_gnd_net_\,
            in3 => \N__4180\,
            lcout => \U712_REG_SM.REG_CYCLE_START_RNITO6SZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011110111"
        )
    port map (
            in0 => \N__4018\,
            in1 => \N__4078\,
            in2 => \N__4187\,
            in3 => \N__4408\,
            lcout => \U712_REG_SM.N_348\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000110010"
        )
    port map (
            in0 => \N__5748\,
            in1 => \N__5722\,
            in2 => \N__5795\,
            in3 => \N__4186\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9817\,
            ce => 'H',
            sr => \N__10805\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__6004\,
            in1 => \N__5884\,
            in2 => \N__6755\,
            in3 => \N__4157\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9817\,
            ce => 'H',
            sr => \N__10805\
        );

    \U712_REG_SM.STATE_COUNT_RNIBMB91_1_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__4407\,
            in1 => \N__5885\,
            in2 => \N__6008\,
            in3 => \N__6747\,
            lcout => \U712_REG_SM.N_319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBRn_ibuf_RNIBAB_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4337\,
            lcout => \DBRn_c_i\,
            ltout => \DBRn_c_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4148\,
            in3 => \N__10824\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001000000000"
        )
    port map (
            in0 => \N__4451\,
            in1 => \N__4373\,
            in2 => \N__5755\,
            in3 => \N__4185\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9808\,
            ce => 'H',
            sr => \N__10800\
        );

    \U712_REG_SM.C1_SYNC_0_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4127\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9811\,
            ce => 'H',
            sr => \N__10793\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__5790\,
            in1 => \N__4688\,
            in2 => \N__5723\,
            in3 => \N__4088\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9811\,
            ce => 'H',
            sr => \N__10793\
        );

    \U712_REG_SM.REGENn_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110101011111010"
        )
    port map (
            in0 => \N__5815\,
            in1 => \N__4087\,
            in2 => \N__4278\,
            in3 => \N__4079\,
            lcout => \REGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9811\,
            ce => 'H',
            sr => \N__10793\
        );

    \U712_REG_SM.C1_SYNC_RNIAS4F1_1_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__5883\,
            in1 => \N__6003\,
            in2 => \N__5957\,
            in3 => \N__5914\,
            lcout => \U712_REG_SM.C1_SYNC_RNIAS4F1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__4446\,
            in1 => \N__4369\,
            in2 => \_gnd_net_\,
            in3 => \N__4240\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9814\,
            ce => 'H',
            sr => \N__10786\
        );

    \U712_REG_SM.ASn_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__4213\,
            in1 => \N__5822\,
            in2 => \_gnd_net_\,
            in3 => \N__4241\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9814\,
            ce => 'H',
            sr => \N__10786\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__7428\,
            in1 => \N__6151\,
            in2 => \N__5459\,
            in3 => \N__4478\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011101011111010"
        )
    port map (
            in0 => \N__6198\,
            in1 => \N__5573\,
            in2 => \N__4202\,
            in3 => \N__8990\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9803\,
            ce => 'H',
            sr => \N__10801\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_0_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111010"
        )
    port map (
            in0 => \N__4472\,
            in1 => \N__7427\,
            in2 => \N__6152\,
            in3 => \N__5455\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_A20_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__11153\,
            in1 => \N__4199\,
            in2 => \N__11075\,
            in3 => \N__4592\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A20C_net\,
            ce => 'H',
            sr => \N__10794\
        );

    \U712_REG_SM.STATE_COUNT_RNI4BRH_3_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4415\,
            in1 => \N__5747\,
            in2 => \_gnd_net_\,
            in3 => \N__4450\,
            lcout => \U712_REG_SM.STATE_COUNT_RNI4BRHZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000001"
        )
    port map (
            in0 => \N__7869\,
            in1 => \N__7969\,
            in2 => \N__7150\,
            in3 => \N__7219\,
            lcout => \U712_CHIP_RAM.N_347\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4184\,
            in1 => \N__4413\,
            in2 => \_gnd_net_\,
            in3 => \N__4441\,
            lcout => \U712_REG_SM.N_400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__5870\,
            in1 => \N__6562\,
            in2 => \_gnd_net_\,
            in3 => \N__5793\,
            lcout => \U712_REG_SM.N_106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_3_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111101110"
        )
    port map (
            in0 => \N__5991\,
            in1 => \N__4440\,
            in2 => \_gnd_net_\,
            in3 => \N__5869\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_346_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_2_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110101"
        )
    port map (
            in0 => \N__4412\,
            in1 => \N__5919\,
            in2 => \N__4454\,
            in3 => \N__5953\,
            lcout => \U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_1_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000010001"
        )
    port map (
            in0 => \N__5794\,
            in1 => \N__4442\,
            in2 => \N__6754\,
            in3 => \N__4414\,
            lcout => \U712_REG_SM.N_379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIS63V_1_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__5948\,
            in1 => \N__5915\,
            in2 => \N__5669\,
            in3 => \N__4930\,
            lcout => OPEN,
            ltout => \U712_REG_SM.STATE_COUNT_srsts_i_i_0_o2_0_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI35EO1_1_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5871\,
            in2 => \N__4376\,
            in3 => \N__5992\,
            lcout => \U712_REG_SM.N_342\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001011"
        )
    port map (
            in0 => \N__10357\,
            in1 => \N__4358\,
            in2 => \N__4352\,
            in3 => \N__4343\,
            lcout => \DS_ENm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9812\,
            ce => 'H',
            sr => \N__10779\
        );

    \DBR_SYNC_0_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4336\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9815\,
            ce => 'H',
            sr => \N__10775\
        );

    \U712_REG_SM.REG_CYCLE_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__4329\,
            in1 => \N__8386\,
            in2 => \_gnd_net_\,
            in3 => \N__4288\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10889\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_0_a3_0_a2_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8125\,
            in2 => \_gnd_net_\,
            in3 => \N__9638\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__4747\,
            in1 => \N__6554\,
            in2 => \_gnd_net_\,
            in3 => \N__7568\,
            lcout => \WRITE_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9794\,
            ce => \N__4493\,
            sr => \N__10802\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10826\,
            in2 => \_gnd_net_\,
            in3 => \N__4977\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10825\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4484\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNISNC52_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__7381\,
            in1 => \N__7740\,
            in2 => \N__7112\,
            in3 => \N__7245\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNO_1_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7247\,
            in1 => \N__6377\,
            in2 => \_gnd_net_\,
            in3 => \N__5092\,
            lcout => \U712_CHIP_RAM.N_409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI71B91_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101100"
        )
    port map (
            in0 => \N__7605\,
            in1 => \N__7950\,
            in2 => \N__7113\,
            in3 => \N__7246\,
            lcout => \U712_CHIP_RAM.N_304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIR9VE1_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__5617\,
            in1 => \N__6881\,
            in2 => \N__7567\,
            in3 => \N__5671\,
            lcout => \U712_CHIP_RAM.N_489\,
            ltout => \U712_CHIP_RAM.N_489_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNO_1_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__4471\,
            in1 => \N__4998\,
            in2 => \N__4460\,
            in3 => \N__5446\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__7951\,
            in1 => \N__7079\,
            in2 => \N__4457\,
            in3 => \N__5093\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_3_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__7970\,
            in1 => \N__7269\,
            in2 => \N__7138\,
            in3 => \N__5095\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_361_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_1_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__6147\,
            in1 => \N__7434\,
            in2 => \N__4619\,
            in3 => \N__5444\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_i_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_2_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11071\,
            in1 => \N__4813\,
            in2 => \N__4616\,
            in3 => \N__5567\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_416_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_0_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__5568\,
            in1 => \N__4591\,
            in2 => \N__4580\,
            in3 => \N__7562\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.BANK0_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__4552\,
            in1 => \N__4978\,
            in2 => \N__4577\,
            in3 => \N__4574\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9804\,
            ce => 'H',
            sr => \N__10787\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_3_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7868\,
            in1 => \N__7432\,
            in2 => \_gnd_net_\,
            in3 => \N__5442\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_3_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7268\,
            in2 => \N__4541\,
            in3 => \N__6375\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_410_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__6146\,
            in1 => \N__7433\,
            in2 => \N__4538\,
            in3 => \N__5443\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_1_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5872\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9807\,
            ce => 'H',
            sr => \N__10780\
        );

    \U712_REG_SM.C3_SYNC_0_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4525\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9807\,
            ce => 'H',
            sr => \N__10780\
        );

    \U712_REG_SM.REG_TACK_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__4687\,
            in1 => \N__4676\,
            in2 => \N__5699\,
            in3 => \N__5353\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9807\,
            ce => 'H',
            sr => \N__10780\
        );

    \U712_REG_SM.C1_SYNC_1_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5920\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9807\,
            ce => 'H',
            sr => \N__10780\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__4648\,
            in1 => \N__5684\,
            in2 => \_gnd_net_\,
            in3 => \N__4670\,
            lcout => \LATCH_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9807\,
            ce => 'H',
            sr => \N__10780\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4902\,
            in2 => \_gnd_net_\,
            in3 => \N__4636\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4637\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9813\,
            ce => 'H',
            sr => \N__10770\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000001010"
        )
    port map (
            in0 => \N__5290\,
            in1 => \N__8481\,
            in2 => \N__5330\,
            in3 => \N__4919\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9813\,
            ce => 'H',
            sr => \N__10770\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__4917\,
            in1 => \_gnd_net_\,
            in2 => \N__8483\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9813\,
            ce => 'H',
            sr => \N__10770\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__4625\,
            in1 => \N__5326\,
            in2 => \N__5309\,
            in3 => \N__4916\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9813\,
            ce => 'H',
            sr => \N__10770\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4904\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9813\,
            ce => 'H',
            sr => \N__10770\
        );

    \DBR_SYNC_1_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4931\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9813\,
            ce => 'H',
            sr => \N__10770\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111000100"
        )
    port map (
            in0 => \N__4918\,
            in1 => \N__4876\,
            in2 => \N__8482\,
            in3 => \N__4903\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9813\,
            ce => 'H',
            sr => \N__10770\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__5325\,
            in1 => \N__8295\,
            in2 => \_gnd_net_\,
            in3 => \N__5291\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9816\,
            ce => \N__5267\,
            sr => \N__10767\
        );

    \CONSTANT_ONE_LUT4_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4850\,
            in1 => \N__4832\,
            in2 => \_gnd_net_\,
            in3 => \N__9464\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__4814\,
            in1 => \N__5572\,
            in2 => \N__9682\,
            in3 => \N__4802\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9792\,
            ce => 'H',
            sr => \N__10795\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011100000101"
        )
    port map (
            in0 => \N__4796\,
            in1 => \N__9637\,
            in2 => \N__4766\,
            in3 => \N__5619\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9792\,
            ce => 'H',
            sr => \N__10795\
        );

    \U712_CHIP_RAM.DBDIR_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011101010101010"
        )
    port map (
            in0 => \N__4699\,
            in1 => \N__4748\,
            in2 => \N__7566\,
            in3 => \N__5002\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9792\,
            ce => 'H',
            sr => \N__10795\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110011"
        )
    port map (
            in0 => \N__5091\,
            in1 => \N__8392\,
            in2 => \N__5483\,
            in3 => \N__5020\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111101100110"
        )
    port map (
            in0 => \N__5041\,
            in1 => \N__7125\,
            in2 => \N__5024\,
            in3 => \N__6842\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9795\,
            ce => \N__6796\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI49DCG_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111011101"
        )
    port map (
            in0 => \N__8390\,
            in1 => \N__5534\,
            in2 => \N__5021\,
            in3 => \N__5090\,
            lcout => \U712_CHIP_RAM.N_62\,
            ltout => \U712_CHIP_RAM.N_62_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__4979\,
            in1 => \N__6671\,
            in2 => \N__5006\,
            in3 => \N__8391\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9795\,
            ce => \N__6796\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIGGM16_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101011111"
        )
    port map (
            in0 => \N__7475\,
            in1 => \N__5672\,
            in2 => \N__5003\,
            in3 => \N__5618\,
            lcout => \U712_CHIP_RAM.N_434_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_3_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7395\,
            in1 => \N__6357\,
            in2 => \N__7867\,
            in3 => \N__5454\,
            lcout => \U712_CHIP_RAM.N_452\,
            ltout => \U712_CHIP_RAM.N_452_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIQ6QH5_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7545\,
            in2 => \N__4982\,
            in3 => \N__5159\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__7098\,
            in1 => \N__5384\,
            in2 => \N__7443\,
            in3 => \N__5365\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010001110101111"
        )
    port map (
            in0 => \N__4942\,
            in1 => \N__9681\,
            in2 => \N__4961\,
            in3 => \N__7973\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9800\,
            ce => 'H',
            sr => \N__10781\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4GV43_2_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__7972\,
            in1 => \N__7871\,
            in2 => \_gnd_net_\,
            in3 => \N__5445\,
            lcout => \U712_CHIP_RAM.N_11_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__5585\,
            in1 => \N__8388\,
            in2 => \N__5102\,
            in3 => \N__5111\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7202\,
            in2 => \_gnd_net_\,
            in3 => \N__6066\,
            lcout => \U712_CHIP_RAM.N_288\,
            ltout => \U712_CHIP_RAM.N_288_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_2_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000010"
        )
    port map (
            in0 => \N__5801\,
            in1 => \N__7971\,
            in2 => \N__5117\,
            in3 => \N__7097\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_372_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIADE59_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__8389\,
            in1 => \N__5498\,
            in2 => \N__5114\,
            in3 => \N__6067\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNILV2DI_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__5584\,
            in1 => \N__8387\,
            in2 => \N__5105\,
            in3 => \N__5094\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_7_1_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__8375\,
            in1 => \N__7217\,
            in2 => \_gnd_net_\,
            in3 => \N__7146\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_4_1_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7436\,
            in1 => \N__6073\,
            in2 => \N__5060\,
            in3 => \N__7741\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_366_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__8374\,
            in1 => \N__5204\,
            in2 => \N__5057\,
            in3 => \N__6088\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__7437\,
            in1 => \N__6383\,
            in2 => \N__5054\,
            in3 => \N__5447\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5213\,
            in2 => \N__5207\,
            in3 => \N__9420\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_5_1_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__7435\,
            in1 => \N__7870\,
            in2 => \_gnd_net_\,
            in3 => \N__6364\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5198\,
            in1 => \N__5180\,
            in2 => \_gnd_net_\,
            in3 => \N__9418\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9419\,
            in1 => \N__9644\,
            in2 => \N__5162\,
            in3 => \N__8513\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIEH9V_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__5647\,
            in1 => \N__5620\,
            in2 => \_gnd_net_\,
            in3 => \N__6880\,
            lcout => \U712_CHIP_RAM.N_448\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000100010"
        )
    port map (
            in0 => \N__7286\,
            in1 => \N__7438\,
            in2 => \_gnd_net_\,
            in3 => \N__7126\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_345_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__9645\,
            in1 => \N__7745\,
            in2 => \N__5150\,
            in3 => \N__6087\,
            lcout => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5147\,
            in1 => \N__5132\,
            in2 => \_gnd_net_\,
            in3 => \N__9417\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011011100"
        )
    port map (
            in0 => \N__7151\,
            in1 => \N__6317\,
            in2 => \N__7445\,
            in3 => \N__7294\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011000101"
        )
    port map (
            in0 => \N__5378\,
            in1 => \N__5339\,
            in2 => \N__5372\,
            in3 => \N__5369\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9809\,
            ce => 'H',
            sr => \N__10768\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5354\,
            in2 => \_gnd_net_\,
            in3 => \N__5338\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__8373\,
            in1 => \N__5305\,
            in2 => \N__5294\,
            in3 => \N__5289\,
            lcout => \U712_CYCLE_TERM.N_316_i_0_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001010101010"
        )
    port map (
            in0 => \N__9704\,
            in1 => \N__10328\,
            in2 => \N__10246\,
            in3 => \N__5261\,
            lcout => \U712_BYTE_ENABLE.un1_CUUBEn_i_0_aZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10822\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5273\,
            lcout => \U712_CYCLE_TERM.N_316_i_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101010"
        )
    port map (
            in0 => \N__9705\,
            in1 => \N__10322\,
            in2 => \N__10244\,
            in3 => \N__5257\,
            lcout => \U712_BYTE_ENABLE.un1_CLMBEn_i_0_aZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_x2_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10055\,
            in2 => \_gnd_net_\,
            in3 => \N__10139\,
            lcout => \U712_BYTE_ENABLE.N_282_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5246\,
            in1 => \N__5231\,
            in2 => \_gnd_net_\,
            in3 => \N__9525\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_0_2_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7832\,
            in2 => \_gnd_net_\,
            in3 => \N__7923\,
            lcout => \U712_CHIP_RAM.N_371_1\,
            ltout => \U712_CHIP_RAM.N_371_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__7378\,
            in1 => \N__7193\,
            in2 => \N__5501\,
            in3 => \N__7072\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__5468\,
            in1 => \N__7380\,
            in2 => \_gnd_net_\,
            in3 => \N__5525\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI27TJ3_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__7194\,
            in1 => \N__5474\,
            in2 => \N__6089\,
            in3 => \N__7379\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5462\,
            in3 => \N__7195\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9789\,
            ce => 'H',
            sr => \N__10788\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7813\,
            in1 => \N__7416\,
            in2 => \N__6376\,
            in3 => \N__5448\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9793\,
            ce => \N__5396\,
            sr => \N__10782\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI68LV_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7588\,
            in1 => \N__7069\,
            in2 => \_gnd_net_\,
            in3 => \N__7808\,
            lcout => \U712_CHIP_RAM.N_436\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111000"
        )
    port map (
            in0 => \N__7812\,
            in1 => \N__7415\,
            in2 => \N__7968\,
            in3 => \N__7121\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_i_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101100"
        )
    port map (
            in0 => \N__7414\,
            in1 => \N__7070\,
            in2 => \N__7967\,
            in3 => \N__7811\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_129_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7810\,
            in1 => \N__7285\,
            in2 => \_gnd_net_\,
            in3 => \N__7945\,
            lcout => \U712_CHIP_RAM.N_329\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_2_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__7413\,
            in1 => \N__7809\,
            in2 => \N__7142\,
            in3 => \N__6074\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_414_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110011"
        )
    port map (
            in0 => \N__7546\,
            in1 => \N__7589\,
            in2 => \N__5687\,
            in3 => \N__5563\,
            lcout => \U712_CHIP_RAM.N_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIIPOI5_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000000000"
        )
    port map (
            in0 => \N__5670\,
            in1 => \N__7468\,
            in2 => \N__5624\,
            in3 => \N__5520\,
            lcout => \U712_CHIP_RAM.N_373\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_3_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6356\,
            in1 => \N__7386\,
            in2 => \N__7848\,
            in3 => \N__6068\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER15\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4F6EB_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__6069\,
            in1 => \N__5507\,
            in2 => \N__5537\,
            in3 => \N__5521\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6619\,
            in1 => \N__6634\,
            in2 => \N__6812\,
            in3 => \N__6649\,
            lcout => \U712_CHIP_RAM.N_286\,
            ltout => \U712_CHIP_RAM.N_286_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI16TJ3_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__7209\,
            in1 => \N__7819\,
            in2 => \N__5528\,
            in3 => \N__6355\,
            lcout => \U712_CHIP_RAM.N_486\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_0_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6354\,
            in1 => \N__7385\,
            in2 => \N__7847\,
            in3 => \N__7210\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_2_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7922\,
            in2 => \_gnd_net_\,
            in3 => \N__7071\,
            lcout => \U712_CHIP_RAM.N_287\,
            ltout => \U712_CHIP_RAM.N_287_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIF74S2_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__7815\,
            in1 => \N__7510\,
            in2 => \N__6161\,
            in3 => \N__6158\,
            lcout => \U712_CHIP_RAM.N_283\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__8362\,
            in1 => \N__7007\,
            in2 => \N__6122\,
            in3 => \N__6082\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9801\,
            ce => \N__6017\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__6081\,
            in1 => \N__8363\,
            in2 => \_gnd_net_\,
            in3 => \N__6110\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9801\,
            ce => \N__6017\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__8364\,
            in1 => \N__6305\,
            in2 => \N__6101\,
            in3 => \N__6083\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9801\,
            ce => \N__6017\,
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIAS4F1_0_1_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5993\,
            in1 => \N__5949\,
            in2 => \N__5924\,
            in3 => \N__5873\,
            lcout => \U712_REG_SM.C1_SYNC_RNIAS4F1_0Z0Z_1\,
            ltout => \U712_REG_SM.C1_SYNC_RNIAS4F1_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIOC3L1_4_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5825\,
            in3 => \N__5791\,
            lcout => \U712_REG_SM.ASn_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIKPND1_3_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__7849\,
            in1 => \N__7426\,
            in2 => \_gnd_net_\,
            in3 => \N__8372\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__6563\,
            in1 => \N__5792\,
            in2 => \N__5759\,
            in3 => \N__5712\,
            lcout => \U712_REG_SM.N_104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_6_1_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7521\,
            in2 => \_gnd_net_\,
            in3 => \N__6869\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_RNO_6Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__7965\,
            in1 => \N__8361\,
            in2 => \N__6386\,
            in3 => \N__7144\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__7287\,
            in1 => \N__7850\,
            in2 => \_gnd_net_\,
            in3 => \N__6374\,
            lcout => \U712_CHIP_RAM.N_388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7966\,
            in1 => \N__7218\,
            in2 => \_gnd_net_\,
            in3 => \N__7145\,
            lcout => \U712_CHIP_RAM.N_370\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_38_i_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__8191\,
            in1 => \N__6299\,
            in2 => \N__6228\,
            in3 => \N__7609\,
            lcout => \N_38_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_1_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7612\,
            in1 => \N__8252\,
            in2 => \_gnd_net_\,
            in3 => \N__6224\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_426_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_47_i_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__6605\,
            in1 => \N__6572\,
            in2 => \N__6269\,
            in3 => \N__10327\,
            lcout => \N_47_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7611\,
            in1 => \N__8251\,
            in2 => \_gnd_net_\,
            in3 => \N__6223\,
            lcout => \U712_BYTE_ENABLE.N_431\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_46_i_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000110011"
        )
    port map (
            in0 => \N__8192\,
            in1 => \N__6242\,
            in2 => \N__6229\,
            in3 => \N__7610\,
            lcout => \N_46_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__10061\,
            in1 => \N__10157\,
            in2 => \_gnd_net_\,
            in3 => \N__9706\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2Z0Z_0\,
            ltout => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_45_i_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__6596\,
            in1 => \N__10326\,
            in2 => \N__6590\,
            in3 => \N__6571\,
            lcout => \N_45_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_1_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__9707\,
            in1 => \N__10245\,
            in2 => \_gnd_net_\,
            in3 => \N__10156\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_0_m2_i_m2_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001111111"
        )
    port map (
            in0 => \N__8172\,
            in1 => \N__6555\,
            in2 => \N__8241\,
            in3 => \N__7304\,
            lcout => \N_344\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DMA_LATCH_EN_0_a2_0_a2_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__8171\,
            in1 => \N__8232\,
            in2 => \_gnd_net_\,
            in3 => \N__7303\,
            lcout => \DMA_LATCH_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9703\,
            in1 => \N__6464\,
            in2 => \N__9527\,
            in3 => \N__9335\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__6458\,
            in1 => \N__9522\,
            in2 => \N__9695\,
            in3 => \N__8975\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__8770\,
            in1 => \N__8719\,
            in2 => \N__6449\,
            in3 => \N__9002\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9786\,
            ce => \N__9127\,
            sr => \N__10783\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6425\,
            in1 => \N__6404\,
            in2 => \_gnd_net_\,
            in3 => \N__9521\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__8501\,
            in1 => \N__9523\,
            in2 => \N__6698\,
            in3 => \N__9661\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__8718\,
            in1 => \N__7715\,
            in2 => \N__6695\,
            in3 => \N__8771\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9786\,
            ce => \N__9127\,
            sr => \N__10783\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_cry_c_0_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7114\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7439\,
            in2 => \_gnd_net_\,
            in3 => \N__6659\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6846\,
            in1 => \N__7949\,
            in2 => \_gnd_net_\,
            in3 => \N__6656\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \N__9790\,
            ce => \N__6797\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6843\,
            in1 => \N__7846\,
            in2 => \_gnd_net_\,
            in3 => \N__6653\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__9790\,
            ce => \N__6797\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6847\,
            in1 => \N__6650\,
            in2 => \_gnd_net_\,
            in3 => \N__6638\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__9790\,
            ce => \N__6797\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6844\,
            in1 => \N__6635\,
            in2 => \_gnd_net_\,
            in3 => \N__6623\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__9790\,
            ce => \N__6797\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6848\,
            in1 => \N__6620\,
            in2 => \_gnd_net_\,
            in3 => \N__6608\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__9790\,
            ce => \N__6797\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6845\,
            in1 => \N__6811\,
            in2 => \_gnd_net_\,
            in3 => \N__6815\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9790\,
            ce => \N__6797\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6962\,
            in2 => \_gnd_net_\,
            in3 => \N__6779\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__6733\,
            ce => 'H',
            sr => \N__7457\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7001\,
            in2 => \_gnd_net_\,
            in3 => \N__6776\,
            lcout => \U712_CHIP_RAM.REFRESH5lto1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__6733\,
            ce => 'H',
            sr => \N__7457\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6976\,
            in2 => \_gnd_net_\,
            in3 => \N__6773\,
            lcout => \U712_CHIP_RAM.REFRESH5lto2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__6733\,
            ce => 'H',
            sr => \N__7457\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6925\,
            in2 => \_gnd_net_\,
            in3 => \N__6770\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__6733\,
            ce => 'H',
            sr => \N__7457\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6989\,
            in2 => \_gnd_net_\,
            in3 => \N__6767\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__6733\,
            ce => 'H',
            sr => \N__7457\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6938\,
            in2 => \_gnd_net_\,
            in3 => \N__6764\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__6733\,
            ce => 'H',
            sr => \N__7457\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6950\,
            in2 => \_gnd_net_\,
            in3 => \N__6761\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__6733\,
            ce => 'H',
            sr => \N__7457\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6901\,
            in2 => \_gnd_net_\,
            in3 => \N__6758\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6733\,
            ce => 'H',
            sr => \N__7457\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110001000"
        )
    port map (
            in0 => \N__7706\,
            in1 => \N__8359\,
            in2 => \N__7616\,
            in3 => \N__7512\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIHSHE1_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6870\,
            in1 => \N__8360\,
            in2 => \_gnd_net_\,
            in3 => \N__7511\,
            lcout => \U712_CHIP_RAM.N_201_i_i_a2_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9860\,
            in1 => \N__9933\,
            in2 => \N__8861\,
            in3 => \N__9442\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111011"
        )
    port map (
            in0 => \N__7444\,
            in1 => \N__7284\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_306_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011100000"
        )
    port map (
            in0 => \N__7851\,
            in1 => \N__7220\,
            in2 => \N__7154\,
            in3 => \N__7143\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100111111"
        )
    port map (
            in0 => \N__7000\,
            in1 => \N__6988\,
            in2 => \N__6977\,
            in3 => \N__6961\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6949\,
            in2 => \_gnd_net_\,
            in3 => \N__6937\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111111011"
        )
    port map (
            in0 => \N__6926\,
            in1 => \N__6911\,
            in2 => \N__6905\,
            in3 => \N__6887\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9802\,
            ce => 'H',
            sr => \N__10761\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8190\,
            in2 => \_gnd_net_\,
            in3 => \N__8250\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9806\,
            ce => 'H',
            sr => \N__10758\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7688\,
            in2 => \_gnd_net_\,
            in3 => \N__7696\,
            lcout => \U712_CHIP_RAM.un3_DMA_CYCLE_START\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7697\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9806\,
            ce => 'H',
            sr => \N__10758\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8717\,
            in1 => \N__9065\,
            in2 => \N__8781\,
            in3 => \N__7682\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9783\,
            ce => \N__9128\,
            sr => \N__10778\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__7658\,
            in1 => \N__9498\,
            in2 => \N__9710\,
            in3 => \N__9353\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10823\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7979\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__9494\,
            in1 => \N__9893\,
            in2 => \_gnd_net_\,
            in3 => \N__9963\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => \U712_CHIP_RAM.CMA_5_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__7639\,
            in1 => \N__9657\,
            in2 => \N__7643\,
            in3 => \N__8524\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110001111"
        )
    port map (
            in0 => \N__7640\,
            in1 => \N__9656\,
            in2 => \N__8602\,
            in3 => \N__8525\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNI8NM9_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9524\,
            in3 => \N__9699\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9889\,
            in2 => \_gnd_net_\,
            in3 => \N__9959\,
            lcout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8003\,
            in1 => \N__9689\,
            in2 => \_gnd_net_\,
            in3 => \N__8492\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_463_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111110000"
        )
    port map (
            in0 => \N__9493\,
            in1 => \_gnd_net_\,
            in2 => \N__7982\,
            in3 => \N__8758\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101001111"
        )
    port map (
            in0 => \N__8757\,
            in1 => \N__10520\,
            in2 => \N__9531\,
            in3 => \N__9690\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100001000"
        )
    port map (
            in0 => \N__10519\,
            in1 => \N__9512\,
            in2 => \N__9708\,
            in3 => \N__8759\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100110001"
        )
    port map (
            in0 => \N__9958\,
            in1 => \N__8871\,
            in2 => \N__9895\,
            in3 => \N__9492\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__7921\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7814\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9323\,
            in1 => \N__11062\,
            in2 => \_gnd_net_\,
            in3 => \N__9040\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10888\,
            ce => \N__10857\,
            sr => \N__10766\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11061\,
            in1 => \N__9322\,
            in2 => \_gnd_net_\,
            in3 => \N__9275\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10888\,
            ce => \N__10857\,
            sr => \N__10766\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10466\,
            in1 => \N__9274\,
            in2 => \_gnd_net_\,
            in3 => \N__11059\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            ce => \N__10855\,
            sr => \N__10760\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11060\,
            in1 => \N__9224\,
            in2 => \_gnd_net_\,
            in3 => \N__9039\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            ce => \N__10855\,
            sr => \N__10760\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9026\,
            in1 => \N__11053\,
            in2 => \_gnd_net_\,
            in3 => \N__9321\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__10853\,
            sr => \N__10757\
        );

    \pll_RNI8MQ3_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8474\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8393\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_DRDENn_0_a2_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__8215\,
            in1 => \N__8189\,
            in2 => \_gnd_net_\,
            in3 => \N__8124\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CRCSn_LC_13_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8876\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9782\,
            ce => 'H',
            sr => \N__10803\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_13_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8720\,
            in1 => \N__10403\,
            in2 => \N__8783\,
            in3 => \N__8039\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9784\,
            ce => \N__9130\,
            sr => \N__10789\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8715\,
            in1 => \N__8930\,
            in2 => \N__8782\,
            in3 => \N__8900\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9787\,
            ce => \N__9129\,
            sr => \N__10784\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__9968\,
            in1 => \N__9894\,
            in2 => \N__9526\,
            in3 => \N__8875\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9787\,
            ce => \N__9129\,
            sr => \N__10784\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8822\,
            in1 => \N__8816\,
            in2 => \_gnd_net_\,
            in3 => \N__8810\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9787\,
            ce => \N__9129\,
            sr => \N__10784\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__8766\,
            in1 => \N__8716\,
            in2 => \N__9053\,
            in3 => \N__9359\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9787\,
            ce => \N__9129\,
            sr => \N__10784\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__9673\,
            in1 => \N__8669\,
            in2 => \N__8603\,
            in3 => \N__10901\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9787\,
            ce => \N__9129\,
            sr => \N__10784\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__9179\,
            in1 => \N__9674\,
            in2 => \N__8627\,
            in3 => \N__8601\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9787\,
            ce => \N__9129\,
            sr => \N__10784\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8561\,
            in1 => \N__8540\,
            in2 => \_gnd_net_\,
            in3 => \N__9519\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9520\,
            in1 => \N__9694\,
            in2 => \N__8528\,
            in3 => \N__9341\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9170\,
            in2 => \N__9164\,
            in3 => \N__9161\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9791\,
            ce => \N__9137\,
            sr => \N__10776\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9101\,
            in1 => \N__9083\,
            in2 => \_gnd_net_\,
            in3 => \N__9502\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10613\,
            in1 => \N__11054\,
            in2 => \_gnd_net_\,
            in3 => \N__10505\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10887\,
            ce => \N__10858\,
            sr => \N__10769\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9267\,
            in1 => \N__11055\,
            in2 => \_gnd_net_\,
            in3 => \N__10465\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10887\,
            ce => \N__10858\,
            sr => \N__10769\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__9223\,
            in1 => \_gnd_net_\,
            in2 => \N__11070\,
            in3 => \N__9041\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10887\,
            ce => \N__10858\,
            sr => \N__10769\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8960\,
            in1 => \N__11049\,
            in2 => \_gnd_net_\,
            in3 => \N__10568\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10856\,
            sr => \N__10762\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__11145\,
            in1 => \_gnd_net_\,
            in2 => \N__11069\,
            in3 => \N__9207\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10856\,
            sr => \N__10762\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11016\,
            in1 => \N__10575\,
            in2 => \_gnd_net_\,
            in3 => \N__8956\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10884\,
            ce => \N__10854\,
            sr => \N__10759\
        );

    \U712_CHIP_RAM.CASn_LC_14_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9532\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9785\,
            ce => 'H',
            sr => \N__10804\
        );

    \U712_CHIP_RAM.WEn_LC_14_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9967\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9785\,
            ce => 'H',
            sr => \N__10804\
        );

    \U712_CHIP_RAM.RASn_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9896\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9788\,
            ce => 'H',
            sr => \N__10796\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9709\,
            in1 => \N__9539\,
            in2 => \N__9533\,
            in3 => \N__9230\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11000\,
            in1 => \N__10608\,
            in2 => \_gnd_net_\,
            in3 => \N__10577\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__10860\,
            sr => \N__10777\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10609\,
            in1 => \N__11001\,
            in2 => \_gnd_net_\,
            in3 => \N__10500\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__10860\,
            sr => \N__10777\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10501\,
            in1 => \N__11002\,
            in2 => \_gnd_net_\,
            in3 => \N__10464\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__10860\,
            sr => \N__10777\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9306\,
            in1 => \N__11003\,
            in2 => \_gnd_net_\,
            in3 => \N__9258\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__10860\,
            sr => \N__10777\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9216\,
            in1 => \N__11012\,
            in2 => \_gnd_net_\,
            in3 => \N__11152\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10885\,
            ce => \N__10859\,
            sr => \N__10771\
        );

    \U712_BYTE_ENABLE.N_357_i_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011100000"
        )
    port map (
            in0 => \N__10276\,
            in1 => \N__10236\,
            in2 => \N__10155\,
            in3 => \N__10035\,
            lcout => \N_357_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_UDSn_i_0_0_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__10241\,
            in1 => \N__10376\,
            in2 => \_gnd_net_\,
            in3 => \N__10122\,
            lcout => \N_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UMBE_i_o2_i_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111000000"
        )
    port map (
            in0 => \N__10240\,
            in1 => \N__10306\,
            in2 => \N__10048\,
            in3 => \N__10121\,
            lcout => \N_231\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10996\,
            in1 => \N__10607\,
            in2 => \_gnd_net_\,
            in3 => \N__10576\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10886\,
            ce => \N__10861\,
            sr => \N__10785\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__10499\,
            in1 => \_gnd_net_\,
            in2 => \N__11032\,
            in3 => \N__10454\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10886\,
            ce => \N__10861\,
            sr => \N__10785\
        );

    \U712_BYTE_ENABLE.N_358_i_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000111000100"
        )
    port map (
            in0 => \N__10291\,
            in1 => \N__10060\,
            in2 => \N__10247\,
            in3 => \N__10147\,
            lcout => \N_358_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011111111"
        )
    port map (
            in0 => \N__10143\,
            in1 => \N__10243\,
            in2 => \_gnd_net_\,
            in3 => \N__10375\,
            lcout => \N_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_0_0_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101110000"
        )
    port map (
            in0 => \N__10307\,
            in1 => \N__10242\,
            in2 => \N__10154\,
            in3 => \N__10059\,
            lcout => \LLBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_22_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__11127\,
            in1 => \N__11084\,
            in2 => \_gnd_net_\,
            in3 => \N__11048\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10883\,
            ce => \N__10862\,
            sr => \N__10807\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     May 6 2025 20:26:24

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DA : out std_logic_vector(2 downto 0);
    A : in std_logic_vector(20 downto 0);
    DBRn : in std_logic;
    RAMENn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    TCIn : out std_logic;
    TBIn : out std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__12772\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7827\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_555_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_390_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_2_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_2_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_2_2\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.m77_0_a2_0_2_cascade_\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \A_c_8\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_3\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_7\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.N_436_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_194_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_20_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER41_0_a3_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.m101_i_1\ : std_logic;
signal \U712_CHIP_RAM.N_305_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_376\ : std_logic;
signal \U712_CHIP_RAM.m101_i_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.m101_i_2\ : std_logic;
signal \U712_CHIP_RAM.N_304_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_312_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.N_39\ : std_logic;
signal \U712_CHIP_RAM.N_326\ : std_logic;
signal \U712_CHIP_RAM.N_39_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.N_307_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_467_cascade_\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_440\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_1\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.un3_DBR_COUNT_cry_1\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.un3_DBR_COUNT_cry_2\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.un3_DBR_COUNT_cry_3\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.un3_DBR_COUNT_cry_4\ : std_logic;
signal \U712_CHIP_RAM.un3_DBR_COUNT_cry_5\ : std_logic;
signal \U712_CHIP_RAM.un3_DBR_COUNT_cry_6\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_7\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_6\ : std_logic;
signal \U712_CHIP_RAM.N_194\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_5_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_378\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDs_0_4\ : std_logic;
signal \U712_CHIP_RAM.N_396_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_0_2\ : std_logic;
signal \U712_CHIP_RAM.N_397\ : std_logic;
signal \U712_CHIP_RAM.N_555\ : std_logic;
signal \U712_CHIP_RAM.N_449\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDs_0_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_1_3\ : std_logic;
signal \U712_CHIP_RAM.N_194_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_i_0_9\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.m123_i_2\ : std_logic;
signal \U712_CHIP_RAM.N_305\ : std_logic;
signal \U712_CHIP_RAM.N_190\ : std_logic;
signal \U712_CHIP_RAM.N_476\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_344\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_307\ : std_logic;
signal \U712_CHIP_RAM.N_551_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_304\ : std_logic;
signal \U712_CHIP_RAM.N_435_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_325\ : std_logic;
signal \U712_CHIP_RAM.N_321\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_551\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER41_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.LATCH_CLK_6\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.m93_i_a2_5\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.m93_i_a2_4\ : std_logic;
signal \U712_CHIP_RAM.N_428_cascade_\ : std_logic;
signal \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_430\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto7_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lt7\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_335_cascade_\ : std_logic;
signal \N_202_i\ : std_logic;
signal \TSn_c\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \N_165_i\ : std_logic;
signal \WEn_c\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA25_0_i_cascade_\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_361\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \A_c_13\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_435\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0\ : std_logic;
signal \U712_CHIP_RAM.N_467\ : std_logic;
signal \U712_CHIP_RAM.DBENn_7_0_0\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.N_367\ : std_logic;
signal \U712_CHIP_RAM.N_419\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_10_10_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \U712_REG_SM.N_402\ : std_logic;
signal \U712_REG_SM.START_RSTZ0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0\ : std_logic;
signal \U712_CHIP_RAM.N_314\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA25_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_REG_SM.N_373_cascade_\ : std_logic;
signal \U712_REG_SM.N_130\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ1Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\ : std_logic;
signal \U712_REG_SM.N_406\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_328_cascade_\ : std_logic;
signal \U712_REG_SM.N_331_cascade_\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\ : std_logic;
signal \U712_REG_SM.N_328\ : std_logic;
signal \U712_REG_SM.N_412\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.REGENn_e_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_0\ : std_logic;
signal \REGENn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.N_332\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.N_455_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \U712_REG_SM.N_373\ : std_logic;
signal \U712_REG_SM.N_330_cascade_\ : std_logic;
signal \U712_REG_SM.N_413\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_410\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_2\ : std_logic;
signal \U712_REG_SM.STATE_COUNTc_0_0\ : std_logic;
signal \U712_REG_SM.N_308\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.N_308_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_1\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_2\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0\ : std_logic;
signal \N_336_i\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_1\ : std_logic;
signal \LDSn_c\ : std_logic;
signal \U712_REG_SM.N_459\ : std_logic;
signal \U712_REG_SM.un1_REGENn_0_sqmuxa_0\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \UDSn_c\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \U712_REG_SM.N_404\ : std_logic;
signal \N_335_i\ : std_logic;
signal \N_337_i\ : std_logic;
signal \N_177_i\ : std_logic;
signal \N_334\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0\ : std_logic;
signal \N_175_i\ : std_logic;
signal \N_336\ : std_logic;
signal \U712_CHIP_RAM.m50_i_a2_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_337_cascade_\ : std_logic;
signal \N_200_i\ : std_logic;
signal \A_c_1\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \N_334_i\ : std_logic;
signal \RnW_c\ : std_logic;
signal \DMA_WRITE_CYCLE\ : std_logic;
signal \N_379\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \N_167_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \DA_wire\ : std_logic_vector(2 downto 0);
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    TBIn <= \TBIn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    ASn <= \ASn_wire\;
    DA <= \DA_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    TCIn <= \TCIn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__4344\,
            RESETB => \N__7365\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12772\,
            DIN => \N__12771\,
            DOUT => \N__12770\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12772\,
            PADOUT => \N__12771\,
            PADIN => \N__12770\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7422\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12763\,
            DIN => \N__12762\,
            DOUT => \N__12761\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12763\,
            PADOUT => \N__12762\,
            PADIN => \N__12761\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12754\,
            DIN => \N__12753\,
            DOUT => \N__12752\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12754\,
            PADOUT => \N__12753\,
            PADIN => \N__12752\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8226\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12745\,
            DIN => \N__12744\,
            DOUT => \N__12743\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12745\,
            PADOUT => \N__12744\,
            PADIN => \N__12743\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11142\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12736\,
            DIN => \N__12735\,
            DOUT => \N__12734\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12736\,
            PADOUT => \N__12735\,
            PADIN => \N__12734\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12727\,
            DIN => \N__12726\,
            DOUT => \N__12725\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12727\,
            PADOUT => \N__12726\,
            PADIN => \N__12725\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12718\,
            DIN => \N__12717\,
            DOUT => \N__12716\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12718\,
            PADOUT => \N__12717\,
            PADIN => \N__12716\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12709\,
            DIN => \N__12708\,
            DOUT => \N__12707\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12709\,
            PADOUT => \N__12708\,
            PADIN => \N__12707\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12700\,
            DIN => \N__12699\,
            DOUT => \N__12698\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12700\,
            PADOUT => \N__12699\,
            PADIN => \N__12698\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12691\,
            DIN => \N__12690\,
            DOUT => \N__12689\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12691\,
            PADOUT => \N__12690\,
            PADIN => \N__12689\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12682\,
            DIN => \N__12681\,
            DOUT => \N__12680\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12682\,
            PADOUT => \N__12681\,
            PADIN => \N__12680\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12673\,
            DIN => \N__12672\,
            DOUT => \N__12671\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12673\,
            PADOUT => \N__12672\,
            PADIN => \N__12671\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7671\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12664\,
            DIN => \N__12663\,
            DOUT => \N__12662\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12664\,
            PADOUT => \N__12663\,
            PADIN => \N__12662\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9408\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12655\,
            DIN => \N__12654\,
            DOUT => \N__12653\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12655\,
            PADOUT => \N__12654\,
            PADIN => \N__12653\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12646\,
            DIN => \N__12645\,
            DOUT => \N__12644\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12646\,
            PADOUT => \N__12645\,
            PADIN => \N__12644\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5910\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12637\,
            DIN => \N__12636\,
            DOUT => \N__12635\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12637\,
            PADOUT => \N__12636\,
            PADIN => \N__12635\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12628\,
            DIN => \N__12627\,
            DOUT => \N__12626\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12628\,
            PADOUT => \N__12627\,
            PADIN => \N__12626\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12619\,
            DIN => \N__12618\,
            DOUT => \N__12617\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12619\,
            PADOUT => \N__12618\,
            PADIN => \N__12617\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4956\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12610\,
            DIN => \N__12609\,
            DOUT => \N__12608\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12610\,
            PADOUT => \N__12609\,
            PADIN => \N__12608\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12601\,
            DIN => \N__12600\,
            DOUT => \N__12599\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12601\,
            PADOUT => \N__12600\,
            PADIN => \N__12599\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12592\,
            DIN => \N__12591\,
            DOUT => \N__12590\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12592\,
            PADOUT => \N__12591\,
            PADIN => \N__12590\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7308\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12583\,
            DIN => \N__12582\,
            DOUT => \N__12581\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12583\,
            PADOUT => \N__12582\,
            PADIN => \N__12581\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12574\,
            DIN => \N__12573\,
            DOUT => \N__12572\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12574\,
            PADOUT => \N__12573\,
            PADIN => \N__12572\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7335\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12565\,
            DIN => \N__12564\,
            DOUT => \N__12563\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12565\,
            PADOUT => \N__12564\,
            PADIN => \N__12563\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12556\,
            DIN => \N__12555\,
            DOUT => \N__12554\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12556\,
            PADOUT => \N__12555\,
            PADIN => \N__12554\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9630\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12547\,
            DIN => \N__12546\,
            DOUT => \N__12545\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12547\,
            PADOUT => \N__12546\,
            PADIN => \N__12545\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8045\,
            DIN0 => OPEN,
            DOUT0 => \N__7289\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12538\,
            DIN => \N__12537\,
            DOUT => \N__12536\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12538\,
            PADOUT => \N__12537\,
            PADIN => \N__12536\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12529\,
            DIN => \N__12528\,
            DOUT => \N__12527\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12529\,
            PADOUT => \N__12528\,
            PADIN => \N__12527\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12520\,
            DIN => \N__12519\,
            DOUT => \N__12518\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12520\,
            PADOUT => \N__12519\,
            PADIN => \N__12518\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12511\,
            DIN => \N__12510\,
            DOUT => \N__12509\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12511\,
            PADOUT => \N__12510\,
            PADIN => \N__12509\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12502\,
            DIN => \N__12501\,
            DOUT => \N__12500\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12502\,
            PADOUT => \N__12501\,
            PADIN => \N__12500\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12493\,
            DIN => \N__12492\,
            DOUT => \N__12491\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12493\,
            PADOUT => \N__12492\,
            PADIN => \N__12491\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6441\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12484\,
            DIN => \N__12483\,
            DOUT => \N__12482\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12484\,
            PADOUT => \N__12483\,
            PADIN => \N__12482\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12475\,
            DIN => \N__12474\,
            DOUT => \N__12473\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12475\,
            PADOUT => \N__12474\,
            PADIN => \N__12473\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12466\,
            DIN => \N__12465\,
            DOUT => \N__12464\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12466\,
            PADOUT => \N__12465\,
            PADIN => \N__12464\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12457\,
            DIN => \N__12456\,
            DOUT => \N__12455\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12457\,
            PADOUT => \N__12456\,
            PADIN => \N__12455\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12448\,
            DIN => \N__12447\,
            DOUT => \N__12446\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12448\,
            PADOUT => \N__12447\,
            PADIN => \N__12446\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12439\,
            DIN => \N__12438\,
            DOUT => \N__12437\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12439\,
            PADOUT => \N__12438\,
            PADIN => \N__12437\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6399\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12430\,
            DIN => \N__12429\,
            DOUT => \N__12428\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12430\,
            PADOUT => \N__12429\,
            PADIN => \N__12428\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12421\,
            DIN => \N__12420\,
            DOUT => \N__12419\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12421\,
            PADOUT => \N__12420\,
            PADIN => \N__12419\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12412\,
            DIN => \N__12411\,
            DOUT => \N__12410\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12412\,
            PADOUT => \N__12411\,
            PADIN => \N__12410\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9435\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12403\,
            DIN => \N__12402\,
            DOUT => \N__12401\,
            PACKAGEPIN => \DA_wire\(0)
        );

    \DA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12403\,
            PADOUT => \N__12402\,
            PADIN => \N__12401\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6563\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12394\,
            DIN => \N__12393\,
            DOUT => \N__12392\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12394\,
            PADOUT => \N__12393\,
            PADIN => \N__12392\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12385\,
            DIN => \N__12384\,
            DOUT => \N__12383\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12385\,
            PADOUT => \N__12384\,
            PADIN => \N__12383\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7878\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12376\,
            DIN => \N__12375\,
            DOUT => \N__12374\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12376\,
            PADOUT => \N__12375\,
            PADIN => \N__12374\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7821\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12367\,
            DIN => \N__12366\,
            DOUT => \N__12365\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12367\,
            PADOUT => \N__12366\,
            PADIN => \N__12365\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8403\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12358\,
            DIN => \N__12357\,
            DOUT => \N__12356\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12358\,
            PADOUT => \N__12357\,
            PADIN => \N__12356\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12349\,
            DIN => \N__12348\,
            DOUT => \N__12347\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12349\,
            PADOUT => \N__12348\,
            PADIN => \N__12347\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12340\,
            DIN => \N__12339\,
            DOUT => \N__12338\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12340\,
            PADOUT => \N__12339\,
            PADIN => \N__12338\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11727\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12331\,
            DIN => \N__12330\,
            DOUT => \N__12329\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12331\,
            PADOUT => \N__12330\,
            PADIN => \N__12329\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8049\,
            DIN0 => OPEN,
            DOUT0 => \N__7290\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12322\,
            DIN => \N__12321\,
            DOUT => \N__12320\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12322\,
            PADOUT => \N__12321\,
            PADIN => \N__12320\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6423\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12313\,
            DIN => \N__12312\,
            DOUT => \N__12311\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12313\,
            PADOUT => \N__12312\,
            PADIN => \N__12311\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6867\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12304\,
            DIN => \N__12303\,
            DOUT => \N__12302\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12304\,
            PADOUT => \N__12303\,
            PADIN => \N__12302\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11844\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12295\,
            DIN => \N__12294\,
            DOUT => \N__12293\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12295\,
            PADOUT => \N__12294\,
            PADIN => \N__12293\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12286\,
            DIN => \N__12285\,
            DOUT => \N__12284\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12286\,
            PADOUT => \N__12285\,
            PADIN => \N__12284\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12277\,
            DIN => \N__12276\,
            DOUT => \N__12275\,
            PACKAGEPIN => \DA_wire\(2)
        );

    \DA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12277\,
            PADOUT => \N__12276\,
            PADIN => \N__12275\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5805\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12268\,
            DIN => \N__12267\,
            DOUT => \N__12266\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12268\,
            PADOUT => \N__12267\,
            PADIN => \N__12266\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12259\,
            DIN => \N__12258\,
            DOUT => \N__12257\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12259\,
            PADOUT => \N__12258\,
            PADIN => \N__12257\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12250\,
            DIN => \N__12249\,
            DOUT => \N__12248\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12250\,
            PADOUT => \N__12249\,
            PADIN => \N__12248\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6747\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12241\,
            DIN => \N__12240\,
            DOUT => \N__12239\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12241\,
            PADOUT => \N__12240\,
            PADIN => \N__12239\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9615\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12232\,
            DIN => \N__12231\,
            DOUT => \N__12230\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12232\,
            PADOUT => \N__12231\,
            PADIN => \N__12230\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12223\,
            DIN => \N__12222\,
            DOUT => \N__12221\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12223\,
            PADOUT => \N__12222\,
            PADIN => \N__12221\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11787\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12214\,
            DIN => \N__12213\,
            DOUT => \N__12212\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12214\,
            PADOUT => \N__12213\,
            PADIN => \N__12212\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8035\,
            DIN0 => OPEN,
            DOUT0 => \N__7285\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12205\,
            DIN => \N__12204\,
            DOUT => \N__12203\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12205\,
            PADOUT => \N__12204\,
            PADIN => \N__12203\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7842\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12196\,
            DIN => \N__12195\,
            DOUT => \N__12194\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12196\,
            PADOUT => \N__12195\,
            PADIN => \N__12194\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12187\,
            DIN => \N__12186\,
            DOUT => \N__12185\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12187\,
            PADOUT => \N__12186\,
            PADIN => \N__12185\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12178\,
            DIN => \N__12177\,
            DOUT => \N__12176\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12178\,
            PADOUT => \N__12177\,
            PADIN => \N__12176\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5700\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12169\,
            DIN => \N__12168\,
            DOUT => \N__12167\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12169\,
            PADOUT => \N__12168\,
            PADIN => \N__12167\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12160\,
            DIN => \N__12159\,
            DOUT => \N__12158\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12160\,
            PADOUT => \N__12159\,
            PADIN => \N__12158\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12151\,
            DIN => \N__12150\,
            DOUT => \N__12149\,
            PACKAGEPIN => \DA_wire\(1)
        );

    \DA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12151\,
            PADOUT => \N__12150\,
            PADIN => \N__12149\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6813\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12142\,
            DIN => \N__12141\,
            DOUT => \N__12140\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12142\,
            PADOUT => \N__12141\,
            PADIN => \N__12140\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12133\,
            DIN => \N__12132\,
            DOUT => \N__12131\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12133\,
            PADOUT => \N__12132\,
            PADIN => \N__12131\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12124\,
            DIN => \N__12123\,
            DOUT => \N__12122\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12124\,
            PADOUT => \N__12123\,
            PADIN => \N__12122\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6837\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12115\,
            DIN => \N__12114\,
            DOUT => \N__12113\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12115\,
            PADOUT => \N__12114\,
            PADIN => \N__12113\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10023\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12106\,
            DIN => \N__12105\,
            DOUT => \N__12104\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12106\,
            PADOUT => \N__12105\,
            PADIN => \N__12104\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11274\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12097\,
            DIN => \N__12096\,
            DOUT => \N__12095\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12097\,
            PADOUT => \N__12096\,
            PADIN => \N__12095\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4446\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12088\,
            DIN => \N__12087\,
            DOUT => \N__12086\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12088\,
            PADOUT => \N__12087\,
            PADIN => \N__12086\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12079\,
            DIN => \N__12078\,
            DOUT => \N__12077\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12079\,
            PADOUT => \N__12078\,
            PADIN => \N__12077\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12070\,
            DIN => \N__12069\,
            DOUT => \N__12068\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12070\,
            PADOUT => \N__12069\,
            PADIN => \N__12068\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5028\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12061\,
            DIN => \N__12060\,
            DOUT => \N__12059\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12061\,
            PADOUT => \N__12060\,
            PADIN => \N__12059\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12052\,
            DIN => \N__12051\,
            DOUT => \N__12050\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12052\,
            PADOUT => \N__12051\,
            PADIN => \N__12050\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12043\,
            DIN => \N__12042\,
            DOUT => \N__12041\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12043\,
            PADOUT => \N__12042\,
            PADIN => \N__12041\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5909\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12034\,
            DIN => \N__12033\,
            DOUT => \N__12032\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12034\,
            PADOUT => \N__12033\,
            PADIN => \N__12032\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10170\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12025\,
            DIN => \N__12024\,
            DOUT => \N__12023\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12025\,
            PADOUT => \N__12024\,
            PADIN => \N__12023\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8520\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12016\,
            DIN => \N__12015\,
            DOUT => \N__12014\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12016\,
            PADOUT => \N__12015\,
            PADIN => \N__12014\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12007\,
            DIN => \N__12006\,
            DOUT => \N__12005\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12007\,
            PADOUT => \N__12006\,
            PADIN => \N__12005\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8513\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11998\,
            DIN => \N__11997\,
            DOUT => \N__11996\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11998\,
            PADOUT => \N__11997\,
            PADIN => \N__11996\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4404\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11989\,
            DIN => \N__11988\,
            DOUT => \N__11987\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11989\,
            PADOUT => \N__11988\,
            PADIN => \N__11987\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6669\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11980\,
            DIN => \N__11979\,
            DOUT => \N__11978\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11980\,
            PADOUT => \N__11979\,
            PADIN => \N__11978\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11971\,
            DIN => \N__11970\,
            DOUT => \N__11969\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11971\,
            PADOUT => \N__11970\,
            PADIN => \N__11969\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11962\,
            DIN => \N__11961\,
            DOUT => \N__11960\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11962\,
            PADOUT => \N__11961\,
            PADIN => \N__11960\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11953\,
            DIN => \N__11952\,
            DOUT => \N__11951\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11953\,
            PADOUT => \N__11952\,
            PADIN => \N__11951\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11944\,
            DIN => \N__11943\,
            DOUT => \N__11942\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11944\,
            PADOUT => \N__11943\,
            PADIN => \N__11942\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8498\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11935\,
            DIN => \N__11934\,
            DOUT => \N__11933\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11935\,
            PADOUT => \N__11934\,
            PADIN => \N__11933\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11859\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11926\,
            DIN => \N__11925\,
            DOUT => \N__11924\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11926\,
            PADOUT => \N__11925\,
            PADIN => \N__11924\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6501\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11917\,
            DIN => \N__11916\,
            DOUT => \N__11915\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11917\,
            PADOUT => \N__11916\,
            PADIN => \N__11915\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5655\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2899\ : InMux
    port map (
            O => \N__11898\,
            I => \N__11894\
        );

    \I__2898\ : InMux
    port map (
            O => \N__11897\,
            I => \N__11891\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__11894\,
            I => \N__11888\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__11891\,
            I => \N__11885\
        );

    \I__2895\ : Span12Mux_v
    port map (
            O => \N__11888\,
            I => \N__11881\
        );

    \I__2894\ : Span4Mux_v
    port map (
            O => \N__11885\,
            I => \N__11878\
        );

    \I__2893\ : CascadeMux
    port map (
            O => \N__11884\,
            I => \N__11875\
        );

    \I__2892\ : Span12Mux_h
    port map (
            O => \N__11881\,
            I => \N__11872\
        );

    \I__2891\ : Span4Mux_v
    port map (
            O => \N__11878\,
            I => \N__11869\
        );

    \I__2890\ : InMux
    port map (
            O => \N__11875\,
            I => \N__11866\
        );

    \I__2889\ : Odrv12
    port map (
            O => \N__11872\,
            I => \REG_CYCLEm\
        );

    \I__2888\ : Odrv4
    port map (
            O => \N__11869\,
            I => \REG_CYCLEm\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__11866\,
            I => \REG_CYCLEm\
        );

    \I__2886\ : IoInMux
    port map (
            O => \N__11859\,
            I => \N__11856\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__11856\,
            I => \N__11853\
        );

    \I__2884\ : Span4Mux_s3_v
    port map (
            O => \N__11853\,
            I => \N__11850\
        );

    \I__2883\ : Span4Mux_v
    port map (
            O => \N__11850\,
            I => \N__11847\
        );

    \I__2882\ : Odrv4
    port map (
            O => \N__11847\,
            I => \N_167_i\
        );

    \I__2881\ : IoInMux
    port map (
            O => \N__11844\,
            I => \N__11841\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__11841\,
            I => \N__11838\
        );

    \I__2879\ : Span4Mux_s3_h
    port map (
            O => \N__11838\,
            I => \N__11835\
        );

    \I__2878\ : Span4Mux_h
    port map (
            O => \N__11835\,
            I => \N__11832\
        );

    \I__2877\ : Span4Mux_h
    port map (
            O => \N__11832\,
            I => \N__11829\
        );

    \I__2876\ : Sp12to4
    port map (
            O => \N__11829\,
            I => \N__11826\
        );

    \I__2875\ : Span12Mux_v
    port map (
            O => \N__11826\,
            I => \N__11823\
        );

    \I__2874\ : Odrv12
    port map (
            O => \N__11823\,
            I => \N_177_i\
        );

    \I__2873\ : CascadeMux
    port map (
            O => \N__11820\,
            I => \N__11817\
        );

    \I__2872\ : InMux
    port map (
            O => \N__11817\,
            I => \N__11814\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__11814\,
            I => \N__11811\
        );

    \I__2870\ : Odrv4
    port map (
            O => \N__11811\,
            I => \N_334\
        );

    \I__2869\ : InMux
    port map (
            O => \N__11808\,
            I => \N__11805\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__11805\,
            I => \N__11801\
        );

    \I__2867\ : InMux
    port map (
            O => \N__11804\,
            I => \N__11798\
        );

    \I__2866\ : Span4Mux_h
    port map (
            O => \N__11801\,
            I => \N__11793\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__11798\,
            I => \N__11793\
        );

    \I__2864\ : Span4Mux_h
    port map (
            O => \N__11793\,
            I => \N__11790\
        );

    \I__2863\ : Odrv4
    port map (
            O => \N__11790\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0\
        );

    \I__2862\ : IoInMux
    port map (
            O => \N__11787\,
            I => \N__11784\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__11784\,
            I => \N__11781\
        );

    \I__2860\ : IoSpan4Mux
    port map (
            O => \N__11781\,
            I => \N__11778\
        );

    \I__2859\ : Span4Mux_s3_h
    port map (
            O => \N__11778\,
            I => \N__11775\
        );

    \I__2858\ : Span4Mux_v
    port map (
            O => \N__11775\,
            I => \N__11772\
        );

    \I__2857\ : Span4Mux_h
    port map (
            O => \N__11772\,
            I => \N__11769\
        );

    \I__2856\ : Odrv4
    port map (
            O => \N__11769\,
            I => \N_175_i\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__11766\,
            I => \N__11763\
        );

    \I__2854\ : InMux
    port map (
            O => \N__11763\,
            I => \N__11760\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__11760\,
            I => \N__11757\
        );

    \I__2852\ : Odrv4
    port map (
            O => \N__11757\,
            I => \N_336\
        );

    \I__2851\ : InMux
    port map (
            O => \N__11754\,
            I => \N__11751\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__11751\,
            I => \N__11748\
        );

    \I__2849\ : Span4Mux_v
    port map (
            O => \N__11748\,
            I => \N__11744\
        );

    \I__2848\ : InMux
    port map (
            O => \N__11747\,
            I => \N__11741\
        );

    \I__2847\ : Sp12to4
    port map (
            O => \N__11744\,
            I => \N__11738\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__11741\,
            I => \N__11735\
        );

    \I__2845\ : Odrv12
    port map (
            O => \N__11738\,
            I => \U712_CHIP_RAM.m50_i_a2_0_0\
        );

    \I__2844\ : Odrv4
    port map (
            O => \N__11735\,
            I => \U712_CHIP_RAM.m50_i_a2_0_0\
        );

    \I__2843\ : CascadeMux
    port map (
            O => \N__11730\,
            I => \U712_CHIP_RAM.N_337_cascade_\
        );

    \I__2842\ : IoInMux
    port map (
            O => \N__11727\,
            I => \N__11724\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__11724\,
            I => \N__11721\
        );

    \I__2840\ : IoSpan4Mux
    port map (
            O => \N__11721\,
            I => \N__11718\
        );

    \I__2839\ : Sp12to4
    port map (
            O => \N__11718\,
            I => \N__11715\
        );

    \I__2838\ : Span12Mux_s7_v
    port map (
            O => \N__11715\,
            I => \N__11712\
        );

    \I__2837\ : Span12Mux_v
    port map (
            O => \N__11712\,
            I => \N__11709\
        );

    \I__2836\ : Odrv12
    port map (
            O => \N__11709\,
            I => \N_200_i\
        );

    \I__2835\ : CascadeMux
    port map (
            O => \N__11706\,
            I => \N__11702\
        );

    \I__2834\ : InMux
    port map (
            O => \N__11705\,
            I => \N__11698\
        );

    \I__2833\ : InMux
    port map (
            O => \N__11702\,
            I => \N__11693\
        );

    \I__2832\ : InMux
    port map (
            O => \N__11701\,
            I => \N__11693\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__11698\,
            I => \N__11685\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__11693\,
            I => \N__11682\
        );

    \I__2829\ : InMux
    port map (
            O => \N__11692\,
            I => \N__11679\
        );

    \I__2828\ : InMux
    port map (
            O => \N__11691\,
            I => \N__11674\
        );

    \I__2827\ : InMux
    port map (
            O => \N__11690\,
            I => \N__11674\
        );

    \I__2826\ : InMux
    port map (
            O => \N__11689\,
            I => \N__11671\
        );

    \I__2825\ : InMux
    port map (
            O => \N__11688\,
            I => \N__11668\
        );

    \I__2824\ : Span4Mux_v
    port map (
            O => \N__11685\,
            I => \N__11665\
        );

    \I__2823\ : Span4Mux_v
    port map (
            O => \N__11682\,
            I => \N__11662\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__11679\,
            I => \N__11659\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__11674\,
            I => \N__11654\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__11671\,
            I => \N__11654\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__11668\,
            I => \N__11651\
        );

    \I__2818\ : Span4Mux_v
    port map (
            O => \N__11665\,
            I => \N__11648\
        );

    \I__2817\ : Span4Mux_v
    port map (
            O => \N__11662\,
            I => \N__11643\
        );

    \I__2816\ : Span4Mux_v
    port map (
            O => \N__11659\,
            I => \N__11643\
        );

    \I__2815\ : Span4Mux_v
    port map (
            O => \N__11654\,
            I => \N__11640\
        );

    \I__2814\ : Span4Mux_v
    port map (
            O => \N__11651\,
            I => \N__11637\
        );

    \I__2813\ : Sp12to4
    port map (
            O => \N__11648\,
            I => \N__11630\
        );

    \I__2812\ : Sp12to4
    port map (
            O => \N__11643\,
            I => \N__11630\
        );

    \I__2811\ : Sp12to4
    port map (
            O => \N__11640\,
            I => \N__11630\
        );

    \I__2810\ : Span4Mux_v
    port map (
            O => \N__11637\,
            I => \N__11627\
        );

    \I__2809\ : Span12Mux_h
    port map (
            O => \N__11630\,
            I => \N__11622\
        );

    \I__2808\ : Sp12to4
    port map (
            O => \N__11627\,
            I => \N__11622\
        );

    \I__2807\ : Odrv12
    port map (
            O => \N__11622\,
            I => \A_c_1\
        );

    \I__2806\ : CascadeMux
    port map (
            O => \N__11619\,
            I => \N__11613\
        );

    \I__2805\ : InMux
    port map (
            O => \N__11618\,
            I => \N__11609\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__11617\,
            I => \N__11604\
        );

    \I__2803\ : InMux
    port map (
            O => \N__11616\,
            I => \N__11598\
        );

    \I__2802\ : InMux
    port map (
            O => \N__11613\,
            I => \N__11595\
        );

    \I__2801\ : InMux
    port map (
            O => \N__11612\,
            I => \N__11592\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__11609\,
            I => \N__11589\
        );

    \I__2799\ : InMux
    port map (
            O => \N__11608\,
            I => \N__11584\
        );

    \I__2798\ : InMux
    port map (
            O => \N__11607\,
            I => \N__11584\
        );

    \I__2797\ : InMux
    port map (
            O => \N__11604\,
            I => \N__11581\
        );

    \I__2796\ : InMux
    port map (
            O => \N__11603\,
            I => \N__11578\
        );

    \I__2795\ : InMux
    port map (
            O => \N__11602\,
            I => \N__11575\
        );

    \I__2794\ : CascadeMux
    port map (
            O => \N__11601\,
            I => \N__11572\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__11598\,
            I => \N__11567\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__11595\,
            I => \N__11567\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__11592\,
            I => \N__11564\
        );

    \I__2790\ : Span4Mux_h
    port map (
            O => \N__11589\,
            I => \N__11557\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__11584\,
            I => \N__11557\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__11581\,
            I => \N__11557\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__11578\,
            I => \N__11552\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__11575\,
            I => \N__11552\
        );

    \I__2785\ : InMux
    port map (
            O => \N__11572\,
            I => \N__11549\
        );

    \I__2784\ : Span4Mux_v
    port map (
            O => \N__11567\,
            I => \N__11546\
        );

    \I__2783\ : Span4Mux_v
    port map (
            O => \N__11564\,
            I => \N__11543\
        );

    \I__2782\ : Span4Mux_v
    port map (
            O => \N__11557\,
            I => \N__11538\
        );

    \I__2781\ : Span4Mux_v
    port map (
            O => \N__11552\,
            I => \N__11538\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__11549\,
            I => \N__11535\
        );

    \I__2779\ : Sp12to4
    port map (
            O => \N__11546\,
            I => \N__11528\
        );

    \I__2778\ : Sp12to4
    port map (
            O => \N__11543\,
            I => \N__11528\
        );

    \I__2777\ : Sp12to4
    port map (
            O => \N__11538\,
            I => \N__11528\
        );

    \I__2776\ : Span4Mux_v
    port map (
            O => \N__11535\,
            I => \N__11525\
        );

    \I__2775\ : Span12Mux_h
    port map (
            O => \N__11528\,
            I => \N__11520\
        );

    \I__2774\ : Sp12to4
    port map (
            O => \N__11525\,
            I => \N__11520\
        );

    \I__2773\ : Odrv12
    port map (
            O => \N__11520\,
            I => \A_c_0\
        );

    \I__2772\ : InMux
    port map (
            O => \N__11517\,
            I => \N__11512\
        );

    \I__2771\ : CascadeMux
    port map (
            O => \N__11516\,
            I => \N__11509\
        );

    \I__2770\ : InMux
    port map (
            O => \N__11515\,
            I => \N__11506\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__11512\,
            I => \N__11503\
        );

    \I__2768\ : InMux
    port map (
            O => \N__11509\,
            I => \N__11500\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__11506\,
            I => \N__11494\
        );

    \I__2766\ : Span4Mux_v
    port map (
            O => \N__11503\,
            I => \N__11491\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__11500\,
            I => \N__11488\
        );

    \I__2764\ : InMux
    port map (
            O => \N__11499\,
            I => \N__11483\
        );

    \I__2763\ : InMux
    port map (
            O => \N__11498\,
            I => \N__11483\
        );

    \I__2762\ : InMux
    port map (
            O => \N__11497\,
            I => \N__11478\
        );

    \I__2761\ : Span4Mux_v
    port map (
            O => \N__11494\,
            I => \N__11475\
        );

    \I__2760\ : Span4Mux_v
    port map (
            O => \N__11491\,
            I => \N__11468\
        );

    \I__2759\ : Span4Mux_h
    port map (
            O => \N__11488\,
            I => \N__11468\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__11483\,
            I => \N__11468\
        );

    \I__2757\ : InMux
    port map (
            O => \N__11482\,
            I => \N__11461\
        );

    \I__2756\ : InMux
    port map (
            O => \N__11481\,
            I => \N__11461\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__11478\,
            I => \N__11458\
        );

    \I__2754\ : Span4Mux_v
    port map (
            O => \N__11475\,
            I => \N__11455\
        );

    \I__2753\ : Span4Mux_h
    port map (
            O => \N__11468\,
            I => \N__11452\
        );

    \I__2752\ : InMux
    port map (
            O => \N__11467\,
            I => \N__11449\
        );

    \I__2751\ : InMux
    port map (
            O => \N__11466\,
            I => \N__11446\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__11461\,
            I => \N__11443\
        );

    \I__2749\ : Sp12to4
    port map (
            O => \N__11458\,
            I => \N__11440\
        );

    \I__2748\ : Span4Mux_v
    port map (
            O => \N__11455\,
            I => \N__11437\
        );

    \I__2747\ : Span4Mux_v
    port map (
            O => \N__11452\,
            I => \N__11434\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__11449\,
            I => \N__11429\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__11446\,
            I => \N__11429\
        );

    \I__2744\ : Span12Mux_v
    port map (
            O => \N__11443\,
            I => \N__11426\
        );

    \I__2743\ : Span12Mux_v
    port map (
            O => \N__11440\,
            I => \N__11423\
        );

    \I__2742\ : Sp12to4
    port map (
            O => \N__11437\,
            I => \N__11416\
        );

    \I__2741\ : Sp12to4
    port map (
            O => \N__11434\,
            I => \N__11416\
        );

    \I__2740\ : Span12Mux_v
    port map (
            O => \N__11429\,
            I => \N__11416\
        );

    \I__2739\ : Span12Mux_h
    port map (
            O => \N__11426\,
            I => \N__11413\
        );

    \I__2738\ : Span12Mux_h
    port map (
            O => \N__11423\,
            I => \N__11410\
        );

    \I__2737\ : Span12Mux_h
    port map (
            O => \N__11416\,
            I => \N__11407\
        );

    \I__2736\ : Odrv12
    port map (
            O => \N__11413\,
            I => \SIZ_c_1\
        );

    \I__2735\ : Odrv12
    port map (
            O => \N__11410\,
            I => \SIZ_c_1\
        );

    \I__2734\ : Odrv12
    port map (
            O => \N__11407\,
            I => \SIZ_c_1\
        );

    \I__2733\ : CascadeMux
    port map (
            O => \N__11400\,
            I => \N__11394\
        );

    \I__2732\ : InMux
    port map (
            O => \N__11399\,
            I => \N__11391\
        );

    \I__2731\ : InMux
    port map (
            O => \N__11398\,
            I => \N__11388\
        );

    \I__2730\ : InMux
    port map (
            O => \N__11397\,
            I => \N__11385\
        );

    \I__2729\ : InMux
    port map (
            O => \N__11394\,
            I => \N__11382\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__11391\,
            I => \N__11374\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__11388\,
            I => \N__11374\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__11385\,
            I => \N__11369\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__11382\,
            I => \N__11369\
        );

    \I__2724\ : CascadeMux
    port map (
            O => \N__11381\,
            I => \N__11365\
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__11380\,
            I => \N__11362\
        );

    \I__2722\ : CascadeMux
    port map (
            O => \N__11379\,
            I => \N__11359\
        );

    \I__2721\ : Span4Mux_v
    port map (
            O => \N__11374\,
            I => \N__11355\
        );

    \I__2720\ : Span4Mux_v
    port map (
            O => \N__11369\,
            I => \N__11352\
        );

    \I__2719\ : InMux
    port map (
            O => \N__11368\,
            I => \N__11349\
        );

    \I__2718\ : InMux
    port map (
            O => \N__11365\,
            I => \N__11344\
        );

    \I__2717\ : InMux
    port map (
            O => \N__11362\,
            I => \N__11344\
        );

    \I__2716\ : InMux
    port map (
            O => \N__11359\,
            I => \N__11340\
        );

    \I__2715\ : InMux
    port map (
            O => \N__11358\,
            I => \N__11337\
        );

    \I__2714\ : Span4Mux_v
    port map (
            O => \N__11355\,
            I => \N__11328\
        );

    \I__2713\ : Span4Mux_v
    port map (
            O => \N__11352\,
            I => \N__11328\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__11349\,
            I => \N__11328\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__11344\,
            I => \N__11328\
        );

    \I__2710\ : InMux
    port map (
            O => \N__11343\,
            I => \N__11325\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__11340\,
            I => \N__11322\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__11337\,
            I => \N__11319\
        );

    \I__2707\ : Span4Mux_h
    port map (
            O => \N__11328\,
            I => \N__11314\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__11325\,
            I => \N__11314\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__11322\,
            I => \N__11311\
        );

    \I__2704\ : Span4Mux_v
    port map (
            O => \N__11319\,
            I => \N__11308\
        );

    \I__2703\ : Span4Mux_h
    port map (
            O => \N__11314\,
            I => \N__11305\
        );

    \I__2702\ : Sp12to4
    port map (
            O => \N__11311\,
            I => \N__11302\
        );

    \I__2701\ : Span4Mux_v
    port map (
            O => \N__11308\,
            I => \N__11299\
        );

    \I__2700\ : Span4Mux_v
    port map (
            O => \N__11305\,
            I => \N__11296\
        );

    \I__2699\ : Span12Mux_h
    port map (
            O => \N__11302\,
            I => \N__11293\
        );

    \I__2698\ : Span4Mux_v
    port map (
            O => \N__11299\,
            I => \N__11290\
        );

    \I__2697\ : Span4Mux_h
    port map (
            O => \N__11296\,
            I => \N__11287\
        );

    \I__2696\ : Span12Mux_v
    port map (
            O => \N__11293\,
            I => \N__11284\
        );

    \I__2695\ : Sp12to4
    port map (
            O => \N__11290\,
            I => \N__11279\
        );

    \I__2694\ : Sp12to4
    port map (
            O => \N__11287\,
            I => \N__11279\
        );

    \I__2693\ : Odrv12
    port map (
            O => \N__11284\,
            I => \SIZ_c_0\
        );

    \I__2692\ : Odrv12
    port map (
            O => \N__11279\,
            I => \SIZ_c_0\
        );

    \I__2691\ : IoInMux
    port map (
            O => \N__11274\,
            I => \N__11271\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__11271\,
            I => \N__11268\
        );

    \I__2689\ : Span4Mux_s2_v
    port map (
            O => \N__11268\,
            I => \N__11265\
        );

    \I__2688\ : Span4Mux_v
    port map (
            O => \N__11265\,
            I => \N__11262\
        );

    \I__2687\ : Odrv4
    port map (
            O => \N__11262\,
            I => \N_334_i\
        );

    \I__2686\ : CascadeMux
    port map (
            O => \N__11259\,
            I => \N__11254\
        );

    \I__2685\ : InMux
    port map (
            O => \N__11258\,
            I => \N__11251\
        );

    \I__2684\ : InMux
    port map (
            O => \N__11257\,
            I => \N__11247\
        );

    \I__2683\ : InMux
    port map (
            O => \N__11254\,
            I => \N__11244\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__11251\,
            I => \N__11241\
        );

    \I__2681\ : InMux
    port map (
            O => \N__11250\,
            I => \N__11238\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__11247\,
            I => \N__11235\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__11244\,
            I => \N__11231\
        );

    \I__2678\ : Span4Mux_v
    port map (
            O => \N__11241\,
            I => \N__11228\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__11238\,
            I => \N__11225\
        );

    \I__2676\ : Span4Mux_v
    port map (
            O => \N__11235\,
            I => \N__11222\
        );

    \I__2675\ : InMux
    port map (
            O => \N__11234\,
            I => \N__11219\
        );

    \I__2674\ : Span4Mux_v
    port map (
            O => \N__11231\,
            I => \N__11216\
        );

    \I__2673\ : Span4Mux_v
    port map (
            O => \N__11228\,
            I => \N__11213\
        );

    \I__2672\ : Span4Mux_v
    port map (
            O => \N__11225\,
            I => \N__11210\
        );

    \I__2671\ : Sp12to4
    port map (
            O => \N__11222\,
            I => \N__11207\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__11219\,
            I => \N__11204\
        );

    \I__2669\ : Span4Mux_h
    port map (
            O => \N__11216\,
            I => \N__11201\
        );

    \I__2668\ : Span4Mux_v
    port map (
            O => \N__11213\,
            I => \N__11196\
        );

    \I__2667\ : Span4Mux_h
    port map (
            O => \N__11210\,
            I => \N__11196\
        );

    \I__2666\ : Span12Mux_h
    port map (
            O => \N__11207\,
            I => \N__11191\
        );

    \I__2665\ : Span12Mux_v
    port map (
            O => \N__11204\,
            I => \N__11191\
        );

    \I__2664\ : Sp12to4
    port map (
            O => \N__11201\,
            I => \N__11186\
        );

    \I__2663\ : Sp12to4
    port map (
            O => \N__11196\,
            I => \N__11186\
        );

    \I__2662\ : Span12Mux_h
    port map (
            O => \N__11191\,
            I => \N__11183\
        );

    \I__2661\ : Span12Mux_h
    port map (
            O => \N__11186\,
            I => \N__11180\
        );

    \I__2660\ : Odrv12
    port map (
            O => \N__11183\,
            I => \RnW_c\
        );

    \I__2659\ : Odrv12
    port map (
            O => \N__11180\,
            I => \RnW_c\
        );

    \I__2658\ : InMux
    port map (
            O => \N__11175\,
            I => \N__11171\
        );

    \I__2657\ : InMux
    port map (
            O => \N__11174\,
            I => \N__11168\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__11171\,
            I => \N__11165\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__11168\,
            I => \N__11162\
        );

    \I__2654\ : Span12Mux_s6_h
    port map (
            O => \N__11165\,
            I => \N__11159\
        );

    \I__2653\ : Sp12to4
    port map (
            O => \N__11162\,
            I => \N__11156\
        );

    \I__2652\ : Span12Mux_v
    port map (
            O => \N__11159\,
            I => \N__11150\
        );

    \I__2651\ : Span12Mux_v
    port map (
            O => \N__11156\,
            I => \N__11150\
        );

    \I__2650\ : InMux
    port map (
            O => \N__11155\,
            I => \N__11147\
        );

    \I__2649\ : Odrv12
    port map (
            O => \N__11150\,
            I => \DMA_WRITE_CYCLE\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__11147\,
            I => \DMA_WRITE_CYCLE\
        );

    \I__2647\ : IoInMux
    port map (
            O => \N__11142\,
            I => \N__11139\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__11139\,
            I => \N__11136\
        );

    \I__2645\ : IoSpan4Mux
    port map (
            O => \N__11136\,
            I => \N__11133\
        );

    \I__2644\ : Span4Mux_s3_h
    port map (
            O => \N__11133\,
            I => \N__11130\
        );

    \I__2643\ : Odrv4
    port map (
            O => \N__11130\,
            I => \N_379\
        );

    \I__2642\ : InMux
    port map (
            O => \N__11127\,
            I => \N__11124\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__11124\,
            I => \N__11117\
        );

    \I__2640\ : InMux
    port map (
            O => \N__11123\,
            I => \N__11114\
        );

    \I__2639\ : InMux
    port map (
            O => \N__11122\,
            I => \N__11111\
        );

    \I__2638\ : InMux
    port map (
            O => \N__11121\,
            I => \N__11105\
        );

    \I__2637\ : InMux
    port map (
            O => \N__11120\,
            I => \N__11105\
        );

    \I__2636\ : Sp12to4
    port map (
            O => \N__11117\,
            I => \N__11102\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__11114\,
            I => \N__11099\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__11111\,
            I => \N__11096\
        );

    \I__2633\ : InMux
    port map (
            O => \N__11110\,
            I => \N__11093\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__11105\,
            I => \N__11090\
        );

    \I__2631\ : Span12Mux_v
    port map (
            O => \N__11102\,
            I => \N__11087\
        );

    \I__2630\ : Span12Mux_h
    port map (
            O => \N__11099\,
            I => \N__11084\
        );

    \I__2629\ : Span12Mux_h
    port map (
            O => \N__11096\,
            I => \N__11079\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__11093\,
            I => \N__11079\
        );

    \I__2627\ : Span4Mux_h
    port map (
            O => \N__11090\,
            I => \N__11076\
        );

    \I__2626\ : Span12Mux_h
    port map (
            O => \N__11087\,
            I => \N__11073\
        );

    \I__2625\ : Span12Mux_v
    port map (
            O => \N__11084\,
            I => \N__11070\
        );

    \I__2624\ : Span12Mux_v
    port map (
            O => \N__11079\,
            I => \N__11067\
        );

    \I__2623\ : Span4Mux_v
    port map (
            O => \N__11076\,
            I => \N__11064\
        );

    \I__2622\ : Odrv12
    port map (
            O => \N__11073\,
            I => \CASUn_c\
        );

    \I__2621\ : Odrv12
    port map (
            O => \N__11070\,
            I => \CASUn_c\
        );

    \I__2620\ : Odrv12
    port map (
            O => \N__11067\,
            I => \CASUn_c\
        );

    \I__2619\ : Odrv4
    port map (
            O => \N__11064\,
            I => \CASUn_c\
        );

    \I__2618\ : InMux
    port map (
            O => \N__11055\,
            I => \N__11052\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__11052\,
            I => \N__11048\
        );

    \I__2616\ : InMux
    port map (
            O => \N__11051\,
            I => \N__11045\
        );

    \I__2615\ : Span4Mux_v
    port map (
            O => \N__11048\,
            I => \N__11040\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__11045\,
            I => \N__11037\
        );

    \I__2613\ : InMux
    port map (
            O => \N__11044\,
            I => \N__11034\
        );

    \I__2612\ : InMux
    port map (
            O => \N__11043\,
            I => \N__11031\
        );

    \I__2611\ : Span4Mux_v
    port map (
            O => \N__11040\,
            I => \N__11024\
        );

    \I__2610\ : Span4Mux_v
    port map (
            O => \N__11037\,
            I => \N__11024\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__11034\,
            I => \N__11024\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__11031\,
            I => \N__11021\
        );

    \I__2607\ : Span4Mux_v
    port map (
            O => \N__11024\,
            I => \N__11017\
        );

    \I__2606\ : Span4Mux_v
    port map (
            O => \N__11021\,
            I => \N__11014\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__11020\,
            I => \N__11010\
        );

    \I__2604\ : Span4Mux_v
    port map (
            O => \N__11017\,
            I => \N__11007\
        );

    \I__2603\ : Sp12to4
    port map (
            O => \N__11014\,
            I => \N__11004\
        );

    \I__2602\ : InMux
    port map (
            O => \N__11013\,
            I => \N__11001\
        );

    \I__2601\ : InMux
    port map (
            O => \N__11010\,
            I => \N__10998\
        );

    \I__2600\ : Sp12to4
    port map (
            O => \N__11007\,
            I => \N__10995\
        );

    \I__2599\ : Span12Mux_h
    port map (
            O => \N__11004\,
            I => \N__10988\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__11001\,
            I => \N__10988\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__10998\,
            I => \N__10988\
        );

    \I__2596\ : Span12Mux_h
    port map (
            O => \N__10995\,
            I => \N__10985\
        );

    \I__2595\ : Span12Mux_v
    port map (
            O => \N__10988\,
            I => \N__10982\
        );

    \I__2594\ : Odrv12
    port map (
            O => \N__10985\,
            I => \CASLn_c\
        );

    \I__2593\ : Odrv12
    port map (
            O => \N__10982\,
            I => \CASLn_c\
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__10977\,
            I => \N__10974\
        );

    \I__2591\ : InMux
    port map (
            O => \N__10974\,
            I => \N__10970\
        );

    \I__2590\ : InMux
    port map (
            O => \N__10973\,
            I => \N__10967\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__10970\,
            I => \N__10962\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__10967\,
            I => \N__10959\
        );

    \I__2587\ : InMux
    port map (
            O => \N__10966\,
            I => \N__10956\
        );

    \I__2586\ : InMux
    port map (
            O => \N__10965\,
            I => \N__10953\
        );

    \I__2585\ : Span4Mux_v
    port map (
            O => \N__10962\,
            I => \N__10941\
        );

    \I__2584\ : Span4Mux_v
    port map (
            O => \N__10959\,
            I => \N__10936\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__10956\,
            I => \N__10936\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__10953\,
            I => \N__10933\
        );

    \I__2581\ : InMux
    port map (
            O => \N__10952\,
            I => \N__10929\
        );

    \I__2580\ : InMux
    port map (
            O => \N__10951\,
            I => \N__10922\
        );

    \I__2579\ : InMux
    port map (
            O => \N__10950\,
            I => \N__10922\
        );

    \I__2578\ : InMux
    port map (
            O => \N__10949\,
            I => \N__10922\
        );

    \I__2577\ : InMux
    port map (
            O => \N__10948\,
            I => \N__10917\
        );

    \I__2576\ : InMux
    port map (
            O => \N__10947\,
            I => \N__10917\
        );

    \I__2575\ : InMux
    port map (
            O => \N__10946\,
            I => \N__10914\
        );

    \I__2574\ : CascadeMux
    port map (
            O => \N__10945\,
            I => \N__10911\
        );

    \I__2573\ : InMux
    port map (
            O => \N__10944\,
            I => \N__10906\
        );

    \I__2572\ : Sp12to4
    port map (
            O => \N__10941\,
            I => \N__10903\
        );

    \I__2571\ : Span4Mux_v
    port map (
            O => \N__10936\,
            I => \N__10900\
        );

    \I__2570\ : Span4Mux_v
    port map (
            O => \N__10933\,
            I => \N__10897\
        );

    \I__2569\ : InMux
    port map (
            O => \N__10932\,
            I => \N__10893\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__10929\,
            I => \N__10883\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__10922\,
            I => \N__10878\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__10917\,
            I => \N__10878\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__10914\,
            I => \N__10875\
        );

    \I__2564\ : InMux
    port map (
            O => \N__10911\,
            I => \N__10872\
        );

    \I__2563\ : InMux
    port map (
            O => \N__10910\,
            I => \N__10867\
        );

    \I__2562\ : InMux
    port map (
            O => \N__10909\,
            I => \N__10867\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__10906\,
            I => \N__10864\
        );

    \I__2560\ : Span12Mux_h
    port map (
            O => \N__10903\,
            I => \N__10861\
        );

    \I__2559\ : Span4Mux_h
    port map (
            O => \N__10900\,
            I => \N__10858\
        );

    \I__2558\ : Span4Mux_h
    port map (
            O => \N__10897\,
            I => \N__10855\
        );

    \I__2557\ : InMux
    port map (
            O => \N__10896\,
            I => \N__10852\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__10893\,
            I => \N__10849\
        );

    \I__2555\ : InMux
    port map (
            O => \N__10892\,
            I => \N__10844\
        );

    \I__2554\ : InMux
    port map (
            O => \N__10891\,
            I => \N__10844\
        );

    \I__2553\ : InMux
    port map (
            O => \N__10890\,
            I => \N__10841\
        );

    \I__2552\ : InMux
    port map (
            O => \N__10889\,
            I => \N__10832\
        );

    \I__2551\ : InMux
    port map (
            O => \N__10888\,
            I => \N__10832\
        );

    \I__2550\ : InMux
    port map (
            O => \N__10887\,
            I => \N__10832\
        );

    \I__2549\ : InMux
    port map (
            O => \N__10886\,
            I => \N__10832\
        );

    \I__2548\ : Span4Mux_v
    port map (
            O => \N__10883\,
            I => \N__10825\
        );

    \I__2547\ : Span4Mux_v
    port map (
            O => \N__10878\,
            I => \N__10825\
        );

    \I__2546\ : Span4Mux_h
    port map (
            O => \N__10875\,
            I => \N__10825\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__10872\,
            I => \N__10818\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__10867\,
            I => \N__10818\
        );

    \I__2543\ : Span4Mux_h
    port map (
            O => \N__10864\,
            I => \N__10818\
        );

    \I__2542\ : Odrv12
    port map (
            O => \N__10861\,
            I => \CPU_CYCLEm\
        );

    \I__2541\ : Odrv4
    port map (
            O => \N__10858\,
            I => \CPU_CYCLEm\
        );

    \I__2540\ : Odrv4
    port map (
            O => \N__10855\,
            I => \CPU_CYCLEm\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__10852\,
            I => \CPU_CYCLEm\
        );

    \I__2538\ : Odrv4
    port map (
            O => \N__10849\,
            I => \CPU_CYCLEm\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__10844\,
            I => \CPU_CYCLEm\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__10841\,
            I => \CPU_CYCLEm\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__10832\,
            I => \CPU_CYCLEm\
        );

    \I__2534\ : Odrv4
    port map (
            O => \N__10825\,
            I => \CPU_CYCLEm\
        );

    \I__2533\ : Odrv4
    port map (
            O => \N__10818\,
            I => \CPU_CYCLEm\
        );

    \I__2532\ : InMux
    port map (
            O => \N__10797\,
            I => \N__10792\
        );

    \I__2531\ : InMux
    port map (
            O => \N__10796\,
            I => \N__10789\
        );

    \I__2530\ : InMux
    port map (
            O => \N__10795\,
            I => \N__10786\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__10792\,
            I => \N__10782\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__10789\,
            I => \N__10777\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__10786\,
            I => \N__10777\
        );

    \I__2526\ : InMux
    port map (
            O => \N__10785\,
            I => \N__10774\
        );

    \I__2525\ : Span4Mux_h
    port map (
            O => \N__10782\,
            I => \N__10771\
        );

    \I__2524\ : Span4Mux_v
    port map (
            O => \N__10777\,
            I => \N__10766\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__10774\,
            I => \N__10766\
        );

    \I__2522\ : Sp12to4
    port map (
            O => \N__10771\,
            I => \N__10763\
        );

    \I__2521\ : Span4Mux_h
    port map (
            O => \N__10766\,
            I => \N__10760\
        );

    \I__2520\ : Span12Mux_v
    port map (
            O => \N__10763\,
            I => \N__10757\
        );

    \I__2519\ : Sp12to4
    port map (
            O => \N__10760\,
            I => \N__10754\
        );

    \I__2518\ : Span12Mux_h
    port map (
            O => \N__10757\,
            I => \N__10751\
        );

    \I__2517\ : Span12Mux_v
    port map (
            O => \N__10754\,
            I => \N__10748\
        );

    \I__2516\ : Odrv12
    port map (
            O => \N__10751\,
            I => \DRA_c_5\
        );

    \I__2515\ : Odrv12
    port map (
            O => \N__10748\,
            I => \DRA_c_5\
        );

    \I__2514\ : CascadeMux
    port map (
            O => \N__10743\,
            I => \N__10738\
        );

    \I__2513\ : CascadeMux
    port map (
            O => \N__10742\,
            I => \N__10730\
        );

    \I__2512\ : InMux
    port map (
            O => \N__10741\,
            I => \N__10726\
        );

    \I__2511\ : InMux
    port map (
            O => \N__10738\,
            I => \N__10723\
        );

    \I__2510\ : CascadeMux
    port map (
            O => \N__10737\,
            I => \N__10717\
        );

    \I__2509\ : InMux
    port map (
            O => \N__10736\,
            I => \N__10709\
        );

    \I__2508\ : InMux
    port map (
            O => \N__10735\,
            I => \N__10706\
        );

    \I__2507\ : InMux
    port map (
            O => \N__10734\,
            I => \N__10703\
        );

    \I__2506\ : InMux
    port map (
            O => \N__10733\,
            I => \N__10698\
        );

    \I__2505\ : InMux
    port map (
            O => \N__10730\,
            I => \N__10693\
        );

    \I__2504\ : InMux
    port map (
            O => \N__10729\,
            I => \N__10693\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__10726\,
            I => \N__10690\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__10723\,
            I => \N__10687\
        );

    \I__2501\ : InMux
    port map (
            O => \N__10722\,
            I => \N__10682\
        );

    \I__2500\ : InMux
    port map (
            O => \N__10721\,
            I => \N__10682\
        );

    \I__2499\ : InMux
    port map (
            O => \N__10720\,
            I => \N__10679\
        );

    \I__2498\ : InMux
    port map (
            O => \N__10717\,
            I => \N__10672\
        );

    \I__2497\ : InMux
    port map (
            O => \N__10716\,
            I => \N__10672\
        );

    \I__2496\ : InMux
    port map (
            O => \N__10715\,
            I => \N__10672\
        );

    \I__2495\ : InMux
    port map (
            O => \N__10714\,
            I => \N__10669\
        );

    \I__2494\ : InMux
    port map (
            O => \N__10713\,
            I => \N__10666\
        );

    \I__2493\ : InMux
    port map (
            O => \N__10712\,
            I => \N__10662\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__10709\,
            I => \N__10659\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__10706\,
            I => \N__10654\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__10703\,
            I => \N__10654\
        );

    \I__2489\ : InMux
    port map (
            O => \N__10702\,
            I => \N__10651\
        );

    \I__2488\ : InMux
    port map (
            O => \N__10701\,
            I => \N__10648\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__10698\,
            I => \N__10643\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__10693\,
            I => \N__10643\
        );

    \I__2485\ : Span4Mux_v
    port map (
            O => \N__10690\,
            I => \N__10631\
        );

    \I__2484\ : Span4Mux_v
    port map (
            O => \N__10687\,
            I => \N__10631\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__10682\,
            I => \N__10631\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__10679\,
            I => \N__10631\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__10672\,
            I => \N__10631\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__10669\,
            I => \N__10626\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__10666\,
            I => \N__10626\
        );

    \I__2478\ : InMux
    port map (
            O => \N__10665\,
            I => \N__10623\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__10662\,
            I => \N__10620\
        );

    \I__2476\ : Span4Mux_h
    port map (
            O => \N__10659\,
            I => \N__10617\
        );

    \I__2475\ : Span4Mux_v
    port map (
            O => \N__10654\,
            I => \N__10610\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__10651\,
            I => \N__10610\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__10648\,
            I => \N__10610\
        );

    \I__2472\ : Span4Mux_v
    port map (
            O => \N__10643\,
            I => \N__10607\
        );

    \I__2471\ : InMux
    port map (
            O => \N__10642\,
            I => \N__10604\
        );

    \I__2470\ : Span4Mux_h
    port map (
            O => \N__10631\,
            I => \N__10595\
        );

    \I__2469\ : Span4Mux_v
    port map (
            O => \N__10626\,
            I => \N__10595\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__10623\,
            I => \N__10595\
        );

    \I__2467\ : Span4Mux_v
    port map (
            O => \N__10620\,
            I => \N__10595\
        );

    \I__2466\ : Sp12to4
    port map (
            O => \N__10617\,
            I => \N__10592\
        );

    \I__2465\ : Sp12to4
    port map (
            O => \N__10610\,
            I => \N__10589\
        );

    \I__2464\ : Sp12to4
    port map (
            O => \N__10607\,
            I => \N__10582\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__10604\,
            I => \N__10582\
        );

    \I__2462\ : Sp12to4
    port map (
            O => \N__10595\,
            I => \N__10582\
        );

    \I__2461\ : Span12Mux_v
    port map (
            O => \N__10592\,
            I => \N__10579\
        );

    \I__2460\ : Span12Mux_v
    port map (
            O => \N__10589\,
            I => \N__10576\
        );

    \I__2459\ : Span12Mux_h
    port map (
            O => \N__10582\,
            I => \N__10573\
        );

    \I__2458\ : Span12Mux_h
    port map (
            O => \N__10579\,
            I => \N__10570\
        );

    \I__2457\ : Span12Mux_h
    port map (
            O => \N__10576\,
            I => \N__10565\
        );

    \I__2456\ : Span12Mux_v
    port map (
            O => \N__10573\,
            I => \N__10565\
        );

    \I__2455\ : Odrv12
    port map (
            O => \N__10570\,
            I => \AGNUS_REV_c\
        );

    \I__2454\ : Odrv12
    port map (
            O => \N__10565\,
            I => \AGNUS_REV_c\
        );

    \I__2453\ : InMux
    port map (
            O => \N__10560\,
            I => \N__10554\
        );

    \I__2452\ : InMux
    port map (
            O => \N__10559\,
            I => \N__10551\
        );

    \I__2451\ : InMux
    port map (
            O => \N__10558\,
            I => \N__10546\
        );

    \I__2450\ : InMux
    port map (
            O => \N__10557\,
            I => \N__10546\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__10554\,
            I => \N__10543\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__10551\,
            I => \N__10540\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__10546\,
            I => \N__10537\
        );

    \I__2446\ : Span4Mux_h
    port map (
            O => \N__10543\,
            I => \N__10532\
        );

    \I__2445\ : Span4Mux_v
    port map (
            O => \N__10540\,
            I => \N__10532\
        );

    \I__2444\ : Sp12to4
    port map (
            O => \N__10537\,
            I => \N__10529\
        );

    \I__2443\ : Span4Mux_v
    port map (
            O => \N__10532\,
            I => \N__10526\
        );

    \I__2442\ : Span12Mux_v
    port map (
            O => \N__10529\,
            I => \N__10521\
        );

    \I__2441\ : Sp12to4
    port map (
            O => \N__10526\,
            I => \N__10521\
        );

    \I__2440\ : Span12Mux_h
    port map (
            O => \N__10521\,
            I => \N__10518\
        );

    \I__2439\ : Odrv12
    port map (
            O => \N__10518\,
            I => \DRA_c_6\
        );

    \I__2438\ : InMux
    port map (
            O => \N__10515\,
            I => \N__10512\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__10512\,
            I => \N__10509\
        );

    \I__2436\ : Odrv12
    port map (
            O => \N__10509\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2435\ : CEMux
    port map (
            O => \N__10506\,
            I => \N__10464\
        );

    \I__2434\ : CEMux
    port map (
            O => \N__10505\,
            I => \N__10464\
        );

    \I__2433\ : CEMux
    port map (
            O => \N__10504\,
            I => \N__10464\
        );

    \I__2432\ : CEMux
    port map (
            O => \N__10503\,
            I => \N__10464\
        );

    \I__2431\ : CEMux
    port map (
            O => \N__10502\,
            I => \N__10464\
        );

    \I__2430\ : CEMux
    port map (
            O => \N__10501\,
            I => \N__10464\
        );

    \I__2429\ : CEMux
    port map (
            O => \N__10500\,
            I => \N__10464\
        );

    \I__2428\ : CEMux
    port map (
            O => \N__10499\,
            I => \N__10464\
        );

    \I__2427\ : CEMux
    port map (
            O => \N__10498\,
            I => \N__10464\
        );

    \I__2426\ : CEMux
    port map (
            O => \N__10497\,
            I => \N__10464\
        );

    \I__2425\ : CEMux
    port map (
            O => \N__10496\,
            I => \N__10464\
        );

    \I__2424\ : CEMux
    port map (
            O => \N__10495\,
            I => \N__10464\
        );

    \I__2423\ : CEMux
    port map (
            O => \N__10494\,
            I => \N__10464\
        );

    \I__2422\ : CEMux
    port map (
            O => \N__10493\,
            I => \N__10464\
        );

    \I__2421\ : GlobalMux
    port map (
            O => \N__10464\,
            I => \N__10461\
        );

    \I__2420\ : gio2CtrlBuf
    port map (
            O => \N__10461\,
            I => \DBRn_c_i_0_g\
        );

    \I__2419\ : InMux
    port map (
            O => \N__10458\,
            I => \N__10455\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__10455\,
            I => \N__10452\
        );

    \I__2417\ : Span12Mux_h
    port map (
            O => \N__10452\,
            I => \N__10449\
        );

    \I__2416\ : Odrv12
    port map (
            O => \N__10449\,
            I => \RAS1n_c\
        );

    \I__2415\ : InMux
    port map (
            O => \N__10446\,
            I => \N__10442\
        );

    \I__2414\ : InMux
    port map (
            O => \N__10445\,
            I => \N__10439\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__10442\,
            I => \N__10436\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__10439\,
            I => \N__10433\
        );

    \I__2411\ : Span4Mux_v
    port map (
            O => \N__10436\,
            I => \N__10428\
        );

    \I__2410\ : Span4Mux_v
    port map (
            O => \N__10433\,
            I => \N__10428\
        );

    \I__2409\ : Sp12to4
    port map (
            O => \N__10428\,
            I => \N__10425\
        );

    \I__2408\ : Span12Mux_h
    port map (
            O => \N__10425\,
            I => \N__10422\
        );

    \I__2407\ : Odrv12
    port map (
            O => \N__10422\,
            I => \RAS0n_c\
        );

    \I__2406\ : CascadeMux
    port map (
            O => \N__10419\,
            I => \N__10414\
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__10418\,
            I => \N__10411\
        );

    \I__2404\ : CascadeMux
    port map (
            O => \N__10417\,
            I => \N__10401\
        );

    \I__2403\ : InMux
    port map (
            O => \N__10414\,
            I => \N__10397\
        );

    \I__2402\ : InMux
    port map (
            O => \N__10411\,
            I => \N__10386\
        );

    \I__2401\ : InMux
    port map (
            O => \N__10410\,
            I => \N__10386\
        );

    \I__2400\ : InMux
    port map (
            O => \N__10409\,
            I => \N__10386\
        );

    \I__2399\ : InMux
    port map (
            O => \N__10408\,
            I => \N__10375\
        );

    \I__2398\ : InMux
    port map (
            O => \N__10407\,
            I => \N__10375\
        );

    \I__2397\ : CascadeMux
    port map (
            O => \N__10406\,
            I => \N__10372\
        );

    \I__2396\ : InMux
    port map (
            O => \N__10405\,
            I => \N__10367\
        );

    \I__2395\ : InMux
    port map (
            O => \N__10404\,
            I => \N__10367\
        );

    \I__2394\ : InMux
    port map (
            O => \N__10401\,
            I => \N__10364\
        );

    \I__2393\ : InMux
    port map (
            O => \N__10400\,
            I => \N__10361\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__10397\,
            I => \N__10358\
        );

    \I__2391\ : InMux
    port map (
            O => \N__10396\,
            I => \N__10351\
        );

    \I__2390\ : InMux
    port map (
            O => \N__10395\,
            I => \N__10351\
        );

    \I__2389\ : InMux
    port map (
            O => \N__10394\,
            I => \N__10351\
        );

    \I__2388\ : InMux
    port map (
            O => \N__10393\,
            I => \N__10347\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__10386\,
            I => \N__10344\
        );

    \I__2386\ : InMux
    port map (
            O => \N__10385\,
            I => \N__10341\
        );

    \I__2385\ : InMux
    port map (
            O => \N__10384\,
            I => \N__10338\
        );

    \I__2384\ : InMux
    port map (
            O => \N__10383\,
            I => \N__10335\
        );

    \I__2383\ : InMux
    port map (
            O => \N__10382\,
            I => \N__10328\
        );

    \I__2382\ : InMux
    port map (
            O => \N__10381\,
            I => \N__10328\
        );

    \I__2381\ : InMux
    port map (
            O => \N__10380\,
            I => \N__10328\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__10375\,
            I => \N__10322\
        );

    \I__2379\ : InMux
    port map (
            O => \N__10372\,
            I => \N__10319\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__10367\,
            I => \N__10312\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__10364\,
            I => \N__10312\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__10361\,
            I => \N__10309\
        );

    \I__2375\ : Span4Mux_h
    port map (
            O => \N__10358\,
            I => \N__10304\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__10351\,
            I => \N__10304\
        );

    \I__2373\ : InMux
    port map (
            O => \N__10350\,
            I => \N__10301\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__10347\,
            I => \N__10297\
        );

    \I__2371\ : Span4Mux_v
    port map (
            O => \N__10344\,
            I => \N__10286\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__10341\,
            I => \N__10286\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__10338\,
            I => \N__10286\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__10335\,
            I => \N__10286\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__10328\,
            I => \N__10286\
        );

    \I__2366\ : InMux
    port map (
            O => \N__10327\,
            I => \N__10283\
        );

    \I__2365\ : InMux
    port map (
            O => \N__10326\,
            I => \N__10280\
        );

    \I__2364\ : InMux
    port map (
            O => \N__10325\,
            I => \N__10277\
        );

    \I__2363\ : Span4Mux_h
    port map (
            O => \N__10322\,
            I => \N__10272\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__10319\,
            I => \N__10272\
        );

    \I__2361\ : InMux
    port map (
            O => \N__10318\,
            I => \N__10269\
        );

    \I__2360\ : InMux
    port map (
            O => \N__10317\,
            I => \N__10266\
        );

    \I__2359\ : Span4Mux_h
    port map (
            O => \N__10312\,
            I => \N__10257\
        );

    \I__2358\ : Span4Mux_v
    port map (
            O => \N__10309\,
            I => \N__10257\
        );

    \I__2357\ : Span4Mux_v
    port map (
            O => \N__10304\,
            I => \N__10257\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__10301\,
            I => \N__10257\
        );

    \I__2355\ : InMux
    port map (
            O => \N__10300\,
            I => \N__10254\
        );

    \I__2354\ : Span4Mux_v
    port map (
            O => \N__10297\,
            I => \N__10247\
        );

    \I__2353\ : Span4Mux_v
    port map (
            O => \N__10286\,
            I => \N__10247\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__10283\,
            I => \N__10240\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__10280\,
            I => \N__10240\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__10277\,
            I => \N__10240\
        );

    \I__2349\ : Span4Mux_h
    port map (
            O => \N__10272\,
            I => \N__10233\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__10269\,
            I => \N__10233\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__10266\,
            I => \N__10233\
        );

    \I__2346\ : Span4Mux_h
    port map (
            O => \N__10257\,
            I => \N__10226\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__10254\,
            I => \N__10226\
        );

    \I__2344\ : InMux
    port map (
            O => \N__10253\,
            I => \N__10221\
        );

    \I__2343\ : InMux
    port map (
            O => \N__10252\,
            I => \N__10221\
        );

    \I__2342\ : Span4Mux_h
    port map (
            O => \N__10247\,
            I => \N__10214\
        );

    \I__2341\ : Span4Mux_v
    port map (
            O => \N__10240\,
            I => \N__10214\
        );

    \I__2340\ : Span4Mux_v
    port map (
            O => \N__10233\,
            I => \N__10214\
        );

    \I__2339\ : InMux
    port map (
            O => \N__10232\,
            I => \N__10209\
        );

    \I__2338\ : InMux
    port map (
            O => \N__10231\,
            I => \N__10209\
        );

    \I__2337\ : Sp12to4
    port map (
            O => \N__10226\,
            I => \N__10206\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__10221\,
            I => \N__10199\
        );

    \I__2335\ : Sp12to4
    port map (
            O => \N__10214\,
            I => \N__10199\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__10209\,
            I => \N__10199\
        );

    \I__2333\ : Span12Mux_v
    port map (
            O => \N__10206\,
            I => \N__10196\
        );

    \I__2332\ : Span12Mux_h
    port map (
            O => \N__10199\,
            I => \N__10193\
        );

    \I__2331\ : Span12Mux_h
    port map (
            O => \N__10196\,
            I => \N__10190\
        );

    \I__2330\ : Odrv12
    port map (
            O => \N__10193\,
            I => \RESETn_c\
        );

    \I__2329\ : Odrv12
    port map (
            O => \N__10190\,
            I => \RESETn_c\
        );

    \I__2328\ : InMux
    port map (
            O => \N__10185\,
            I => \N__10182\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__10182\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2326\ : InMux
    port map (
            O => \N__10179\,
            I => \N__10176\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__10176\,
            I => \N__10173\
        );

    \I__2324\ : Odrv4
    port map (
            O => \N__10173\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__2323\ : IoInMux
    port map (
            O => \N__10170\,
            I => \N__10167\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__10167\,
            I => \N__10164\
        );

    \I__2321\ : Span4Mux_s1_v
    port map (
            O => \N__10164\,
            I => \N__10161\
        );

    \I__2320\ : Sp12to4
    port map (
            O => \N__10161\,
            I => \N__10158\
        );

    \I__2319\ : Span12Mux_h
    port map (
            O => \N__10158\,
            I => \N__10155\
        );

    \I__2318\ : Span12Mux_v
    port map (
            O => \N__10155\,
            I => \N__10151\
        );

    \I__2317\ : InMux
    port map (
            O => \N__10154\,
            I => \N__10148\
        );

    \I__2316\ : Odrv12
    port map (
            O => \N__10151\,
            I => \LDSn_c\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__10148\,
            I => \LDSn_c\
        );

    \I__2314\ : InMux
    port map (
            O => \N__10143\,
            I => \N__10140\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__10140\,
            I => \U712_REG_SM.N_459\
        );

    \I__2312\ : CascadeMux
    port map (
            O => \N__10137\,
            I => \N__10133\
        );

    \I__2311\ : InMux
    port map (
            O => \N__10136\,
            I => \N__10128\
        );

    \I__2310\ : InMux
    port map (
            O => \N__10133\,
            I => \N__10128\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__10128\,
            I => \N__10124\
        );

    \I__2308\ : InMux
    port map (
            O => \N__10127\,
            I => \N__10121\
        );

    \I__2307\ : Odrv12
    port map (
            O => \N__10124\,
            I => \U712_REG_SM.un1_REGENn_0_sqmuxa_0\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__10121\,
            I => \U712_REG_SM.un1_REGENn_0_sqmuxa_0\
        );

    \I__2305\ : InMux
    port map (
            O => \N__10116\,
            I => \N__10110\
        );

    \I__2304\ : InMux
    port map (
            O => \N__10115\,
            I => \N__10105\
        );

    \I__2303\ : InMux
    port map (
            O => \N__10114\,
            I => \N__10105\
        );

    \I__2302\ : CascadeMux
    port map (
            O => \N__10113\,
            I => \N__10093\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__10110\,
            I => \N__10088\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__10105\,
            I => \N__10088\
        );

    \I__2299\ : CascadeMux
    port map (
            O => \N__10104\,
            I => \N__10085\
        );

    \I__2298\ : InMux
    port map (
            O => \N__10103\,
            I => \N__10082\
        );

    \I__2297\ : InMux
    port map (
            O => \N__10102\,
            I => \N__10079\
        );

    \I__2296\ : InMux
    port map (
            O => \N__10101\,
            I => \N__10076\
        );

    \I__2295\ : InMux
    port map (
            O => \N__10100\,
            I => \N__10071\
        );

    \I__2294\ : InMux
    port map (
            O => \N__10099\,
            I => \N__10071\
        );

    \I__2293\ : InMux
    port map (
            O => \N__10098\,
            I => \N__10066\
        );

    \I__2292\ : InMux
    port map (
            O => \N__10097\,
            I => \N__10066\
        );

    \I__2291\ : CascadeMux
    port map (
            O => \N__10096\,
            I => \N__10062\
        );

    \I__2290\ : InMux
    port map (
            O => \N__10093\,
            I => \N__10059\
        );

    \I__2289\ : Span4Mux_h
    port map (
            O => \N__10088\,
            I => \N__10056\
        );

    \I__2288\ : InMux
    port map (
            O => \N__10085\,
            I => \N__10053\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__10082\,
            I => \N__10044\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__10079\,
            I => \N__10044\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__10076\,
            I => \N__10044\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__10071\,
            I => \N__10044\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__10066\,
            I => \N__10041\
        );

    \I__2282\ : InMux
    port map (
            O => \N__10065\,
            I => \N__10036\
        );

    \I__2281\ : InMux
    port map (
            O => \N__10062\,
            I => \N__10036\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__10059\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2279\ : Odrv4
    port map (
            O => \N__10056\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__10053\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2277\ : Odrv4
    port map (
            O => \N__10044\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2276\ : Odrv12
    port map (
            O => \N__10041\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__10036\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2274\ : IoInMux
    port map (
            O => \N__10023\,
            I => \N__10020\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__10020\,
            I => \N__10017\
        );

    \I__2272\ : IoSpan4Mux
    port map (
            O => \N__10017\,
            I => \N__10014\
        );

    \I__2271\ : Span4Mux_s2_v
    port map (
            O => \N__10014\,
            I => \N__10011\
        );

    \I__2270\ : Sp12to4
    port map (
            O => \N__10011\,
            I => \N__10007\
        );

    \I__2269\ : CascadeMux
    port map (
            O => \N__10010\,
            I => \N__10004\
        );

    \I__2268\ : Span12Mux_v
    port map (
            O => \N__10007\,
            I => \N__10001\
        );

    \I__2267\ : InMux
    port map (
            O => \N__10004\,
            I => \N__9998\
        );

    \I__2266\ : Odrv12
    port map (
            O => \N__10001\,
            I => \UDSn_c\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__9998\,
            I => \UDSn_c\
        );

    \I__2264\ : InMux
    port map (
            O => \N__9993\,
            I => \N__9990\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__9990\,
            I => \N__9950\
        );

    \I__2262\ : ClkMux
    port map (
            O => \N__9989\,
            I => \N__9831\
        );

    \I__2261\ : ClkMux
    port map (
            O => \N__9988\,
            I => \N__9831\
        );

    \I__2260\ : ClkMux
    port map (
            O => \N__9987\,
            I => \N__9831\
        );

    \I__2259\ : ClkMux
    port map (
            O => \N__9986\,
            I => \N__9831\
        );

    \I__2258\ : ClkMux
    port map (
            O => \N__9985\,
            I => \N__9831\
        );

    \I__2257\ : ClkMux
    port map (
            O => \N__9984\,
            I => \N__9831\
        );

    \I__2256\ : ClkMux
    port map (
            O => \N__9983\,
            I => \N__9831\
        );

    \I__2255\ : ClkMux
    port map (
            O => \N__9982\,
            I => \N__9831\
        );

    \I__2254\ : ClkMux
    port map (
            O => \N__9981\,
            I => \N__9831\
        );

    \I__2253\ : ClkMux
    port map (
            O => \N__9980\,
            I => \N__9831\
        );

    \I__2252\ : ClkMux
    port map (
            O => \N__9979\,
            I => \N__9831\
        );

    \I__2251\ : ClkMux
    port map (
            O => \N__9978\,
            I => \N__9831\
        );

    \I__2250\ : ClkMux
    port map (
            O => \N__9977\,
            I => \N__9831\
        );

    \I__2249\ : ClkMux
    port map (
            O => \N__9976\,
            I => \N__9831\
        );

    \I__2248\ : ClkMux
    port map (
            O => \N__9975\,
            I => \N__9831\
        );

    \I__2247\ : ClkMux
    port map (
            O => \N__9974\,
            I => \N__9831\
        );

    \I__2246\ : ClkMux
    port map (
            O => \N__9973\,
            I => \N__9831\
        );

    \I__2245\ : ClkMux
    port map (
            O => \N__9972\,
            I => \N__9831\
        );

    \I__2244\ : ClkMux
    port map (
            O => \N__9971\,
            I => \N__9831\
        );

    \I__2243\ : ClkMux
    port map (
            O => \N__9970\,
            I => \N__9831\
        );

    \I__2242\ : ClkMux
    port map (
            O => \N__9969\,
            I => \N__9831\
        );

    \I__2241\ : ClkMux
    port map (
            O => \N__9968\,
            I => \N__9831\
        );

    \I__2240\ : ClkMux
    port map (
            O => \N__9967\,
            I => \N__9831\
        );

    \I__2239\ : ClkMux
    port map (
            O => \N__9966\,
            I => \N__9831\
        );

    \I__2238\ : ClkMux
    port map (
            O => \N__9965\,
            I => \N__9831\
        );

    \I__2237\ : ClkMux
    port map (
            O => \N__9964\,
            I => \N__9831\
        );

    \I__2236\ : ClkMux
    port map (
            O => \N__9963\,
            I => \N__9831\
        );

    \I__2235\ : ClkMux
    port map (
            O => \N__9962\,
            I => \N__9831\
        );

    \I__2234\ : ClkMux
    port map (
            O => \N__9961\,
            I => \N__9831\
        );

    \I__2233\ : ClkMux
    port map (
            O => \N__9960\,
            I => \N__9831\
        );

    \I__2232\ : ClkMux
    port map (
            O => \N__9959\,
            I => \N__9831\
        );

    \I__2231\ : ClkMux
    port map (
            O => \N__9958\,
            I => \N__9831\
        );

    \I__2230\ : ClkMux
    port map (
            O => \N__9957\,
            I => \N__9831\
        );

    \I__2229\ : ClkMux
    port map (
            O => \N__9956\,
            I => \N__9831\
        );

    \I__2228\ : ClkMux
    port map (
            O => \N__9955\,
            I => \N__9831\
        );

    \I__2227\ : ClkMux
    port map (
            O => \N__9954\,
            I => \N__9831\
        );

    \I__2226\ : ClkMux
    port map (
            O => \N__9953\,
            I => \N__9831\
        );

    \I__2225\ : Glb2LocalMux
    port map (
            O => \N__9950\,
            I => \N__9831\
        );

    \I__2224\ : ClkMux
    port map (
            O => \N__9949\,
            I => \N__9831\
        );

    \I__2223\ : ClkMux
    port map (
            O => \N__9948\,
            I => \N__9831\
        );

    \I__2222\ : ClkMux
    port map (
            O => \N__9947\,
            I => \N__9831\
        );

    \I__2221\ : ClkMux
    port map (
            O => \N__9946\,
            I => \N__9831\
        );

    \I__2220\ : ClkMux
    port map (
            O => \N__9945\,
            I => \N__9831\
        );

    \I__2219\ : ClkMux
    port map (
            O => \N__9944\,
            I => \N__9831\
        );

    \I__2218\ : ClkMux
    port map (
            O => \N__9943\,
            I => \N__9831\
        );

    \I__2217\ : ClkMux
    port map (
            O => \N__9942\,
            I => \N__9831\
        );

    \I__2216\ : ClkMux
    port map (
            O => \N__9941\,
            I => \N__9831\
        );

    \I__2215\ : ClkMux
    port map (
            O => \N__9940\,
            I => \N__9831\
        );

    \I__2214\ : ClkMux
    port map (
            O => \N__9939\,
            I => \N__9831\
        );

    \I__2213\ : ClkMux
    port map (
            O => \N__9938\,
            I => \N__9831\
        );

    \I__2212\ : ClkMux
    port map (
            O => \N__9937\,
            I => \N__9831\
        );

    \I__2211\ : ClkMux
    port map (
            O => \N__9936\,
            I => \N__9831\
        );

    \I__2210\ : GlobalMux
    port map (
            O => \N__9831\,
            I => \CLK80_PLL\
        );

    \I__2209\ : InMux
    port map (
            O => \N__9828\,
            I => \N__9820\
        );

    \I__2208\ : InMux
    port map (
            O => \N__9827\,
            I => \N__9817\
        );

    \I__2207\ : InMux
    port map (
            O => \N__9826\,
            I => \N__9814\
        );

    \I__2206\ : InMux
    port map (
            O => \N__9825\,
            I => \N__9811\
        );

    \I__2205\ : InMux
    port map (
            O => \N__9824\,
            I => \N__9808\
        );

    \I__2204\ : InMux
    port map (
            O => \N__9823\,
            I => \N__9805\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__9820\,
            I => \N__9802\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__9817\,
            I => \N__9796\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__9814\,
            I => \N__9788\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__9811\,
            I => \N__9781\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__9808\,
            I => \N__9770\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__9805\,
            I => \N__9746\
        );

    \I__2197\ : Glb2LocalMux
    port map (
            O => \N__9802\,
            I => \N__9642\
        );

    \I__2196\ : SRMux
    port map (
            O => \N__9801\,
            I => \N__9642\
        );

    \I__2195\ : SRMux
    port map (
            O => \N__9800\,
            I => \N__9642\
        );

    \I__2194\ : SRMux
    port map (
            O => \N__9799\,
            I => \N__9642\
        );

    \I__2193\ : Glb2LocalMux
    port map (
            O => \N__9796\,
            I => \N__9642\
        );

    \I__2192\ : SRMux
    port map (
            O => \N__9795\,
            I => \N__9642\
        );

    \I__2191\ : SRMux
    port map (
            O => \N__9794\,
            I => \N__9642\
        );

    \I__2190\ : SRMux
    port map (
            O => \N__9793\,
            I => \N__9642\
        );

    \I__2189\ : SRMux
    port map (
            O => \N__9792\,
            I => \N__9642\
        );

    \I__2188\ : SRMux
    port map (
            O => \N__9791\,
            I => \N__9642\
        );

    \I__2187\ : Glb2LocalMux
    port map (
            O => \N__9788\,
            I => \N__9642\
        );

    \I__2186\ : SRMux
    port map (
            O => \N__9787\,
            I => \N__9642\
        );

    \I__2185\ : SRMux
    port map (
            O => \N__9786\,
            I => \N__9642\
        );

    \I__2184\ : SRMux
    port map (
            O => \N__9785\,
            I => \N__9642\
        );

    \I__2183\ : SRMux
    port map (
            O => \N__9784\,
            I => \N__9642\
        );

    \I__2182\ : Glb2LocalMux
    port map (
            O => \N__9781\,
            I => \N__9642\
        );

    \I__2181\ : SRMux
    port map (
            O => \N__9780\,
            I => \N__9642\
        );

    \I__2180\ : SRMux
    port map (
            O => \N__9779\,
            I => \N__9642\
        );

    \I__2179\ : SRMux
    port map (
            O => \N__9778\,
            I => \N__9642\
        );

    \I__2178\ : SRMux
    port map (
            O => \N__9777\,
            I => \N__9642\
        );

    \I__2177\ : SRMux
    port map (
            O => \N__9776\,
            I => \N__9642\
        );

    \I__2176\ : SRMux
    port map (
            O => \N__9775\,
            I => \N__9642\
        );

    \I__2175\ : SRMux
    port map (
            O => \N__9774\,
            I => \N__9642\
        );

    \I__2174\ : SRMux
    port map (
            O => \N__9773\,
            I => \N__9642\
        );

    \I__2173\ : Glb2LocalMux
    port map (
            O => \N__9770\,
            I => \N__9642\
        );

    \I__2172\ : SRMux
    port map (
            O => \N__9769\,
            I => \N__9642\
        );

    \I__2171\ : SRMux
    port map (
            O => \N__9768\,
            I => \N__9642\
        );

    \I__2170\ : SRMux
    port map (
            O => \N__9767\,
            I => \N__9642\
        );

    \I__2169\ : SRMux
    port map (
            O => \N__9766\,
            I => \N__9642\
        );

    \I__2168\ : SRMux
    port map (
            O => \N__9765\,
            I => \N__9642\
        );

    \I__2167\ : SRMux
    port map (
            O => \N__9764\,
            I => \N__9642\
        );

    \I__2166\ : SRMux
    port map (
            O => \N__9763\,
            I => \N__9642\
        );

    \I__2165\ : SRMux
    port map (
            O => \N__9762\,
            I => \N__9642\
        );

    \I__2164\ : SRMux
    port map (
            O => \N__9761\,
            I => \N__9642\
        );

    \I__2163\ : SRMux
    port map (
            O => \N__9760\,
            I => \N__9642\
        );

    \I__2162\ : SRMux
    port map (
            O => \N__9759\,
            I => \N__9642\
        );

    \I__2161\ : SRMux
    port map (
            O => \N__9758\,
            I => \N__9642\
        );

    \I__2160\ : SRMux
    port map (
            O => \N__9757\,
            I => \N__9642\
        );

    \I__2159\ : SRMux
    port map (
            O => \N__9756\,
            I => \N__9642\
        );

    \I__2158\ : SRMux
    port map (
            O => \N__9755\,
            I => \N__9642\
        );

    \I__2157\ : SRMux
    port map (
            O => \N__9754\,
            I => \N__9642\
        );

    \I__2156\ : SRMux
    port map (
            O => \N__9753\,
            I => \N__9642\
        );

    \I__2155\ : SRMux
    port map (
            O => \N__9752\,
            I => \N__9642\
        );

    \I__2154\ : SRMux
    port map (
            O => \N__9751\,
            I => \N__9642\
        );

    \I__2153\ : SRMux
    port map (
            O => \N__9750\,
            I => \N__9642\
        );

    \I__2152\ : SRMux
    port map (
            O => \N__9749\,
            I => \N__9642\
        );

    \I__2151\ : Glb2LocalMux
    port map (
            O => \N__9746\,
            I => \N__9642\
        );

    \I__2150\ : SRMux
    port map (
            O => \N__9745\,
            I => \N__9642\
        );

    \I__2149\ : SRMux
    port map (
            O => \N__9744\,
            I => \N__9642\
        );

    \I__2148\ : SRMux
    port map (
            O => \N__9743\,
            I => \N__9642\
        );

    \I__2147\ : GlobalMux
    port map (
            O => \N__9642\,
            I => \N__9639\
        );

    \I__2146\ : gio2CtrlBuf
    port map (
            O => \N__9639\,
            I => \RESETn_c_i_g\
        );

    \I__2145\ : InMux
    port map (
            O => \N__9636\,
            I => \N__9633\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__9633\,
            I => \U712_REG_SM.N_404\
        );

    \I__2143\ : IoInMux
    port map (
            O => \N__9630\,
            I => \N__9627\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__9627\,
            I => \N__9624\
        );

    \I__2141\ : Span4Mux_s0_v
    port map (
            O => \N__9624\,
            I => \N__9621\
        );

    \I__2140\ : Span4Mux_v
    port map (
            O => \N__9621\,
            I => \N__9618\
        );

    \I__2139\ : Odrv4
    port map (
            O => \N__9618\,
            I => \N_335_i\
        );

    \I__2138\ : IoInMux
    port map (
            O => \N__9615\,
            I => \N__9612\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__9612\,
            I => \N__9609\
        );

    \I__2136\ : Span4Mux_s3_v
    port map (
            O => \N__9609\,
            I => \N__9606\
        );

    \I__2135\ : Odrv4
    port map (
            O => \N__9606\,
            I => \N_337_i\
        );

    \I__2134\ : InMux
    port map (
            O => \N__9603\,
            I => \N__9598\
        );

    \I__2133\ : InMux
    port map (
            O => \N__9602\,
            I => \N__9593\
        );

    \I__2132\ : InMux
    port map (
            O => \N__9601\,
            I => \N__9593\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__9598\,
            I => \N__9590\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__9593\,
            I => \N__9586\
        );

    \I__2129\ : Span4Mux_v
    port map (
            O => \N__9590\,
            I => \N__9583\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9589\,
            I => \N__9580\
        );

    \I__2127\ : Span4Mux_h
    port map (
            O => \N__9586\,
            I => \N__9577\
        );

    \I__2126\ : Sp12to4
    port map (
            O => \N__9583\,
            I => \N__9574\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__9580\,
            I => \N__9569\
        );

    \I__2124\ : Sp12to4
    port map (
            O => \N__9577\,
            I => \N__9569\
        );

    \I__2123\ : Span12Mux_h
    port map (
            O => \N__9574\,
            I => \N__9566\
        );

    \I__2122\ : Span12Mux_v
    port map (
            O => \N__9569\,
            I => \N__9563\
        );

    \I__2121\ : Span12Mux_v
    port map (
            O => \N__9566\,
            I => \N__9560\
        );

    \I__2120\ : Span12Mux_h
    port map (
            O => \N__9563\,
            I => \N__9557\
        );

    \I__2119\ : Odrv12
    port map (
            O => \N__9560\,
            I => \DRA_c_3\
        );

    \I__2118\ : Odrv12
    port map (
            O => \N__9557\,
            I => \DRA_c_3\
        );

    \I__2117\ : InMux
    port map (
            O => \N__9552\,
            I => \N__9548\
        );

    \I__2116\ : InMux
    port map (
            O => \N__9551\,
            I => \N__9545\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__9548\,
            I => \N__9538\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__9545\,
            I => \N__9538\
        );

    \I__2113\ : InMux
    port map (
            O => \N__9544\,
            I => \N__9535\
        );

    \I__2112\ : InMux
    port map (
            O => \N__9543\,
            I => \N__9532\
        );

    \I__2111\ : Span4Mux_v
    port map (
            O => \N__9538\,
            I => \N__9529\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__9535\,
            I => \N__9526\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__9532\,
            I => \N__9521\
        );

    \I__2108\ : Sp12to4
    port map (
            O => \N__9529\,
            I => \N__9521\
        );

    \I__2107\ : Span12Mux_h
    port map (
            O => \N__9526\,
            I => \N__9518\
        );

    \I__2106\ : Span12Mux_h
    port map (
            O => \N__9521\,
            I => \N__9515\
        );

    \I__2105\ : Span12Mux_v
    port map (
            O => \N__9518\,
            I => \N__9512\
        );

    \I__2104\ : Span12Mux_v
    port map (
            O => \N__9515\,
            I => \N__9509\
        );

    \I__2103\ : Odrv12
    port map (
            O => \N__9512\,
            I => \DRA_c_2\
        );

    \I__2102\ : Odrv12
    port map (
            O => \N__9509\,
            I => \DRA_c_2\
        );

    \I__2101\ : InMux
    port map (
            O => \N__9504\,
            I => \N__9501\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__9501\,
            I => \N__9498\
        );

    \I__2099\ : Odrv4
    port map (
            O => \N__9498\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__2098\ : InMux
    port map (
            O => \N__9495\,
            I => \N__9490\
        );

    \I__2097\ : InMux
    port map (
            O => \N__9494\,
            I => \N__9487\
        );

    \I__2096\ : InMux
    port map (
            O => \N__9493\,
            I => \N__9484\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__9490\,
            I => \N__9480\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__9487\,
            I => \N__9475\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__9484\,
            I => \N__9475\
        );

    \I__2092\ : InMux
    port map (
            O => \N__9483\,
            I => \N__9472\
        );

    \I__2091\ : Span4Mux_v
    port map (
            O => \N__9480\,
            I => \N__9469\
        );

    \I__2090\ : Sp12to4
    port map (
            O => \N__9475\,
            I => \N__9464\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__9472\,
            I => \N__9464\
        );

    \I__2088\ : Sp12to4
    port map (
            O => \N__9469\,
            I => \N__9461\
        );

    \I__2087\ : Span12Mux_v
    port map (
            O => \N__9464\,
            I => \N__9458\
        );

    \I__2086\ : Span12Mux_h
    port map (
            O => \N__9461\,
            I => \N__9455\
        );

    \I__2085\ : Span12Mux_h
    port map (
            O => \N__9458\,
            I => \N__9452\
        );

    \I__2084\ : Odrv12
    port map (
            O => \N__9455\,
            I => \DRA_c_8\
        );

    \I__2083\ : Odrv12
    port map (
            O => \N__9452\,
            I => \DRA_c_8\
        );

    \I__2082\ : InMux
    port map (
            O => \N__9447\,
            I => \N__9444\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__9444\,
            I => \N__9441\
        );

    \I__2080\ : Span4Mux_h
    port map (
            O => \N__9441\,
            I => \N__9438\
        );

    \I__2079\ : Odrv4
    port map (
            O => \N__9438\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__2078\ : IoInMux
    port map (
            O => \N__9435\,
            I => \N__9432\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__9432\,
            I => \N__9429\
        );

    \I__2076\ : IoSpan4Mux
    port map (
            O => \N__9429\,
            I => \N__9426\
        );

    \I__2075\ : Sp12to4
    port map (
            O => \N__9426\,
            I => \N__9423\
        );

    \I__2074\ : Span12Mux_v
    port map (
            O => \N__9423\,
            I => \N__9420\
        );

    \I__2073\ : Span12Mux_h
    port map (
            O => \N__9420\,
            I => \N__9417\
        );

    \I__2072\ : Odrv12
    port map (
            O => \N__9417\,
            I => \ASn_c\
        );

    \I__2071\ : CEMux
    port map (
            O => \N__9414\,
            I => \N__9411\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__9411\,
            I => \U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0\
        );

    \I__2069\ : IoInMux
    port map (
            O => \N__9408\,
            I => \N__9405\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__9405\,
            I => \N__9402\
        );

    \I__2067\ : Span4Mux_s3_v
    port map (
            O => \N__9402\,
            I => \N__9399\
        );

    \I__2066\ : Odrv4
    port map (
            O => \N__9399\,
            I => \N_336_i\
        );

    \I__2065\ : InMux
    port map (
            O => \N__9396\,
            I => \N__9393\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__9393\,
            I => \N__9389\
        );

    \I__2063\ : InMux
    port map (
            O => \N__9392\,
            I => \N__9386\
        );

    \I__2062\ : Span4Mux_v
    port map (
            O => \N__9389\,
            I => \N__9383\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__9386\,
            I => \N__9380\
        );

    \I__2060\ : Span4Mux_v
    port map (
            O => \N__9383\,
            I => \N__9377\
        );

    \I__2059\ : Span4Mux_v
    port map (
            O => \N__9380\,
            I => \N__9374\
        );

    \I__2058\ : Sp12to4
    port map (
            O => \N__9377\,
            I => \N__9371\
        );

    \I__2057\ : Sp12to4
    port map (
            O => \N__9374\,
            I => \N__9368\
        );

    \I__2056\ : Span12Mux_h
    port map (
            O => \N__9371\,
            I => \N__9365\
        );

    \I__2055\ : Span12Mux_v
    port map (
            O => \N__9368\,
            I => \N__9362\
        );

    \I__2054\ : Span12Mux_v
    port map (
            O => \N__9365\,
            I => \N__9359\
        );

    \I__2053\ : Span12Mux_h
    port map (
            O => \N__9362\,
            I => \N__9356\
        );

    \I__2052\ : Odrv12
    port map (
            O => \N__9359\,
            I => \DRA_c_0\
        );

    \I__2051\ : Odrv12
    port map (
            O => \N__9356\,
            I => \DRA_c_0\
        );

    \I__2050\ : InMux
    port map (
            O => \N__9351\,
            I => \N__9346\
        );

    \I__2049\ : InMux
    port map (
            O => \N__9350\,
            I => \N__9343\
        );

    \I__2048\ : InMux
    port map (
            O => \N__9349\,
            I => \N__9340\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__9346\,
            I => \N__9336\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__9343\,
            I => \N__9331\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__9340\,
            I => \N__9331\
        );

    \I__2044\ : InMux
    port map (
            O => \N__9339\,
            I => \N__9328\
        );

    \I__2043\ : Span4Mux_v
    port map (
            O => \N__9336\,
            I => \N__9325\
        );

    \I__2042\ : Span4Mux_h
    port map (
            O => \N__9331\,
            I => \N__9320\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__9328\,
            I => \N__9320\
        );

    \I__2040\ : Span4Mux_h
    port map (
            O => \N__9325\,
            I => \N__9317\
        );

    \I__2039\ : Span4Mux_h
    port map (
            O => \N__9320\,
            I => \N__9314\
        );

    \I__2038\ : Sp12to4
    port map (
            O => \N__9317\,
            I => \N__9311\
        );

    \I__2037\ : Span4Mux_v
    port map (
            O => \N__9314\,
            I => \N__9308\
        );

    \I__2036\ : Span12Mux_s10_h
    port map (
            O => \N__9311\,
            I => \N__9303\
        );

    \I__2035\ : Sp12to4
    port map (
            O => \N__9308\,
            I => \N__9303\
        );

    \I__2034\ : Span12Mux_v
    port map (
            O => \N__9303\,
            I => \N__9300\
        );

    \I__2033\ : Odrv12
    port map (
            O => \N__9300\,
            I => \DRA_c_1\
        );

    \I__2032\ : InMux
    port map (
            O => \N__9297\,
            I => \N__9294\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__9294\,
            I => \N__9291\
        );

    \I__2030\ : Odrv12
    port map (
            O => \N__9291\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9288\,
            I => \N__9283\
        );

    \I__2028\ : InMux
    port map (
            O => \N__9287\,
            I => \N__9279\
        );

    \I__2027\ : InMux
    port map (
            O => \N__9286\,
            I => \N__9276\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__9283\,
            I => \N__9273\
        );

    \I__2025\ : InMux
    port map (
            O => \N__9282\,
            I => \N__9270\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__9279\,
            I => \N__9265\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__9276\,
            I => \N__9265\
        );

    \I__2022\ : Span4Mux_v
    port map (
            O => \N__9273\,
            I => \N__9262\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__9270\,
            I => \N__9259\
        );

    \I__2020\ : Span4Mux_v
    port map (
            O => \N__9265\,
            I => \N__9256\
        );

    \I__2019\ : Span4Mux_v
    port map (
            O => \N__9262\,
            I => \N__9251\
        );

    \I__2018\ : Span4Mux_v
    port map (
            O => \N__9259\,
            I => \N__9251\
        );

    \I__2017\ : Span4Mux_v
    port map (
            O => \N__9256\,
            I => \N__9248\
        );

    \I__2016\ : Sp12to4
    port map (
            O => \N__9251\,
            I => \N__9243\
        );

    \I__2015\ : Sp12to4
    port map (
            O => \N__9248\,
            I => \N__9243\
        );

    \I__2014\ : Span12Mux_h
    port map (
            O => \N__9243\,
            I => \N__9240\
        );

    \I__2013\ : Span12Mux_v
    port map (
            O => \N__9240\,
            I => \N__9237\
        );

    \I__2012\ : Odrv12
    port map (
            O => \N__9237\,
            I => \DRA_c_9\
        );

    \I__2011\ : InMux
    port map (
            O => \N__9234\,
            I => \N__9231\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__9231\,
            I => \N__9228\
        );

    \I__2009\ : Span4Mux_h
    port map (
            O => \N__9228\,
            I => \N__9225\
        );

    \I__2008\ : Odrv4
    port map (
            O => \N__9225\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2007\ : ClkMux
    port map (
            O => \N__9222\,
            I => \N__9201\
        );

    \I__2006\ : ClkMux
    port map (
            O => \N__9221\,
            I => \N__9201\
        );

    \I__2005\ : ClkMux
    port map (
            O => \N__9220\,
            I => \N__9201\
        );

    \I__2004\ : ClkMux
    port map (
            O => \N__9219\,
            I => \N__9201\
        );

    \I__2003\ : ClkMux
    port map (
            O => \N__9218\,
            I => \N__9201\
        );

    \I__2002\ : ClkMux
    port map (
            O => \N__9217\,
            I => \N__9201\
        );

    \I__2001\ : ClkMux
    port map (
            O => \N__9216\,
            I => \N__9201\
        );

    \I__2000\ : GlobalMux
    port map (
            O => \N__9201\,
            I => \N__9198\
        );

    \I__1999\ : gio2CtrlBuf
    port map (
            O => \N__9198\,
            I => \C3_c_g\
        );

    \I__1998\ : IoInMux
    port map (
            O => \N__9195\,
            I => \N__9192\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__9192\,
            I => \N__9189\
        );

    \I__1996\ : Span12Mux_s6_v
    port map (
            O => \N__9189\,
            I => \N__9186\
        );

    \I__1995\ : Odrv12
    port map (
            O => \N__9186\,
            I => \RESETn_c_i\
        );

    \I__1994\ : CascadeMux
    port map (
            O => \N__9183\,
            I => \N__9180\
        );

    \I__1993\ : InMux
    port map (
            O => \N__9180\,
            I => \N__9177\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__9177\,
            I => \N__9174\
        );

    \I__1991\ : Odrv12
    port map (
            O => \N__9174\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__1990\ : InMux
    port map (
            O => \N__9171\,
            I => \N__9167\
        );

    \I__1989\ : InMux
    port map (
            O => \N__9170\,
            I => \N__9164\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__9167\,
            I => \N__9158\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__9164\,
            I => \N__9158\
        );

    \I__1986\ : InMux
    port map (
            O => \N__9163\,
            I => \N__9155\
        );

    \I__1985\ : Span4Mux_v
    port map (
            O => \N__9158\,
            I => \N__9151\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__9155\,
            I => \N__9148\
        );

    \I__1983\ : InMux
    port map (
            O => \N__9154\,
            I => \N__9145\
        );

    \I__1982\ : Sp12to4
    port map (
            O => \N__9151\,
            I => \N__9142\
        );

    \I__1981\ : Sp12to4
    port map (
            O => \N__9148\,
            I => \N__9137\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__9145\,
            I => \N__9137\
        );

    \I__1979\ : Span12Mux_h
    port map (
            O => \N__9142\,
            I => \N__9134\
        );

    \I__1978\ : Span12Mux_v
    port map (
            O => \N__9137\,
            I => \N__9131\
        );

    \I__1977\ : Span12Mux_v
    port map (
            O => \N__9134\,
            I => \N__9126\
        );

    \I__1976\ : Span12Mux_h
    port map (
            O => \N__9131\,
            I => \N__9126\
        );

    \I__1975\ : Odrv12
    port map (
            O => \N__9126\,
            I => \DRA_c_4\
        );

    \I__1974\ : InMux
    port map (
            O => \N__9123\,
            I => \N__9120\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__9120\,
            I => \N__9117\
        );

    \I__1972\ : Span4Mux_h
    port map (
            O => \N__9117\,
            I => \N__9114\
        );

    \I__1971\ : Odrv4
    port map (
            O => \N__9114\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__1970\ : InMux
    port map (
            O => \N__9111\,
            I => \N__9108\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__9108\,
            I => \N__9105\
        );

    \I__1968\ : Span4Mux_h
    port map (
            O => \N__9105\,
            I => \N__9102\
        );

    \I__1967\ : Odrv4
    port map (
            O => \N__9102\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__1966\ : InMux
    port map (
            O => \N__9099\,
            I => \N__9096\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__9096\,
            I => \N__9093\
        );

    \I__1964\ : Odrv12
    port map (
            O => \N__9093\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__1963\ : InMux
    port map (
            O => \N__9090\,
            I => \N__9087\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__9087\,
            I => \N__9084\
        );

    \I__1961\ : Odrv12
    port map (
            O => \N__9084\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__1960\ : InMux
    port map (
            O => \N__9081\,
            I => \N__9078\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__9078\,
            I => \N__9075\
        );

    \I__1958\ : Span4Mux_v
    port map (
            O => \N__9075\,
            I => \N__9072\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__9072\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__1956\ : InMux
    port map (
            O => \N__9069\,
            I => \N__9063\
        );

    \I__1955\ : InMux
    port map (
            O => \N__9068\,
            I => \N__9060\
        );

    \I__1954\ : InMux
    port map (
            O => \N__9067\,
            I => \N__9057\
        );

    \I__1953\ : InMux
    port map (
            O => \N__9066\,
            I => \N__9054\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__9063\,
            I => \N__9049\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__9060\,
            I => \N__9049\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__9057\,
            I => \N__9044\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__9054\,
            I => \N__9044\
        );

    \I__1948\ : Span4Mux_v
    port map (
            O => \N__9049\,
            I => \N__9039\
        );

    \I__1947\ : Span4Mux_v
    port map (
            O => \N__9044\,
            I => \N__9039\
        );

    \I__1946\ : Sp12to4
    port map (
            O => \N__9039\,
            I => \N__9036\
        );

    \I__1945\ : Span12Mux_h
    port map (
            O => \N__9036\,
            I => \N__9033\
        );

    \I__1944\ : Odrv12
    port map (
            O => \N__9033\,
            I => \DRA_c_7\
        );

    \I__1943\ : InMux
    port map (
            O => \N__9030\,
            I => \N__9027\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__9027\,
            I => \N__9024\
        );

    \I__1941\ : Odrv4
    port map (
            O => \N__9024\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__1940\ : InMux
    port map (
            O => \N__9021\,
            I => \N__9018\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__9018\,
            I => \N__9015\
        );

    \I__1938\ : Odrv12
    port map (
            O => \N__9015\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\
        );

    \I__1937\ : InMux
    port map (
            O => \N__9012\,
            I => \N__9009\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__9009\,
            I => \U712_REG_SM.N_373\
        );

    \I__1935\ : CascadeMux
    port map (
            O => \N__9006\,
            I => \U712_REG_SM.N_330_cascade_\
        );

    \I__1934\ : InMux
    port map (
            O => \N__9003\,
            I => \N__9000\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__9000\,
            I => \U712_REG_SM.N_413\
        );

    \I__1932\ : InMux
    port map (
            O => \N__8997\,
            I => \N__8990\
        );

    \I__1931\ : InMux
    port map (
            O => \N__8996\,
            I => \N__8987\
        );

    \I__1930\ : InMux
    port map (
            O => \N__8995\,
            I => \N__8984\
        );

    \I__1929\ : InMux
    port map (
            O => \N__8994\,
            I => \N__8979\
        );

    \I__1928\ : InMux
    port map (
            O => \N__8993\,
            I => \N__8979\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__8990\,
            I => \N__8976\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__8987\,
            I => \N__8973\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__8984\,
            I => \N__8968\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__8979\,
            I => \N__8968\
        );

    \I__1923\ : Odrv4
    port map (
            O => \N__8976\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1922\ : Odrv4
    port map (
            O => \N__8973\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1921\ : Odrv4
    port map (
            O => \N__8968\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1920\ : InMux
    port map (
            O => \N__8961\,
            I => \N__8958\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__8958\,
            I => \U712_REG_SM.N_410\
        );

    \I__1918\ : CascadeMux
    port map (
            O => \N__8955\,
            I => \N__8950\
        );

    \I__1917\ : InMux
    port map (
            O => \N__8954\,
            I => \N__8942\
        );

    \I__1916\ : InMux
    port map (
            O => \N__8953\,
            I => \N__8942\
        );

    \I__1915\ : InMux
    port map (
            O => \N__8950\,
            I => \N__8942\
        );

    \I__1914\ : InMux
    port map (
            O => \N__8949\,
            I => \N__8939\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__8942\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__8939\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1911\ : InMux
    port map (
            O => \N__8934\,
            I => \N__8931\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__8931\,
            I => \U712_REG_SM.STATE_COUNTc_0_0\
        );

    \I__1909\ : InMux
    port map (
            O => \N__8928\,
            I => \N__8925\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8925\,
            I => \U712_REG_SM.N_308\
        );

    \I__1907\ : InMux
    port map (
            O => \N__8922\,
            I => \N__8918\
        );

    \I__1906\ : InMux
    port map (
            O => \N__8921\,
            I => \N__8915\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__8918\,
            I => \N__8906\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__8915\,
            I => \N__8906\
        );

    \I__1903\ : InMux
    port map (
            O => \N__8914\,
            I => \N__8903\
        );

    \I__1902\ : InMux
    port map (
            O => \N__8913\,
            I => \N__8898\
        );

    \I__1901\ : InMux
    port map (
            O => \N__8912\,
            I => \N__8898\
        );

    \I__1900\ : InMux
    port map (
            O => \N__8911\,
            I => \N__8895\
        );

    \I__1899\ : Odrv4
    port map (
            O => \N__8906\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__8903\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__8898\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__8895\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1895\ : CascadeMux
    port map (
            O => \N__8886\,
            I => \U712_REG_SM.N_308_cascade_\
        );

    \I__1894\ : InMux
    port map (
            O => \N__8883\,
            I => \N__8878\
        );

    \I__1893\ : InMux
    port map (
            O => \N__8882\,
            I => \N__8873\
        );

    \I__1892\ : InMux
    port map (
            O => \N__8881\,
            I => \N__8870\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__8878\,
            I => \N__8867\
        );

    \I__1890\ : InMux
    port map (
            O => \N__8877\,
            I => \N__8862\
        );

    \I__1889\ : InMux
    port map (
            O => \N__8876\,
            I => \N__8862\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__8873\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__8870\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1886\ : Odrv4
    port map (
            O => \N__8867\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__8862\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1884\ : CascadeMux
    port map (
            O => \N__8853\,
            I => \N__8849\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__8852\,
            I => \N__8838\
        );

    \I__1882\ : InMux
    port map (
            O => \N__8849\,
            I => \N__8833\
        );

    \I__1881\ : InMux
    port map (
            O => \N__8848\,
            I => \N__8830\
        );

    \I__1880\ : InMux
    port map (
            O => \N__8847\,
            I => \N__8825\
        );

    \I__1879\ : InMux
    port map (
            O => \N__8846\,
            I => \N__8825\
        );

    \I__1878\ : InMux
    port map (
            O => \N__8845\,
            I => \N__8822\
        );

    \I__1877\ : InMux
    port map (
            O => \N__8844\,
            I => \N__8819\
        );

    \I__1876\ : InMux
    port map (
            O => \N__8843\,
            I => \N__8810\
        );

    \I__1875\ : InMux
    port map (
            O => \N__8842\,
            I => \N__8810\
        );

    \I__1874\ : InMux
    port map (
            O => \N__8841\,
            I => \N__8810\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8838\,
            I => \N__8810\
        );

    \I__1872\ : InMux
    port map (
            O => \N__8837\,
            I => \N__8805\
        );

    \I__1871\ : InMux
    port map (
            O => \N__8836\,
            I => \N__8805\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__8833\,
            I => \N__8796\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__8830\,
            I => \N__8796\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__8825\,
            I => \N__8796\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__8822\,
            I => \N__8796\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__8819\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__8810\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__8805\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1863\ : Odrv4
    port map (
            O => \N__8796\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__8787\,
            I => \N__8782\
        );

    \I__1861\ : CascadeMux
    port map (
            O => \N__8786\,
            I => \N__8779\
        );

    \I__1860\ : InMux
    port map (
            O => \N__8785\,
            I => \N__8773\
        );

    \I__1859\ : InMux
    port map (
            O => \N__8782\,
            I => \N__8770\
        );

    \I__1858\ : InMux
    port map (
            O => \N__8779\,
            I => \N__8767\
        );

    \I__1857\ : InMux
    port map (
            O => \N__8778\,
            I => \N__8762\
        );

    \I__1856\ : InMux
    port map (
            O => \N__8777\,
            I => \N__8762\
        );

    \I__1855\ : InMux
    port map (
            O => \N__8776\,
            I => \N__8759\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__8773\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__8770\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__8767\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__8762\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__8759\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__1849\ : InMux
    port map (
            O => \N__8748\,
            I => \N__8745\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__8745\,
            I => \N__8742\
        );

    \I__1847\ : Span4Mux_h
    port map (
            O => \N__8742\,
            I => \N__8739\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__8739\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__1845\ : InMux
    port map (
            O => \N__8736\,
            I => \N__8733\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__8733\,
            I => \N__8730\
        );

    \I__1843\ : Odrv4
    port map (
            O => \N__8730\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1842\ : InMux
    port map (
            O => \N__8727\,
            I => \N__8724\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__8724\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1840\ : InMux
    port map (
            O => \N__8721\,
            I => \N__8718\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__8718\,
            I => \U712_CYCLE_TERM.N_332\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8715\,
            I => \N__8705\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8714\,
            I => \N__8705\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8713\,
            I => \N__8705\
        );

    \I__1835\ : CascadeMux
    port map (
            O => \N__8712\,
            I => \N__8702\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__8705\,
            I => \N__8699\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8702\,
            I => \N__8696\
        );

    \I__1832\ : Span4Mux_h
    port map (
            O => \N__8699\,
            I => \N__8693\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__8696\,
            I => \CPU_TACKm\
        );

    \I__1830\ : Odrv4
    port map (
            O => \N__8693\,
            I => \CPU_TACKm\
        );

    \I__1829\ : InMux
    port map (
            O => \N__8688\,
            I => \N__8682\
        );

    \I__1828\ : InMux
    port map (
            O => \N__8687\,
            I => \N__8675\
        );

    \I__1827\ : InMux
    port map (
            O => \N__8686\,
            I => \N__8675\
        );

    \I__1826\ : InMux
    port map (
            O => \N__8685\,
            I => \N__8675\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__8682\,
            I => \REG_TACK\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__8675\,
            I => \REG_TACK\
        );

    \I__1823\ : CascadeMux
    port map (
            O => \N__8670\,
            I => \N__8667\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8667\,
            I => \N__8662\
        );

    \I__1821\ : InMux
    port map (
            O => \N__8666\,
            I => \N__8657\
        );

    \I__1820\ : InMux
    port map (
            O => \N__8665\,
            I => \N__8657\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__8662\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__8657\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1817\ : CascadeMux
    port map (
            O => \N__8652\,
            I => \U712_CYCLE_TERM.N_455_cascade_\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8649\,
            I => \N__8645\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8648\,
            I => \N__8642\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__8645\,
            I => \N__8637\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__8642\,
            I => \N__8634\
        );

    \I__1812\ : InMux
    port map (
            O => \N__8641\,
            I => \N__8631\
        );

    \I__1811\ : InMux
    port map (
            O => \N__8640\,
            I => \N__8628\
        );

    \I__1810\ : Odrv4
    port map (
            O => \N__8637\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1809\ : Odrv4
    port map (
            O => \N__8634\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__8631\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__8628\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1806\ : InMux
    port map (
            O => \N__8619\,
            I => \N__8616\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__8616\,
            I => \N__8612\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8615\,
            I => \N__8609\
        );

    \I__1803\ : Span4Mux_v
    port map (
            O => \N__8612\,
            I => \N__8606\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8609\,
            I => \N__8603\
        );

    \I__1801\ : Span4Mux_h
    port map (
            O => \N__8606\,
            I => \N__8598\
        );

    \I__1800\ : Span4Mux_h
    port map (
            O => \N__8603\,
            I => \N__8598\
        );

    \I__1799\ : Odrv4
    port map (
            O => \N__8598\,
            I => \DBRn_c_i\
        );

    \I__1798\ : InMux
    port map (
            O => \N__8595\,
            I => \N__8591\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__8594\,
            I => \N__8588\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__8591\,
            I => \N__8585\
        );

    \I__1795\ : InMux
    port map (
            O => \N__8588\,
            I => \N__8582\
        );

    \I__1794\ : Span4Mux_h
    port map (
            O => \N__8585\,
            I => \N__8579\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__8582\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1792\ : Odrv4
    port map (
            O => \N__8579\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8574\,
            I => \N__8570\
        );

    \I__1790\ : InMux
    port map (
            O => \N__8573\,
            I => \N__8565\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__8570\,
            I => \N__8562\
        );

    \I__1788\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8559\
        );

    \I__1787\ : InMux
    port map (
            O => \N__8568\,
            I => \N__8556\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__8565\,
            I => \N__8553\
        );

    \I__1785\ : Span4Mux_v
    port map (
            O => \N__8562\,
            I => \N__8550\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__8559\,
            I => \N__8543\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__8556\,
            I => \N__8543\
        );

    \I__1782\ : Span4Mux_h
    port map (
            O => \N__8553\,
            I => \N__8543\
        );

    \I__1781\ : Span4Mux_v
    port map (
            O => \N__8550\,
            I => \N__8540\
        );

    \I__1780\ : Span4Mux_v
    port map (
            O => \N__8543\,
            I => \N__8537\
        );

    \I__1779\ : Span4Mux_v
    port map (
            O => \N__8540\,
            I => \N__8534\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__8537\,
            I => \N__8531\
        );

    \I__1777\ : IoSpan4Mux
    port map (
            O => \N__8534\,
            I => \N__8528\
        );

    \I__1776\ : Span4Mux_v
    port map (
            O => \N__8531\,
            I => \N__8525\
        );

    \I__1775\ : Odrv4
    port map (
            O => \N__8528\,
            I => \CLK40_PLL_i\
        );

    \I__1774\ : Odrv4
    port map (
            O => \N__8525\,
            I => \CLK40_PLL_i\
        );

    \I__1773\ : IoInMux
    port map (
            O => \N__8520\,
            I => \N__8517\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__8517\,
            I => \N__8514\
        );

    \I__1771\ : IoSpan4Mux
    port map (
            O => \N__8514\,
            I => \N__8510\
        );

    \I__1770\ : IoInMux
    port map (
            O => \N__8513\,
            I => \N__8507\
        );

    \I__1769\ : Span4Mux_s3_h
    port map (
            O => \N__8510\,
            I => \N__8502\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__8507\,
            I => \N__8502\
        );

    \I__1767\ : Span4Mux_s2_v
    port map (
            O => \N__8502\,
            I => \N__8499\
        );

    \I__1766\ : Span4Mux_v
    port map (
            O => \N__8499\,
            I => \N__8495\
        );

    \I__1765\ : IoInMux
    port map (
            O => \N__8498\,
            I => \N__8492\
        );

    \I__1764\ : Sp12to4
    port map (
            O => \N__8495\,
            I => \N__8489\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__8492\,
            I => \N__8486\
        );

    \I__1762\ : Span12Mux_h
    port map (
            O => \N__8489\,
            I => \N__8483\
        );

    \I__1761\ : Span12Mux_s9_h
    port map (
            O => \N__8486\,
            I => \N__8480\
        );

    \I__1760\ : Odrv12
    port map (
            O => \N__8483\,
            I => \CLK40_PLL_i_i\
        );

    \I__1759\ : Odrv12
    port map (
            O => \N__8480\,
            I => \CLK40_PLL_i_i\
        );

    \I__1758\ : InMux
    port map (
            O => \N__8475\,
            I => \N__8472\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__8472\,
            I => \U712_REG_SM.N_412\
        );

    \I__1756\ : InMux
    port map (
            O => \N__8469\,
            I => \N__8465\
        );

    \I__1755\ : IoInMux
    port map (
            O => \N__8468\,
            I => \N__8462\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__8465\,
            I => \N__8459\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__8462\,
            I => \N__8456\
        );

    \I__1752\ : Sp12to4
    port map (
            O => \N__8459\,
            I => \N__8453\
        );

    \I__1751\ : IoSpan4Mux
    port map (
            O => \N__8456\,
            I => \N__8450\
        );

    \I__1750\ : Span12Mux_v
    port map (
            O => \N__8453\,
            I => \N__8447\
        );

    \I__1749\ : IoSpan4Mux
    port map (
            O => \N__8450\,
            I => \N__8444\
        );

    \I__1748\ : Span12Mux_h
    port map (
            O => \N__8447\,
            I => \N__8441\
        );

    \I__1747\ : IoSpan4Mux
    port map (
            O => \N__8444\,
            I => \N__8438\
        );

    \I__1746\ : Odrv12
    port map (
            O => \N__8441\,
            I => \C1_c\
        );

    \I__1745\ : Odrv4
    port map (
            O => \N__8438\,
            I => \C1_c\
        );

    \I__1744\ : InMux
    port map (
            O => \N__8433\,
            I => \N__8430\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__8430\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1742\ : InMux
    port map (
            O => \N__8427\,
            I => \N__8424\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__8424\,
            I => \N__8421\
        );

    \I__1740\ : Odrv4
    port map (
            O => \N__8421\,
            I => \U712_REG_SM.REGENn_e_1\
        );

    \I__1739\ : InMux
    port map (
            O => \N__8418\,
            I => \N__8415\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__8415\,
            I => \N__8411\
        );

    \I__1737\ : InMux
    port map (
            O => \N__8414\,
            I => \N__8408\
        );

    \I__1736\ : Odrv4
    port map (
            O => \N__8411\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__8408\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__1734\ : IoInMux
    port map (
            O => \N__8403\,
            I => \N__8400\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__8400\,
            I => \N__8397\
        );

    \I__1732\ : Span4Mux_s0_v
    port map (
            O => \N__8397\,
            I => \N__8394\
        );

    \I__1731\ : Sp12to4
    port map (
            O => \N__8394\,
            I => \N__8390\
        );

    \I__1730\ : InMux
    port map (
            O => \N__8393\,
            I => \N__8386\
        );

    \I__1729\ : Span12Mux_h
    port map (
            O => \N__8390\,
            I => \N__8383\
        );

    \I__1728\ : InMux
    port map (
            O => \N__8389\,
            I => \N__8380\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__8386\,
            I => \N__8377\
        );

    \I__1726\ : Odrv12
    port map (
            O => \N__8383\,
            I => \REGENn_c\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__8380\,
            I => \REGENn_c\
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__8377\,
            I => \REGENn_c\
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__8370\,
            I => \N__8362\
        );

    \I__1722\ : CascadeMux
    port map (
            O => \N__8369\,
            I => \N__8359\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__8368\,
            I => \N__8355\
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__8367\,
            I => \N__8350\
        );

    \I__1719\ : InMux
    port map (
            O => \N__8366\,
            I => \N__8347\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8365\,
            I => \N__8342\
        );

    \I__1717\ : InMux
    port map (
            O => \N__8362\,
            I => \N__8342\
        );

    \I__1716\ : InMux
    port map (
            O => \N__8359\,
            I => \N__8339\
        );

    \I__1715\ : InMux
    port map (
            O => \N__8358\,
            I => \N__8335\
        );

    \I__1714\ : InMux
    port map (
            O => \N__8355\,
            I => \N__8321\
        );

    \I__1713\ : InMux
    port map (
            O => \N__8354\,
            I => \N__8321\
        );

    \I__1712\ : InMux
    port map (
            O => \N__8353\,
            I => \N__8321\
        );

    \I__1711\ : InMux
    port map (
            O => \N__8350\,
            I => \N__8321\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__8347\,
            I => \N__8316\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__8342\,
            I => \N__8316\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__8339\,
            I => \N__8310\
        );

    \I__1707\ : CascadeMux
    port map (
            O => \N__8338\,
            I => \N__8307\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__8335\,
            I => \N__8301\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8334\,
            I => \N__8298\
        );

    \I__1704\ : InMux
    port map (
            O => \N__8333\,
            I => \N__8291\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8332\,
            I => \N__8291\
        );

    \I__1702\ : InMux
    port map (
            O => \N__8331\,
            I => \N__8291\
        );

    \I__1701\ : CascadeMux
    port map (
            O => \N__8330\,
            I => \N__8287\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8321\,
            I => \N__8279\
        );

    \I__1699\ : Span4Mux_v
    port map (
            O => \N__8316\,
            I => \N__8279\
        );

    \I__1698\ : InMux
    port map (
            O => \N__8315\,
            I => \N__8272\
        );

    \I__1697\ : InMux
    port map (
            O => \N__8314\,
            I => \N__8272\
        );

    \I__1696\ : InMux
    port map (
            O => \N__8313\,
            I => \N__8272\
        );

    \I__1695\ : Span4Mux_h
    port map (
            O => \N__8310\,
            I => \N__8269\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8307\,
            I => \N__8260\
        );

    \I__1693\ : InMux
    port map (
            O => \N__8306\,
            I => \N__8260\
        );

    \I__1692\ : InMux
    port map (
            O => \N__8305\,
            I => \N__8260\
        );

    \I__1691\ : InMux
    port map (
            O => \N__8304\,
            I => \N__8260\
        );

    \I__1690\ : Span4Mux_v
    port map (
            O => \N__8301\,
            I => \N__8257\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__8298\,
            I => \N__8252\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__8291\,
            I => \N__8252\
        );

    \I__1687\ : InMux
    port map (
            O => \N__8290\,
            I => \N__8241\
        );

    \I__1686\ : InMux
    port map (
            O => \N__8287\,
            I => \N__8241\
        );

    \I__1685\ : InMux
    port map (
            O => \N__8286\,
            I => \N__8241\
        );

    \I__1684\ : InMux
    port map (
            O => \N__8285\,
            I => \N__8241\
        );

    \I__1683\ : InMux
    port map (
            O => \N__8284\,
            I => \N__8241\
        );

    \I__1682\ : Odrv4
    port map (
            O => \N__8279\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__8272\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1680\ : Odrv4
    port map (
            O => \N__8269\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__8260\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1678\ : Odrv4
    port map (
            O => \N__8257\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1677\ : Odrv4
    port map (
            O => \N__8252\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__8241\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1675\ : IoInMux
    port map (
            O => \N__8226\,
            I => \N__8223\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__8223\,
            I => \N__8220\
        );

    \I__1673\ : Span12Mux_s8_v
    port map (
            O => \N__8220\,
            I => \N__8217\
        );

    \I__1672\ : Span12Mux_h
    port map (
            O => \N__8217\,
            I => \N__8214\
        );

    \I__1671\ : Odrv12
    port map (
            O => \N__8214\,
            I => \CASn_c\
        );

    \I__1670\ : InMux
    port map (
            O => \N__8211\,
            I => \N__8208\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__8208\,
            I => \N__8205\
        );

    \I__1668\ : Odrv4
    port map (
            O => \N__8205\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1667\ : InMux
    port map (
            O => \N__8202\,
            I => \N__8199\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__8199\,
            I => \N__8195\
        );

    \I__1665\ : InMux
    port map (
            O => \N__8198\,
            I => \N__8192\
        );

    \I__1664\ : Span4Mux_v
    port map (
            O => \N__8195\,
            I => \N__8187\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__8192\,
            I => \N__8187\
        );

    \I__1662\ : Odrv4
    port map (
            O => \N__8187\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__1661\ : InMux
    port map (
            O => \N__8184\,
            I => \N__8181\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__8181\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__1659\ : InMux
    port map (
            O => \N__8178\,
            I => \N__8175\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__8175\,
            I => \N__8172\
        );

    \I__1657\ : Odrv4
    port map (
            O => \N__8172\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__1656\ : IoInMux
    port map (
            O => \N__8169\,
            I => \N__8166\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__8166\,
            I => \N__8163\
        );

    \I__1654\ : IoSpan4Mux
    port map (
            O => \N__8163\,
            I => \N__8160\
        );

    \I__1653\ : Span4Mux_s3_h
    port map (
            O => \N__8160\,
            I => \N__8157\
        );

    \I__1652\ : Span4Mux_h
    port map (
            O => \N__8157\,
            I => \N__8154\
        );

    \I__1651\ : Sp12to4
    port map (
            O => \N__8154\,
            I => \N__8150\
        );

    \I__1650\ : InMux
    port map (
            O => \N__8153\,
            I => \N__8147\
        );

    \I__1649\ : Span12Mux_h
    port map (
            O => \N__8150\,
            I => \N__8142\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__8147\,
            I => \N__8142\
        );

    \I__1647\ : Span12Mux_h
    port map (
            O => \N__8142\,
            I => \N__8139\
        );

    \I__1646\ : Span12Mux_v
    port map (
            O => \N__8139\,
            I => \N__8136\
        );

    \I__1645\ : Odrv12
    port map (
            O => \N__8136\,
            I => \C3_c\
        );

    \I__1644\ : InMux
    port map (
            O => \N__8133\,
            I => \N__8129\
        );

    \I__1643\ : InMux
    port map (
            O => \N__8132\,
            I => \N__8126\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__8129\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__8126\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__1640\ : InMux
    port map (
            O => \N__8121\,
            I => \N__8118\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__8118\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1638\ : CascadeMux
    port map (
            O => \N__8115\,
            I => \U712_REG_SM.N_328_cascade_\
        );

    \I__1637\ : CascadeMux
    port map (
            O => \N__8112\,
            I => \U712_REG_SM.N_331_cascade_\
        );

    \I__1636\ : InMux
    port map (
            O => \N__8109\,
            I => \N__8103\
        );

    \I__1635\ : InMux
    port map (
            O => \N__8108\,
            I => \N__8100\
        );

    \I__1634\ : InMux
    port map (
            O => \N__8107\,
            I => \N__8095\
        );

    \I__1633\ : InMux
    port map (
            O => \N__8106\,
            I => \N__8095\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__8103\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__8100\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__8095\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1629\ : InMux
    port map (
            O => \N__8088\,
            I => \N__8083\
        );

    \I__1628\ : InMux
    port map (
            O => \N__8087\,
            I => \N__8080\
        );

    \I__1627\ : InMux
    port map (
            O => \N__8086\,
            I => \N__8077\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__8083\,
            I => \N__8074\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__8080\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__8077\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__1623\ : Odrv4
    port map (
            O => \N__8074\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__8067\,
            I => \N__8063\
        );

    \I__1621\ : InMux
    port map (
            O => \N__8066\,
            I => \N__8060\
        );

    \I__1620\ : InMux
    port map (
            O => \N__8063\,
            I => \N__8057\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__8060\,
            I => \N__8054\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__8057\,
            I => \U712_REG_SM.N_328\
        );

    \I__1617\ : Odrv4
    port map (
            O => \N__8054\,
            I => \U712_REG_SM.N_328\
        );

    \I__1616\ : IoInMux
    port map (
            O => \N__8049\,
            I => \N__8046\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__8046\,
            I => \N__8042\
        );

    \I__1614\ : IoInMux
    port map (
            O => \N__8045\,
            I => \N__8039\
        );

    \I__1613\ : IoSpan4Mux
    port map (
            O => \N__8042\,
            I => \N__8036\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__8039\,
            I => \N__8032\
        );

    \I__1611\ : Span4Mux_s2_v
    port map (
            O => \N__8036\,
            I => \N__8029\
        );

    \I__1610\ : IoInMux
    port map (
            O => \N__8035\,
            I => \N__8026\
        );

    \I__1609\ : IoSpan4Mux
    port map (
            O => \N__8032\,
            I => \N__8023\
        );

    \I__1608\ : Sp12to4
    port map (
            O => \N__8029\,
            I => \N__8020\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__8026\,
            I => \N__8017\
        );

    \I__1606\ : Span4Mux_s3_v
    port map (
            O => \N__8023\,
            I => \N__8014\
        );

    \I__1605\ : Span12Mux_h
    port map (
            O => \N__8020\,
            I => \N__8011\
        );

    \I__1604\ : Span12Mux_s7_h
    port map (
            O => \N__8017\,
            I => \N__8008\
        );

    \I__1603\ : Sp12to4
    port map (
            O => \N__8014\,
            I => \N__8005\
        );

    \I__1602\ : Span12Mux_v
    port map (
            O => \N__8011\,
            I => \N__7997\
        );

    \I__1601\ : Span12Mux_v
    port map (
            O => \N__8008\,
            I => \N__7997\
        );

    \I__1600\ : Span12Mux_v
    port map (
            O => \N__8005\,
            I => \N__7997\
        );

    \I__1599\ : InMux
    port map (
            O => \N__8004\,
            I => \N__7994\
        );

    \I__1598\ : Odrv12
    port map (
            O => \N__7997\,
            I => \TACK_EN\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__7994\,
            I => \TACK_EN\
        );

    \I__1596\ : InMux
    port map (
            O => \N__7989\,
            I => \N__7986\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__7986\,
            I => \N__7982\
        );

    \I__1594\ : InMux
    port map (
            O => \N__7985\,
            I => \N__7979\
        );

    \I__1593\ : Odrv4
    port map (
            O => \N__7982\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__7979\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__7974\,
            I => \U712_REG_SM.N_373_cascade_\
        );

    \I__1590\ : InMux
    port map (
            O => \N__7971\,
            I => \N__7968\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__7968\,
            I => \U712_REG_SM.N_130\
        );

    \I__1588\ : CascadeMux
    port map (
            O => \N__7965\,
            I => \N__7962\
        );

    \I__1587\ : InMux
    port map (
            O => \N__7962\,
            I => \N__7958\
        );

    \I__1586\ : CascadeMux
    port map (
            O => \N__7961\,
            I => \N__7955\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__7958\,
            I => \N__7951\
        );

    \I__1584\ : InMux
    port map (
            O => \N__7955\,
            I => \N__7946\
        );

    \I__1583\ : InMux
    port map (
            O => \N__7954\,
            I => \N__7946\
        );

    \I__1582\ : Odrv4
    port map (
            O => \N__7951\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__7946\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1580\ : InMux
    port map (
            O => \N__7941\,
            I => \N__7935\
        );

    \I__1579\ : InMux
    port map (
            O => \N__7940\,
            I => \N__7935\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__7935\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__1577\ : CascadeMux
    port map (
            O => \N__7932\,
            I => \N__7929\
        );

    \I__1576\ : InMux
    port map (
            O => \N__7929\,
            I => \N__7926\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__7926\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\
        );

    \I__1574\ : CascadeMux
    port map (
            O => \N__7923\,
            I => \N__7920\
        );

    \I__1573\ : InMux
    port map (
            O => \N__7920\,
            I => \N__7917\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__7917\,
            I => \U712_REG_SM.N_406\
        );

    \I__1571\ : InMux
    port map (
            O => \N__7914\,
            I => \N__7910\
        );

    \I__1570\ : InMux
    port map (
            O => \N__7913\,
            I => \N__7907\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__7910\,
            I => \N__7899\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__7907\,
            I => \N__7899\
        );

    \I__1567\ : InMux
    port map (
            O => \N__7906\,
            I => \N__7896\
        );

    \I__1566\ : InMux
    port map (
            O => \N__7905\,
            I => \N__7893\
        );

    \I__1565\ : InMux
    port map (
            O => \N__7904\,
            I => \N__7890\
        );

    \I__1564\ : Span4Mux_v
    port map (
            O => \N__7899\,
            I => \N__7883\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__7896\,
            I => \N__7883\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__7893\,
            I => \N__7883\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__7890\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__7883\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1559\ : IoInMux
    port map (
            O => \N__7878\,
            I => \N__7875\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__7875\,
            I => \N__7872\
        );

    \I__1557\ : Span4Mux_s3_v
    port map (
            O => \N__7872\,
            I => \N__7869\
        );

    \I__1556\ : Span4Mux_v
    port map (
            O => \N__7869\,
            I => \N__7866\
        );

    \I__1555\ : Span4Mux_h
    port map (
            O => \N__7866\,
            I => \N__7863\
        );

    \I__1554\ : Span4Mux_h
    port map (
            O => \N__7863\,
            I => \N__7860\
        );

    \I__1553\ : Odrv4
    port map (
            O => \N__7860\,
            I => \CMA_c_10\
        );

    \I__1552\ : InMux
    port map (
            O => \N__7857\,
            I => \N__7854\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__7854\,
            I => \N__7851\
        );

    \I__1550\ : Span4Mux_h
    port map (
            O => \N__7851\,
            I => \N__7848\
        );

    \I__1549\ : Odrv4
    port map (
            O => \N__7848\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\
        );

    \I__1548\ : CascadeMux
    port map (
            O => \N__7845\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_\
        );

    \I__1547\ : IoInMux
    port map (
            O => \N__7842\,
            I => \N__7839\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__7839\,
            I => \N__7836\
        );

    \I__1545\ : Span12Mux_s5_v
    port map (
            O => \N__7836\,
            I => \N__7833\
        );

    \I__1544\ : Odrv12
    port map (
            O => \N__7833\,
            I => \CMA_c_2\
        );

    \I__1543\ : InMux
    port map (
            O => \N__7830\,
            I => \N__7827\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__7827\,
            I => \N__7824\
        );

    \I__1541\ : Odrv4
    port map (
            O => \N__7824\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__1540\ : IoInMux
    port map (
            O => \N__7821\,
            I => \N__7818\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__7818\,
            I => \N__7815\
        );

    \I__1538\ : IoSpan4Mux
    port map (
            O => \N__7815\,
            I => \N__7812\
        );

    \I__1537\ : Span4Mux_s3_h
    port map (
            O => \N__7812\,
            I => \N__7809\
        );

    \I__1536\ : Sp12to4
    port map (
            O => \N__7809\,
            I => \N__7806\
        );

    \I__1535\ : Span12Mux_h
    port map (
            O => \N__7806\,
            I => \N__7803\
        );

    \I__1534\ : Odrv12
    port map (
            O => \N__7803\,
            I => \CMA_c_4\
        );

    \I__1533\ : InMux
    port map (
            O => \N__7800\,
            I => \N__7793\
        );

    \I__1532\ : InMux
    port map (
            O => \N__7799\,
            I => \N__7793\
        );

    \I__1531\ : InMux
    port map (
            O => \N__7798\,
            I => \N__7790\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__7793\,
            I => \N__7783\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__7790\,
            I => \N__7780\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7789\,
            I => \N__7777\
        );

    \I__1527\ : InMux
    port map (
            O => \N__7788\,
            I => \N__7772\
        );

    \I__1526\ : InMux
    port map (
            O => \N__7787\,
            I => \N__7772\
        );

    \I__1525\ : InMux
    port map (
            O => \N__7786\,
            I => \N__7769\
        );

    \I__1524\ : Odrv4
    port map (
            O => \N__7783\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0\
        );

    \I__1523\ : Odrv12
    port map (
            O => \N__7780\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7777\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__7772\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__7769\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__7758\,
            I => \N__7750\
        );

    \I__1518\ : CascadeMux
    port map (
            O => \N__7757\,
            I => \N__7747\
        );

    \I__1517\ : CascadeMux
    port map (
            O => \N__7756\,
            I => \N__7744\
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__7755\,
            I => \N__7741\
        );

    \I__1515\ : CascadeMux
    port map (
            O => \N__7754\,
            I => \N__7737\
        );

    \I__1514\ : CascadeMux
    port map (
            O => \N__7753\,
            I => \N__7733\
        );

    \I__1513\ : InMux
    port map (
            O => \N__7750\,
            I => \N__7728\
        );

    \I__1512\ : InMux
    port map (
            O => \N__7747\,
            I => \N__7728\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7744\,
            I => \N__7725\
        );

    \I__1510\ : InMux
    port map (
            O => \N__7741\,
            I => \N__7722\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7740\,
            I => \N__7716\
        );

    \I__1508\ : InMux
    port map (
            O => \N__7737\,
            I => \N__7713\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7736\,
            I => \N__7708\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7733\,
            I => \N__7708\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__7728\,
            I => \N__7705\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__7725\,
            I => \N__7700\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7722\,
            I => \N__7700\
        );

    \I__1502\ : InMux
    port map (
            O => \N__7721\,
            I => \N__7695\
        );

    \I__1501\ : InMux
    port map (
            O => \N__7720\,
            I => \N__7695\
        );

    \I__1500\ : InMux
    port map (
            O => \N__7719\,
            I => \N__7692\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__7716\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__7713\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__7708\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__1496\ : Odrv4
    port map (
            O => \N__7705\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__1495\ : Odrv4
    port map (
            O => \N__7700\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__7695\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__7692\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7677\,
            I => \N__7674\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__7674\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__1490\ : IoInMux
    port map (
            O => \N__7671\,
            I => \N__7668\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__7668\,
            I => \N__7665\
        );

    \I__1488\ : Span12Mux_s5_h
    port map (
            O => \N__7665\,
            I => \N__7662\
        );

    \I__1487\ : Span12Mux_h
    port map (
            O => \N__7662\,
            I => \N__7659\
        );

    \I__1486\ : Odrv12
    port map (
            O => \N__7659\,
            I => \CMA_c_7\
        );

    \I__1485\ : CEMux
    port map (
            O => \N__7656\,
            I => \N__7651\
        );

    \I__1484\ : CEMux
    port map (
            O => \N__7655\,
            I => \N__7647\
        );

    \I__1483\ : CEMux
    port map (
            O => \N__7654\,
            I => \N__7644\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__7651\,
            I => \N__7640\
        );

    \I__1481\ : CEMux
    port map (
            O => \N__7650\,
            I => \N__7637\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__7647\,
            I => \N__7634\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7644\,
            I => \N__7631\
        );

    \I__1478\ : CEMux
    port map (
            O => \N__7643\,
            I => \N__7628\
        );

    \I__1477\ : Span4Mux_v
    port map (
            O => \N__7640\,
            I => \N__7625\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__7637\,
            I => \N__7622\
        );

    \I__1475\ : Span4Mux_v
    port map (
            O => \N__7634\,
            I => \N__7619\
        );

    \I__1474\ : Span4Mux_v
    port map (
            O => \N__7631\,
            I => \N__7616\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__7628\,
            I => \N__7609\
        );

    \I__1472\ : Span4Mux_v
    port map (
            O => \N__7625\,
            I => \N__7609\
        );

    \I__1471\ : Span4Mux_h
    port map (
            O => \N__7622\,
            I => \N__7609\
        );

    \I__1470\ : Odrv4
    port map (
            O => \N__7619\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__1469\ : Odrv4
    port map (
            O => \N__7616\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__1468\ : Odrv4
    port map (
            O => \N__7609\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7602\,
            I => \N__7599\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7599\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7596\,
            I => \N__7593\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__7593\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__1463\ : InMux
    port map (
            O => \N__7590\,
            I => \N__7587\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__7587\,
            I => \N__7584\
        );

    \I__1461\ : Span4Mux_h
    port map (
            O => \N__7584\,
            I => \N__7581\
        );

    \I__1460\ : Span4Mux_v
    port map (
            O => \N__7581\,
            I => \N__7578\
        );

    \I__1459\ : Sp12to4
    port map (
            O => \N__7578\,
            I => \N__7575\
        );

    \I__1458\ : Span12Mux_h
    port map (
            O => \N__7575\,
            I => \N__7572\
        );

    \I__1457\ : Odrv12
    port map (
            O => \N__7572\,
            I => \A_c_6\
        );

    \I__1456\ : InMux
    port map (
            O => \N__7569\,
            I => \N__7566\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__7566\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\
        );

    \I__1454\ : CEMux
    port map (
            O => \N__7563\,
            I => \N__7560\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__7560\,
            I => \N__7555\
        );

    \I__1452\ : CEMux
    port map (
            O => \N__7559\,
            I => \N__7552\
        );

    \I__1451\ : CEMux
    port map (
            O => \N__7558\,
            I => \N__7548\
        );

    \I__1450\ : Span4Mux_h
    port map (
            O => \N__7555\,
            I => \N__7543\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__7552\,
            I => \N__7543\
        );

    \I__1448\ : CEMux
    port map (
            O => \N__7551\,
            I => \N__7540\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__7548\,
            I => \N__7537\
        );

    \I__1446\ : Span4Mux_v
    port map (
            O => \N__7543\,
            I => \N__7534\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__7540\,
            I => \N__7531\
        );

    \I__1444\ : Odrv12
    port map (
            O => \N__7537\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\
        );

    \I__1443\ : Odrv4
    port map (
            O => \N__7534\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__7531\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\
        );

    \I__1441\ : InMux
    port map (
            O => \N__7524\,
            I => \N__7520\
        );

    \I__1440\ : InMux
    port map (
            O => \N__7523\,
            I => \N__7517\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__7520\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__7517\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1437\ : InMux
    port map (
            O => \N__7512\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__1436\ : InMux
    port map (
            O => \N__7509\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7506\,
            I => \N__7502\
        );

    \I__1434\ : InMux
    port map (
            O => \N__7505\,
            I => \N__7499\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__7502\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__7499\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1431\ : ClkMux
    port map (
            O => \N__7494\,
            I => \N__7467\
        );

    \I__1430\ : ClkMux
    port map (
            O => \N__7493\,
            I => \N__7467\
        );

    \I__1429\ : ClkMux
    port map (
            O => \N__7492\,
            I => \N__7467\
        );

    \I__1428\ : ClkMux
    port map (
            O => \N__7491\,
            I => \N__7467\
        );

    \I__1427\ : ClkMux
    port map (
            O => \N__7490\,
            I => \N__7467\
        );

    \I__1426\ : ClkMux
    port map (
            O => \N__7489\,
            I => \N__7467\
        );

    \I__1425\ : ClkMux
    port map (
            O => \N__7488\,
            I => \N__7467\
        );

    \I__1424\ : ClkMux
    port map (
            O => \N__7487\,
            I => \N__7467\
        );

    \I__1423\ : ClkMux
    port map (
            O => \N__7486\,
            I => \N__7467\
        );

    \I__1422\ : GlobalMux
    port map (
            O => \N__7467\,
            I => \N__7464\
        );

    \I__1421\ : gio2CtrlBuf
    port map (
            O => \N__7464\,
            I => \C1_c_g\
        );

    \I__1420\ : SRMux
    port map (
            O => \N__7461\,
            I => \N__7458\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__7458\,
            I => \N__7455\
        );

    \I__1418\ : Odrv12
    port map (
            O => \N__7455\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1417\ : InMux
    port map (
            O => \N__7452\,
            I => \N__7449\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__7449\,
            I => \N__7445\
        );

    \I__1415\ : InMux
    port map (
            O => \N__7448\,
            I => \N__7442\
        );

    \I__1414\ : Span4Mux_h
    port map (
            O => \N__7445\,
            I => \N__7435\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__7442\,
            I => \N__7435\
        );

    \I__1412\ : InMux
    port map (
            O => \N__7441\,
            I => \N__7432\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7440\,
            I => \N__7429\
        );

    \I__1410\ : Odrv4
    port map (
            O => \N__7435\,
            I => \DMA_CYCLEm\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__7432\,
            I => \DMA_CYCLEm\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__7429\,
            I => \DMA_CYCLEm\
        );

    \I__1407\ : IoInMux
    port map (
            O => \N__7422\,
            I => \N__7419\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__7419\,
            I => \N__7416\
        );

    \I__1405\ : Sp12to4
    port map (
            O => \N__7416\,
            I => \N__7411\
        );

    \I__1404\ : InMux
    port map (
            O => \N__7415\,
            I => \N__7408\
        );

    \I__1403\ : InMux
    port map (
            O => \N__7414\,
            I => \N__7405\
        );

    \I__1402\ : Span12Mux_v
    port map (
            O => \N__7411\,
            I => \N__7401\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__7408\,
            I => \N__7396\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__7405\,
            I => \N__7396\
        );

    \I__1399\ : InMux
    port map (
            O => \N__7404\,
            I => \N__7393\
        );

    \I__1398\ : Odrv12
    port map (
            O => \N__7401\,
            I => \DBENn_c\
        );

    \I__1397\ : Odrv4
    port map (
            O => \N__7396\,
            I => \DBENn_c\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__7393\,
            I => \DBENn_c\
        );

    \I__1395\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7383\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__7383\,
            I => \N__7380\
        );

    \I__1393\ : Odrv12
    port map (
            O => \N__7380\,
            I => \U712_REG_SM.N_402\
        );

    \I__1392\ : InMux
    port map (
            O => \N__7377\,
            I => \N__7373\
        );

    \I__1391\ : InMux
    port map (
            O => \N__7376\,
            I => \N__7370\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__7373\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__7370\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__1388\ : IoInMux
    port map (
            O => \N__7365\,
            I => \N__7361\
        );

    \I__1387\ : InMux
    port map (
            O => \N__7364\,
            I => \N__7358\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__7361\,
            I => \N__7355\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__7358\,
            I => \N__7352\
        );

    \I__1384\ : Span4Mux_s2_v
    port map (
            O => \N__7355\,
            I => \N__7349\
        );

    \I__1383\ : Span4Mux_v
    port map (
            O => \N__7352\,
            I => \N__7346\
        );

    \I__1382\ : Span4Mux_h
    port map (
            O => \N__7349\,
            I => \N__7343\
        );

    \I__1381\ : Span4Mux_v
    port map (
            O => \N__7346\,
            I => \N__7340\
        );

    \I__1380\ : Odrv4
    port map (
            O => \N__7343\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1379\ : Odrv4
    port map (
            O => \N__7340\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1378\ : IoInMux
    port map (
            O => \N__7335\,
            I => \N__7332\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__7332\,
            I => \N__7329\
        );

    \I__1376\ : Span4Mux_s2_v
    port map (
            O => \N__7329\,
            I => \N__7326\
        );

    \I__1375\ : Span4Mux_v
    port map (
            O => \N__7326\,
            I => \N__7323\
        );

    \I__1374\ : Span4Mux_h
    port map (
            O => \N__7323\,
            I => \N__7320\
        );

    \I__1373\ : Span4Mux_h
    port map (
            O => \N__7320\,
            I => \N__7317\
        );

    \I__1372\ : Odrv4
    port map (
            O => \N__7317\,
            I => \CRCSn_c\
        );

    \I__1371\ : InMux
    port map (
            O => \N__7314\,
            I => \N__7311\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__7311\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__1369\ : IoInMux
    port map (
            O => \N__7308\,
            I => \N__7305\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__7305\,
            I => \N__7302\
        );

    \I__1367\ : Span4Mux_s0_v
    port map (
            O => \N__7302\,
            I => \N__7299\
        );

    \I__1366\ : Sp12to4
    port map (
            O => \N__7299\,
            I => \N__7296\
        );

    \I__1365\ : Span12Mux_h
    port map (
            O => \N__7296\,
            I => \N__7293\
        );

    \I__1364\ : Odrv12
    port map (
            O => \N__7293\,
            I => \CMA_c_0\
        );

    \I__1363\ : IoInMux
    port map (
            O => \N__7290\,
            I => \N__7286\
        );

    \I__1362\ : IoInMux
    port map (
            O => \N__7289\,
            I => \N__7282\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__7286\,
            I => \N__7279\
        );

    \I__1360\ : IoInMux
    port map (
            O => \N__7285\,
            I => \N__7276\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__7282\,
            I => \N__7273\
        );

    \I__1358\ : Span4Mux_s1_v
    port map (
            O => \N__7279\,
            I => \N__7270\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7276\,
            I => \N__7267\
        );

    \I__1356\ : IoSpan4Mux
    port map (
            O => \N__7273\,
            I => \N__7264\
        );

    \I__1355\ : Sp12to4
    port map (
            O => \N__7270\,
            I => \N__7261\
        );

    \I__1354\ : Span4Mux_s2_h
    port map (
            O => \N__7267\,
            I => \N__7258\
        );

    \I__1353\ : Span4Mux_s0_v
    port map (
            O => \N__7264\,
            I => \N__7255\
        );

    \I__1352\ : Span12Mux_h
    port map (
            O => \N__7261\,
            I => \N__7252\
        );

    \I__1351\ : Sp12to4
    port map (
            O => \N__7258\,
            I => \N__7249\
        );

    \I__1350\ : Sp12to4
    port map (
            O => \N__7255\,
            I => \N__7246\
        );

    \I__1349\ : Span12Mux_v
    port map (
            O => \N__7252\,
            I => \N__7238\
        );

    \I__1348\ : Span12Mux_v
    port map (
            O => \N__7249\,
            I => \N__7238\
        );

    \I__1347\ : Span12Mux_v
    port map (
            O => \N__7246\,
            I => \N__7238\
        );

    \I__1346\ : InMux
    port map (
            O => \N__7245\,
            I => \N__7235\
        );

    \I__1345\ : Odrv12
    port map (
            O => \N__7238\,
            I => \TACK_OUTn\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__7235\,
            I => \TACK_OUTn\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7230\,
            I => \N__7227\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__7227\,
            I => \N__7224\
        );

    \I__1341\ : Odrv12
    port map (
            O => \N__7224\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\
        );

    \I__1340\ : InMux
    port map (
            O => \N__7221\,
            I => \N__7218\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__7218\,
            I => \N__7215\
        );

    \I__1338\ : Odrv4
    port map (
            O => \N__7215\,
            I => \U712_CHIP_RAM.N_367\
        );

    \I__1337\ : InMux
    port map (
            O => \N__7212\,
            I => \N__7209\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__7209\,
            I => \N__7206\
        );

    \I__1335\ : Span4Mux_v
    port map (
            O => \N__7206\,
            I => \N__7203\
        );

    \I__1334\ : Odrv4
    port map (
            O => \N__7203\,
            I => \U712_CHIP_RAM.N_419\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__7200\,
            I => \N__7197\
        );

    \I__1332\ : InMux
    port map (
            O => \N__7197\,
            I => \N__7193\
        );

    \I__1331\ : InMux
    port map (
            O => \N__7196\,
            I => \N__7189\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__7193\,
            I => \N__7186\
        );

    \I__1329\ : InMux
    port map (
            O => \N__7192\,
            I => \N__7183\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__7189\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1327\ : Odrv4
    port map (
            O => \N__7186\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__7183\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1325\ : InMux
    port map (
            O => \N__7176\,
            I => \N__7173\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__7173\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__1323\ : InMux
    port map (
            O => \N__7170\,
            I => \bfn_10_10_0_\
        );

    \I__1322\ : InMux
    port map (
            O => \N__7167\,
            I => \N__7163\
        );

    \I__1321\ : InMux
    port map (
            O => \N__7166\,
            I => \N__7160\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__7163\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__7160\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__1318\ : InMux
    port map (
            O => \N__7155\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__1317\ : InMux
    port map (
            O => \N__7152\,
            I => \N__7148\
        );

    \I__1316\ : InMux
    port map (
            O => \N__7151\,
            I => \N__7145\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__7148\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__7145\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__1313\ : InMux
    port map (
            O => \N__7140\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__1312\ : InMux
    port map (
            O => \N__7137\,
            I => \N__7133\
        );

    \I__1311\ : InMux
    port map (
            O => \N__7136\,
            I => \N__7130\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__7133\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__7130\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1308\ : InMux
    port map (
            O => \N__7125\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__1307\ : CascadeMux
    port map (
            O => \N__7122\,
            I => \N__7118\
        );

    \I__1306\ : InMux
    port map (
            O => \N__7121\,
            I => \N__7115\
        );

    \I__1305\ : InMux
    port map (
            O => \N__7118\,
            I => \N__7112\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__7115\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__7112\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1302\ : InMux
    port map (
            O => \N__7107\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__1301\ : InMux
    port map (
            O => \N__7104\,
            I => \N__7100\
        );

    \I__1300\ : InMux
    port map (
            O => \N__7103\,
            I => \N__7097\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__7100\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__7097\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1297\ : InMux
    port map (
            O => \N__7092\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__1296\ : InMux
    port map (
            O => \N__7089\,
            I => \N__7086\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__7086\,
            I => \N__7083\
        );

    \I__1294\ : Span4Mux_v
    port map (
            O => \N__7083\,
            I => \N__7080\
        );

    \I__1293\ : Span4Mux_v
    port map (
            O => \N__7080\,
            I => \N__7077\
        );

    \I__1292\ : Sp12to4
    port map (
            O => \N__7077\,
            I => \N__7074\
        );

    \I__1291\ : Span12Mux_h
    port map (
            O => \N__7074\,
            I => \N__7071\
        );

    \I__1290\ : Odrv12
    port map (
            O => \N__7071\,
            I => \A_c_15\
        );

    \I__1289\ : InMux
    port map (
            O => \N__7068\,
            I => \N__7065\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__7065\,
            I => \N__7062\
        );

    \I__1287\ : Span4Mux_v
    port map (
            O => \N__7062\,
            I => \N__7059\
        );

    \I__1286\ : Odrv4
    port map (
            O => \N__7059\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__7056\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\
        );

    \I__1284\ : InMux
    port map (
            O => \N__7053\,
            I => \N__7050\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__7050\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__1282\ : InMux
    port map (
            O => \N__7047\,
            I => \N__7044\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__7044\,
            I => \N__7041\
        );

    \I__1280\ : Span12Mux_v
    port map (
            O => \N__7041\,
            I => \N__7038\
        );

    \I__1279\ : Span12Mux_h
    port map (
            O => \N__7038\,
            I => \N__7035\
        );

    \I__1278\ : Odrv12
    port map (
            O => \N__7035\,
            I => \A_c_20\
        );

    \I__1277\ : InMux
    port map (
            O => \N__7032\,
            I => \N__7028\
        );

    \I__1276\ : InMux
    port map (
            O => \N__7031\,
            I => \N__7025\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__7028\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__7025\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__1273\ : InMux
    port map (
            O => \N__7020\,
            I => \N__7014\
        );

    \I__1272\ : InMux
    port map (
            O => \N__7019\,
            I => \N__7014\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__7014\,
            I => \N__7011\
        );

    \I__1270\ : Odrv4
    port map (
            O => \N__7011\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__1269\ : InMux
    port map (
            O => \N__7008\,
            I => \N__7005\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__7005\,
            I => \U712_CHIP_RAM.N_435\
        );

    \I__1267\ : InMux
    port map (
            O => \N__7002\,
            I => \N__6999\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__6999\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0\
        );

    \I__1265\ : CascadeMux
    port map (
            O => \N__6996\,
            I => \N__6992\
        );

    \I__1264\ : CascadeMux
    port map (
            O => \N__6995\,
            I => \N__6989\
        );

    \I__1263\ : InMux
    port map (
            O => \N__6992\,
            I => \N__6983\
        );

    \I__1262\ : InMux
    port map (
            O => \N__6989\,
            I => \N__6980\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__6988\,
            I => \N__6976\
        );

    \I__1260\ : CascadeMux
    port map (
            O => \N__6987\,
            I => \N__6973\
        );

    \I__1259\ : CascadeMux
    port map (
            O => \N__6986\,
            I => \N__6970\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__6983\,
            I => \N__6967\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__6980\,
            I => \N__6964\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6979\,
            I => \N__6957\
        );

    \I__1255\ : InMux
    port map (
            O => \N__6976\,
            I => \N__6957\
        );

    \I__1254\ : InMux
    port map (
            O => \N__6973\,
            I => \N__6957\
        );

    \I__1253\ : InMux
    port map (
            O => \N__6970\,
            I => \N__6954\
        );

    \I__1252\ : Odrv4
    port map (
            O => \N__6967\,
            I => \U712_CHIP_RAM.N_467\
        );

    \I__1251\ : Odrv4
    port map (
            O => \N__6964\,
            I => \U712_CHIP_RAM.N_467\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__6957\,
            I => \U712_CHIP_RAM.N_467\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__6954\,
            I => \U712_CHIP_RAM.N_467\
        );

    \I__1248\ : InMux
    port map (
            O => \N__6945\,
            I => \N__6942\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__6942\,
            I => \N__6939\
        );

    \I__1246\ : Span4Mux_h
    port map (
            O => \N__6939\,
            I => \N__6936\
        );

    \I__1245\ : Odrv4
    port map (
            O => \N__6936\,
            I => \U712_CHIP_RAM.DBENn_7_0_0\
        );

    \I__1244\ : InMux
    port map (
            O => \N__6933\,
            I => \N__6929\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6932\,
            I => \N__6926\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__6929\,
            I => \N__6922\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__6926\,
            I => \N__6919\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6925\,
            I => \N__6916\
        );

    \I__1239\ : Span4Mux_v
    port map (
            O => \N__6922\,
            I => \N__6913\
        );

    \I__1238\ : Span4Mux_v
    port map (
            O => \N__6919\,
            I => \N__6910\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__6916\,
            I => \N__6907\
        );

    \I__1236\ : Sp12to4
    port map (
            O => \N__6913\,
            I => \N__6902\
        );

    \I__1235\ : Sp12to4
    port map (
            O => \N__6910\,
            I => \N__6902\
        );

    \I__1234\ : Span12Mux_h
    port map (
            O => \N__6907\,
            I => \N__6899\
        );

    \I__1233\ : Span12Mux_h
    port map (
            O => \N__6902\,
            I => \N__6896\
        );

    \I__1232\ : Span12Mux_v
    port map (
            O => \N__6899\,
            I => \N__6893\
        );

    \I__1231\ : Span12Mux_v
    port map (
            O => \N__6896\,
            I => \N__6890\
        );

    \I__1230\ : Odrv12
    port map (
            O => \N__6893\,
            I => \AWEn_c\
        );

    \I__1229\ : Odrv12
    port map (
            O => \N__6890\,
            I => \AWEn_c\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6885\,
            I => \N__6880\
        );

    \I__1227\ : InMux
    port map (
            O => \N__6884\,
            I => \N__6877\
        );

    \I__1226\ : InMux
    port map (
            O => \N__6883\,
            I => \N__6874\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__6880\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__6877\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__6874\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__1222\ : IoInMux
    port map (
            O => \N__6867\,
            I => \N__6864\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__6864\,
            I => \N__6861\
        );

    \I__1220\ : IoSpan4Mux
    port map (
            O => \N__6861\,
            I => \N__6858\
        );

    \I__1219\ : Sp12to4
    port map (
            O => \N__6858\,
            I => \N__6855\
        );

    \I__1218\ : Span12Mux_s7_v
    port map (
            O => \N__6855\,
            I => \N__6851\
        );

    \I__1217\ : InMux
    port map (
            O => \N__6854\,
            I => \N__6848\
        );

    \I__1216\ : Odrv12
    port map (
            O => \N__6851\,
            I => \DBDIR_c\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__6848\,
            I => \DBDIR_c\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6843\,
            I => \N__6840\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__6840\,
            I => \U712_CHIP_RAM.N_361\
        );

    \I__1212\ : IoInMux
    port map (
            O => \N__6837\,
            I => \N__6834\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__6834\,
            I => \N__6831\
        );

    \I__1210\ : Span4Mux_s3_h
    port map (
            O => \N__6831\,
            I => \N__6828\
        );

    \I__1209\ : Span4Mux_v
    port map (
            O => \N__6828\,
            I => \N__6825\
        );

    \I__1208\ : Span4Mux_v
    port map (
            O => \N__6825\,
            I => \N__6822\
        );

    \I__1207\ : Sp12to4
    port map (
            O => \N__6822\,
            I => \N__6819\
        );

    \I__1206\ : Span12Mux_s10_h
    port map (
            O => \N__6819\,
            I => \N__6816\
        );

    \I__1205\ : Odrv12
    port map (
            O => \N__6816\,
            I => \CMA_c_5\
        );

    \I__1204\ : IoInMux
    port map (
            O => \N__6813\,
            I => \N__6810\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__6810\,
            I => \N__6807\
        );

    \I__1202\ : Span4Mux_s0_v
    port map (
            O => \N__6807\,
            I => \N__6804\
        );

    \I__1201\ : Span4Mux_v
    port map (
            O => \N__6804\,
            I => \N__6801\
        );

    \I__1200\ : Span4Mux_v
    port map (
            O => \N__6801\,
            I => \N__6798\
        );

    \I__1199\ : Sp12to4
    port map (
            O => \N__6798\,
            I => \N__6794\
        );

    \I__1198\ : InMux
    port map (
            O => \N__6797\,
            I => \N__6791\
        );

    \I__1197\ : Span12Mux_h
    port map (
            O => \N__6794\,
            I => \N__6788\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__6791\,
            I => \N__6785\
        );

    \I__1195\ : Span12Mux_v
    port map (
            O => \N__6788\,
            I => \N__6780\
        );

    \I__1194\ : Span12Mux_h
    port map (
            O => \N__6785\,
            I => \N__6780\
        );

    \I__1193\ : Odrv12
    port map (
            O => \N__6780\,
            I => \A_c_10\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6777\,
            I => \N__6774\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__6774\,
            I => \N__6771\
        );

    \I__1190\ : Span4Mux_h
    port map (
            O => \N__6771\,
            I => \N__6768\
        );

    \I__1189\ : Odrv4
    port map (
            O => \N__6768\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\
        );

    \I__1188\ : CascadeMux
    port map (
            O => \N__6765\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6762\,
            I => \N__6759\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__6759\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__1185\ : CascadeMux
    port map (
            O => \N__6756\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_\
        );

    \I__1184\ : InMux
    port map (
            O => \N__6753\,
            I => \N__6750\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__6750\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__1182\ : IoInMux
    port map (
            O => \N__6747\,
            I => \N__6744\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__6744\,
            I => \N__6741\
        );

    \I__1180\ : Span4Mux_s3_v
    port map (
            O => \N__6741\,
            I => \N__6738\
        );

    \I__1179\ : Span4Mux_v
    port map (
            O => \N__6738\,
            I => \N__6735\
        );

    \I__1178\ : Span4Mux_v
    port map (
            O => \N__6735\,
            I => \N__6732\
        );

    \I__1177\ : Odrv4
    port map (
            O => \N__6732\,
            I => \CMA_c_1\
        );

    \I__1176\ : InMux
    port map (
            O => \N__6729\,
            I => \N__6726\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6726\,
            I => \N__6723\
        );

    \I__1174\ : Odrv4
    port map (
            O => \N__6723\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6720\,
            I => \N__6717\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__6717\,
            I => \N__6714\
        );

    \I__1171\ : Span4Mux_v
    port map (
            O => \N__6714\,
            I => \N__6711\
        );

    \I__1170\ : Sp12to4
    port map (
            O => \N__6711\,
            I => \N__6708\
        );

    \I__1169\ : Span12Mux_h
    port map (
            O => \N__6708\,
            I => \N__6705\
        );

    \I__1168\ : Odrv12
    port map (
            O => \N__6705\,
            I => \A_c_13\
        );

    \I__1167\ : InMux
    port map (
            O => \N__6702\,
            I => \N__6699\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6699\,
            I => \N__6696\
        );

    \I__1165\ : Span4Mux_h
    port map (
            O => \N__6696\,
            I => \N__6693\
        );

    \I__1164\ : Sp12to4
    port map (
            O => \N__6693\,
            I => \N__6690\
        );

    \I__1163\ : Span12Mux_v
    port map (
            O => \N__6690\,
            I => \N__6687\
        );

    \I__1162\ : Odrv12
    port map (
            O => \N__6687\,
            I => \A_c_17\
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__6684\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6681\,
            I => \N__6678\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__6678\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\
        );

    \I__1158\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6672\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__6672\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1156\ : IoInMux
    port map (
            O => \N__6669\,
            I => \N__6666\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__6666\,
            I => \N__6663\
        );

    \I__1154\ : Span4Mux_s0_h
    port map (
            O => \N__6663\,
            I => \N__6660\
        );

    \I__1153\ : Sp12to4
    port map (
            O => \N__6660\,
            I => \N__6657\
        );

    \I__1152\ : Span12Mux_s9_v
    port map (
            O => \N__6657\,
            I => \N__6654\
        );

    \I__1151\ : Span12Mux_h
    port map (
            O => \N__6654\,
            I => \N__6651\
        );

    \I__1150\ : Odrv12
    port map (
            O => \N__6651\,
            I => \CMA_c_3\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6648\,
            I => \N__6645\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__6645\,
            I => \N__6642\
        );

    \I__1147\ : Span12Mux_v
    port map (
            O => \N__6642\,
            I => \N__6639\
        );

    \I__1146\ : Span12Mux_h
    port map (
            O => \N__6639\,
            I => \N__6636\
        );

    \I__1145\ : Odrv12
    port map (
            O => \N__6636\,
            I => \A_c_14\
        );

    \I__1144\ : InMux
    port map (
            O => \N__6633\,
            I => \N__6628\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__6632\,
            I => \N__6623\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6631\,
            I => \N__6620\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__6628\,
            I => \N__6617\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6627\,
            I => \N__6614\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6626\,
            I => \N__6609\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6623\,
            I => \N__6609\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__6620\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1136\ : Odrv4
    port map (
            O => \N__6617\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__6614\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__6609\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__6600\,
            I => \U712_CHIP_RAM.REFRESH_RST_cascade_\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6597\,
            I => \N__6593\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6596\,
            I => \N__6590\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__6593\,
            I => \N__6584\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6590\,
            I => \N__6581\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6589\,
            I => \N__6574\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6588\,
            I => \N__6574\
        );

    \I__1126\ : InMux
    port map (
            O => \N__6587\,
            I => \N__6574\
        );

    \I__1125\ : Odrv4
    port map (
            O => \N__6584\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1124\ : Odrv4
    port map (
            O => \N__6581\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6574\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1122\ : CascadeMux
    port map (
            O => \N__6567\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_cascade_\
        );

    \I__1121\ : InMux
    port map (
            O => \N__6564\,
            I => \N__6560\
        );

    \I__1120\ : IoInMux
    port map (
            O => \N__6563\,
            I => \N__6557\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__6560\,
            I => \N__6554\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6557\,
            I => \N__6551\
        );

    \I__1117\ : Span4Mux_v
    port map (
            O => \N__6554\,
            I => \N__6548\
        );

    \I__1116\ : Span12Mux_s4_v
    port map (
            O => \N__6551\,
            I => \N__6545\
        );

    \I__1115\ : Span4Mux_v
    port map (
            O => \N__6548\,
            I => \N__6542\
        );

    \I__1114\ : Span12Mux_v
    port map (
            O => \N__6545\,
            I => \N__6537\
        );

    \I__1113\ : Sp12to4
    port map (
            O => \N__6542\,
            I => \N__6537\
        );

    \I__1112\ : Span12Mux_h
    port map (
            O => \N__6537\,
            I => \N__6534\
        );

    \I__1111\ : Odrv12
    port map (
            O => \N__6534\,
            I => \A_c_9\
        );

    \I__1110\ : InMux
    port map (
            O => \N__6531\,
            I => \N__6528\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__6528\,
            I => \N__6525\
        );

    \I__1108\ : Span4Mux_h
    port map (
            O => \N__6525\,
            I => \N__6522\
        );

    \I__1107\ : Odrv4
    port map (
            O => \N__6522\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__6519\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\
        );

    \I__1105\ : InMux
    port map (
            O => \N__6516\,
            I => \N__6513\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__6513\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1103\ : InMux
    port map (
            O => \N__6510\,
            I => \N__6507\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__6507\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__1101\ : CascadeMux
    port map (
            O => \N__6504\,
            I => \U712_CHIP_RAM.N_335_cascade_\
        );

    \I__1100\ : IoInMux
    port map (
            O => \N__6501\,
            I => \N__6498\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__6498\,
            I => \N__6495\
        );

    \I__1098\ : Span12Mux_s7_v
    port map (
            O => \N__6495\,
            I => \N__6492\
        );

    \I__1097\ : Span12Mux_v
    port map (
            O => \N__6492\,
            I => \N__6489\
        );

    \I__1096\ : Odrv12
    port map (
            O => \N__6489\,
            I => \N_202_i\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6486\,
            I => \N__6483\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6483\,
            I => \N__6479\
        );

    \I__1093\ : InMux
    port map (
            O => \N__6482\,
            I => \N__6476\
        );

    \I__1092\ : Span4Mux_h
    port map (
            O => \N__6479\,
            I => \N__6471\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__6476\,
            I => \N__6471\
        );

    \I__1090\ : Span4Mux_v
    port map (
            O => \N__6471\,
            I => \N__6468\
        );

    \I__1089\ : Sp12to4
    port map (
            O => \N__6468\,
            I => \N__6465\
        );

    \I__1088\ : Span12Mux_h
    port map (
            O => \N__6465\,
            I => \N__6462\
        );

    \I__1087\ : Odrv12
    port map (
            O => \N__6462\,
            I => \TSn_c\
        );

    \I__1086\ : InMux
    port map (
            O => \N__6459\,
            I => \N__6456\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__6456\,
            I => \N__6453\
        );

    \I__1084\ : Span4Mux_h
    port map (
            O => \N__6453\,
            I => \N__6450\
        );

    \I__1083\ : Span4Mux_v
    port map (
            O => \N__6450\,
            I => \N__6447\
        );

    \I__1082\ : Span4Mux_v
    port map (
            O => \N__6447\,
            I => \N__6444\
        );

    \I__1081\ : Odrv4
    port map (
            O => \N__6444\,
            I => \RAMSPACEn_c\
        );

    \I__1080\ : IoInMux
    port map (
            O => \N__6441\,
            I => \N__6438\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__6438\,
            I => \N__6435\
        );

    \I__1078\ : IoSpan4Mux
    port map (
            O => \N__6435\,
            I => \N__6432\
        );

    \I__1077\ : Span4Mux_s3_v
    port map (
            O => \N__6432\,
            I => \N__6429\
        );

    \I__1076\ : Span4Mux_v
    port map (
            O => \N__6429\,
            I => \N__6426\
        );

    \I__1075\ : Odrv4
    port map (
            O => \N__6426\,
            I => \N_165_i\
        );

    \I__1074\ : IoInMux
    port map (
            O => \N__6423\,
            I => \N__6420\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__6420\,
            I => \N__6417\
        );

    \I__1072\ : Span4Mux_s2_h
    port map (
            O => \N__6417\,
            I => \N__6414\
        );

    \I__1071\ : Span4Mux_v
    port map (
            O => \N__6414\,
            I => \N__6411\
        );

    \I__1070\ : Span4Mux_h
    port map (
            O => \N__6411\,
            I => \N__6408\
        );

    \I__1069\ : Sp12to4
    port map (
            O => \N__6408\,
            I => \N__6405\
        );

    \I__1068\ : Span12Mux_h
    port map (
            O => \N__6405\,
            I => \N__6402\
        );

    \I__1067\ : Odrv12
    port map (
            O => \N__6402\,
            I => \WEn_c\
        );

    \I__1066\ : IoInMux
    port map (
            O => \N__6399\,
            I => \N__6396\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__6396\,
            I => \N__6393\
        );

    \I__1064\ : Span4Mux_s0_v
    port map (
            O => \N__6393\,
            I => \N__6390\
        );

    \I__1063\ : Sp12to4
    port map (
            O => \N__6390\,
            I => \N__6387\
        );

    \I__1062\ : Span12Mux_h
    port map (
            O => \N__6387\,
            I => \N__6384\
        );

    \I__1061\ : Odrv12
    port map (
            O => \N__6384\,
            I => \RASn_c\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__6381\,
            I => \U712_CHIP_RAM.N_428_cascade_\
        );

    \I__1059\ : InMux
    port map (
            O => \N__6378\,
            I => \N__6373\
        );

    \I__1058\ : InMux
    port map (
            O => \N__6377\,
            I => \N__6368\
        );

    \I__1057\ : InMux
    port map (
            O => \N__6376\,
            I => \N__6368\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__6373\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__6368\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\
        );

    \I__1054\ : SRMux
    port map (
            O => \N__6363\,
            I => \N__6359\
        );

    \I__1053\ : SRMux
    port map (
            O => \N__6362\,
            I => \N__6356\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6359\,
            I => \N__6353\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__6356\,
            I => \N__6350\
        );

    \I__1050\ : Odrv4
    port map (
            O => \N__6353\,
            I => \U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1\
        );

    \I__1049\ : Odrv4
    port map (
            O => \N__6350\,
            I => \U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1\
        );

    \I__1048\ : InMux
    port map (
            O => \N__6345\,
            I => \N__6342\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__6342\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6339\,
            I => \N__6333\
        );

    \I__1045\ : InMux
    port map (
            O => \N__6338\,
            I => \N__6333\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__6333\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\
        );

    \I__1043\ : InMux
    port map (
            O => \N__6330\,
            I => \N__6327\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__6327\,
            I => \U712_CHIP_RAM.N_430\
        );

    \I__1041\ : CascadeMux
    port map (
            O => \N__6324\,
            I => \U712_CHIP_RAM.REFRESH5lto7_0_cascade_\
        );

    \I__1040\ : InMux
    port map (
            O => \N__6321\,
            I => \N__6318\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__6318\,
            I => \U712_CHIP_RAM.REFRESH5lt7\
        );

    \I__1038\ : CascadeMux
    port map (
            O => \N__6315\,
            I => \N__6312\
        );

    \I__1037\ : InMux
    port map (
            O => \N__6312\,
            I => \N__6308\
        );

    \I__1036\ : CascadeMux
    port map (
            O => \N__6311\,
            I => \N__6304\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__6308\,
            I => \N__6301\
        );

    \I__1034\ : InMux
    port map (
            O => \N__6307\,
            I => \N__6296\
        );

    \I__1033\ : InMux
    port map (
            O => \N__6304\,
            I => \N__6296\
        );

    \I__1032\ : Odrv12
    port map (
            O => \N__6301\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__6296\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6291\,
            I => \N__6288\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6288\,
            I => \N__6283\
        );

    \I__1028\ : InMux
    port map (
            O => \N__6287\,
            I => \N__6278\
        );

    \I__1027\ : InMux
    port map (
            O => \N__6286\,
            I => \N__6278\
        );

    \I__1026\ : Odrv4
    port map (
            O => \N__6283\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__6278\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1024\ : CascadeMux
    port map (
            O => \N__6273\,
            I => \U712_CHIP_RAM.N_435_cascade_\
        );

    \I__1023\ : CascadeMux
    port map (
            O => \N__6270\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_cascade_\
        );

    \I__1022\ : CEMux
    port map (
            O => \N__6267\,
            I => \N__6264\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__6264\,
            I => \N__6261\
        );

    \I__1020\ : Odrv12
    port map (
            O => \N__6261\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_0\
        );

    \I__1019\ : InMux
    port map (
            O => \N__6258\,
            I => \N__6255\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__6255\,
            I => \N__6251\
        );

    \I__1017\ : InMux
    port map (
            O => \N__6254\,
            I => \N__6248\
        );

    \I__1016\ : Span4Mux_h
    port map (
            O => \N__6251\,
            I => \N__6245\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__6248\,
            I => \U712_CHIP_RAM.N_325\
        );

    \I__1014\ : Odrv4
    port map (
            O => \N__6245\,
            I => \U712_CHIP_RAM.N_325\
        );

    \I__1013\ : InMux
    port map (
            O => \N__6240\,
            I => \N__6236\
        );

    \I__1012\ : InMux
    port map (
            O => \N__6239\,
            I => \N__6233\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__6236\,
            I => \N__6230\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__6233\,
            I => \U712_CHIP_RAM.N_321\
        );

    \I__1009\ : Odrv4
    port map (
            O => \N__6230\,
            I => \U712_CHIP_RAM.N_321\
        );

    \I__1008\ : InMux
    port map (
            O => \N__6225\,
            I => \N__6217\
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__6224\,
            I => \N__6206\
        );

    \I__1006\ : CascadeMux
    port map (
            O => \N__6223\,
            I => \N__6203\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6222\,
            I => \N__6191\
        );

    \I__1004\ : InMux
    port map (
            O => \N__6221\,
            I => \N__6191\
        );

    \I__1003\ : InMux
    port map (
            O => \N__6220\,
            I => \N__6188\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__6217\,
            I => \N__6185\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6216\,
            I => \N__6182\
        );

    \I__1000\ : InMux
    port map (
            O => \N__6215\,
            I => \N__6173\
        );

    \I__999\ : InMux
    port map (
            O => \N__6214\,
            I => \N__6173\
        );

    \I__998\ : InMux
    port map (
            O => \N__6213\,
            I => \N__6173\
        );

    \I__997\ : InMux
    port map (
            O => \N__6212\,
            I => \N__6173\
        );

    \I__996\ : InMux
    port map (
            O => \N__6211\,
            I => \N__6168\
        );

    \I__995\ : InMux
    port map (
            O => \N__6210\,
            I => \N__6168\
        );

    \I__994\ : InMux
    port map (
            O => \N__6209\,
            I => \N__6160\
        );

    \I__993\ : InMux
    port map (
            O => \N__6206\,
            I => \N__6155\
        );

    \I__992\ : InMux
    port map (
            O => \N__6203\,
            I => \N__6155\
        );

    \I__991\ : InMux
    port map (
            O => \N__6202\,
            I => \N__6150\
        );

    \I__990\ : InMux
    port map (
            O => \N__6201\,
            I => \N__6150\
        );

    \I__989\ : InMux
    port map (
            O => \N__6200\,
            I => \N__6139\
        );

    \I__988\ : InMux
    port map (
            O => \N__6199\,
            I => \N__6139\
        );

    \I__987\ : InMux
    port map (
            O => \N__6198\,
            I => \N__6139\
        );

    \I__986\ : InMux
    port map (
            O => \N__6197\,
            I => \N__6139\
        );

    \I__985\ : InMux
    port map (
            O => \N__6196\,
            I => \N__6139\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__6191\,
            I => \N__6136\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__6188\,
            I => \N__6125\
        );

    \I__982\ : Span4Mux_v
    port map (
            O => \N__6185\,
            I => \N__6125\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__6182\,
            I => \N__6125\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__6173\,
            I => \N__6125\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__6168\,
            I => \N__6125\
        );

    \I__978\ : InMux
    port map (
            O => \N__6167\,
            I => \N__6114\
        );

    \I__977\ : InMux
    port map (
            O => \N__6166\,
            I => \N__6114\
        );

    \I__976\ : InMux
    port map (
            O => \N__6165\,
            I => \N__6114\
        );

    \I__975\ : InMux
    port map (
            O => \N__6164\,
            I => \N__6114\
        );

    \I__974\ : InMux
    port map (
            O => \N__6163\,
            I => \N__6114\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__6160\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__6155\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__6150\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__6139\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__969\ : Odrv4
    port map (
            O => \N__6136\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__968\ : Odrv4
    port map (
            O => \N__6125\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__6114\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__966\ : CascadeMux
    port map (
            O => \N__6099\,
            I => \N__6090\
        );

    \I__965\ : InMux
    port map (
            O => \N__6098\,
            I => \N__6085\
        );

    \I__964\ : CascadeMux
    port map (
            O => \N__6097\,
            I => \N__6082\
        );

    \I__963\ : CascadeMux
    port map (
            O => \N__6096\,
            I => \N__6078\
        );

    \I__962\ : CascadeMux
    port map (
            O => \N__6095\,
            I => \N__6074\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__6094\,
            I => \N__6071\
        );

    \I__960\ : CascadeMux
    port map (
            O => \N__6093\,
            I => \N__6066\
        );

    \I__959\ : InMux
    port map (
            O => \N__6090\,
            I => \N__6063\
        );

    \I__958\ : CascadeMux
    port map (
            O => \N__6089\,
            I => \N__6057\
        );

    \I__957\ : InMux
    port map (
            O => \N__6088\,
            I => \N__6054\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__6085\,
            I => \N__6051\
        );

    \I__955\ : InMux
    port map (
            O => \N__6082\,
            I => \N__6040\
        );

    \I__954\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6040\
        );

    \I__953\ : InMux
    port map (
            O => \N__6078\,
            I => \N__6040\
        );

    \I__952\ : InMux
    port map (
            O => \N__6077\,
            I => \N__6040\
        );

    \I__951\ : InMux
    port map (
            O => \N__6074\,
            I => \N__6031\
        );

    \I__950\ : InMux
    port map (
            O => \N__6071\,
            I => \N__6031\
        );

    \I__949\ : InMux
    port map (
            O => \N__6070\,
            I => \N__6031\
        );

    \I__948\ : InMux
    port map (
            O => \N__6069\,
            I => \N__6031\
        );

    \I__947\ : InMux
    port map (
            O => \N__6066\,
            I => \N__6018\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__6063\,
            I => \N__6015\
        );

    \I__945\ : InMux
    port map (
            O => \N__6062\,
            I => \N__6008\
        );

    \I__944\ : InMux
    port map (
            O => \N__6061\,
            I => \N__6008\
        );

    \I__943\ : InMux
    port map (
            O => \N__6060\,
            I => \N__6008\
        );

    \I__942\ : InMux
    port map (
            O => \N__6057\,
            I => \N__6005\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__6054\,
            I => \N__6000\
        );

    \I__940\ : Span4Mux_h
    port map (
            O => \N__6051\,
            I => \N__6000\
        );

    \I__939\ : InMux
    port map (
            O => \N__6050\,
            I => \N__5995\
        );

    \I__938\ : InMux
    port map (
            O => \N__6049\,
            I => \N__5995\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__6040\,
            I => \N__5990\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__6031\,
            I => \N__5990\
        );

    \I__935\ : InMux
    port map (
            O => \N__6030\,
            I => \N__5983\
        );

    \I__934\ : InMux
    port map (
            O => \N__6029\,
            I => \N__5983\
        );

    \I__933\ : InMux
    port map (
            O => \N__6028\,
            I => \N__5983\
        );

    \I__932\ : InMux
    port map (
            O => \N__6027\,
            I => \N__5976\
        );

    \I__931\ : InMux
    port map (
            O => \N__6026\,
            I => \N__5976\
        );

    \I__930\ : InMux
    port map (
            O => \N__6025\,
            I => \N__5976\
        );

    \I__929\ : InMux
    port map (
            O => \N__6024\,
            I => \N__5967\
        );

    \I__928\ : InMux
    port map (
            O => \N__6023\,
            I => \N__5967\
        );

    \I__927\ : InMux
    port map (
            O => \N__6022\,
            I => \N__5967\
        );

    \I__926\ : InMux
    port map (
            O => \N__6021\,
            I => \N__5967\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__6018\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__924\ : Odrv4
    port map (
            O => \N__6015\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__6008\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__6005\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__921\ : Odrv4
    port map (
            O => \N__6000\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__5995\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__919\ : Odrv4
    port map (
            O => \N__5990\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5983\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__5976\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__5967\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__915\ : InMux
    port map (
            O => \N__5946\,
            I => \N__5942\
        );

    \I__914\ : InMux
    port map (
            O => \N__5945\,
            I => \N__5938\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__5942\,
            I => \N__5935\
        );

    \I__912\ : InMux
    port map (
            O => \N__5941\,
            I => \N__5932\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__5938\,
            I => \U712_CHIP_RAM.N_551\
        );

    \I__910\ : Odrv4
    port map (
            O => \N__5935\,
            I => \U712_CHIP_RAM.N_551\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5932\,
            I => \U712_CHIP_RAM.N_551\
        );

    \I__908\ : CascadeMux
    port map (
            O => \N__5925\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_2_0_cascade_\
        );

    \I__907\ : InMux
    port map (
            O => \N__5922\,
            I => \N__5919\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__5919\,
            I => \N__5916\
        );

    \I__905\ : Span4Mux_h
    port map (
            O => \N__5916\,
            I => \N__5913\
        );

    \I__904\ : Odrv4
    port map (
            O => \N__5913\,
            I => \U712_CHIP_RAM.LATCH_CLK_6\
        );

    \I__903\ : IoInMux
    port map (
            O => \N__5910\,
            I => \N__5906\
        );

    \I__902\ : IoInMux
    port map (
            O => \N__5909\,
            I => \N__5903\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__5906\,
            I => \N__5898\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__5903\,
            I => \N__5898\
        );

    \I__899\ : IoSpan4Mux
    port map (
            O => \N__5898\,
            I => \N__5895\
        );

    \I__898\ : IoSpan4Mux
    port map (
            O => \N__5895\,
            I => \N__5892\
        );

    \I__897\ : Sp12to4
    port map (
            O => \N__5892\,
            I => \N__5889\
        );

    \I__896\ : Span12Mux_s6_v
    port map (
            O => \N__5889\,
            I => \N__5885\
        );

    \I__895\ : InMux
    port map (
            O => \N__5888\,
            I => \N__5882\
        );

    \I__894\ : Odrv12
    port map (
            O => \N__5885\,
            I => \RAMENn_c\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__5882\,
            I => \RAMENn_c\
        );

    \I__892\ : InMux
    port map (
            O => \N__5877\,
            I => \N__5873\
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__5876\,
            I => \N__5868\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__5873\,
            I => \N__5865\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__5872\,
            I => \N__5861\
        );

    \I__888\ : InMux
    port map (
            O => \N__5871\,
            I => \N__5854\
        );

    \I__887\ : InMux
    port map (
            O => \N__5868\,
            I => \N__5851\
        );

    \I__886\ : Span4Mux_v
    port map (
            O => \N__5865\,
            I => \N__5848\
        );

    \I__885\ : InMux
    port map (
            O => \N__5864\,
            I => \N__5843\
        );

    \I__884\ : InMux
    port map (
            O => \N__5861\,
            I => \N__5843\
        );

    \I__883\ : InMux
    port map (
            O => \N__5860\,
            I => \N__5836\
        );

    \I__882\ : InMux
    port map (
            O => \N__5859\,
            I => \N__5836\
        );

    \I__881\ : InMux
    port map (
            O => \N__5858\,
            I => \N__5836\
        );

    \I__880\ : InMux
    port map (
            O => \N__5857\,
            I => \N__5833\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__5854\,
            I => \N__5830\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__5851\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__877\ : Odrv4
    port map (
            O => \N__5848\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__5843\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5836\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__5833\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__873\ : Odrv4
    port map (
            O => \N__5830\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__872\ : InMux
    port map (
            O => \N__5817\,
            I => \N__5813\
        );

    \I__871\ : InMux
    port map (
            O => \N__5816\,
            I => \N__5810\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__5813\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__5810\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3\
        );

    \I__868\ : IoInMux
    port map (
            O => \N__5805\,
            I => \N__5802\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__5802\,
            I => \N__5799\
        );

    \I__866\ : IoSpan4Mux
    port map (
            O => \N__5799\,
            I => \N__5796\
        );

    \I__865\ : Span4Mux_s0_v
    port map (
            O => \N__5796\,
            I => \N__5793\
        );

    \I__864\ : Sp12to4
    port map (
            O => \N__5793\,
            I => \N__5789\
        );

    \I__863\ : InMux
    port map (
            O => \N__5792\,
            I => \N__5786\
        );

    \I__862\ : Span12Mux_s8_v
    port map (
            O => \N__5789\,
            I => \N__5783\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__5786\,
            I => \N__5780\
        );

    \I__860\ : Span12Mux_v
    port map (
            O => \N__5783\,
            I => \N__5777\
        );

    \I__859\ : Span4Mux_v
    port map (
            O => \N__5780\,
            I => \N__5774\
        );

    \I__858\ : Span12Mux_h
    port map (
            O => \N__5777\,
            I => \N__5769\
        );

    \I__857\ : Sp12to4
    port map (
            O => \N__5774\,
            I => \N__5769\
        );

    \I__856\ : Odrv12
    port map (
            O => \N__5769\,
            I => \A_c_11\
        );

    \I__855\ : InMux
    port map (
            O => \N__5766\,
            I => \N__5763\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__5763\,
            I => \N__5760\
        );

    \I__853\ : Odrv4
    port map (
            O => \N__5760\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\
        );

    \I__852\ : InMux
    port map (
            O => \N__5757\,
            I => \N__5753\
        );

    \I__851\ : InMux
    port map (
            O => \N__5756\,
            I => \N__5750\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__5753\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_6\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__5750\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_6\
        );

    \I__848\ : InMux
    port map (
            O => \N__5745\,
            I => \N__5742\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__5742\,
            I => \U712_CHIP_RAM.m93_i_a2_5\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__5739\,
            I => \N__5736\
        );

    \I__845\ : InMux
    port map (
            O => \N__5736\,
            I => \N__5733\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__5733\,
            I => \N__5727\
        );

    \I__843\ : CascadeMux
    port map (
            O => \N__5732\,
            I => \N__5724\
        );

    \I__842\ : InMux
    port map (
            O => \N__5731\,
            I => \N__5719\
        );

    \I__841\ : InMux
    port map (
            O => \N__5730\,
            I => \N__5719\
        );

    \I__840\ : Span4Mux_h
    port map (
            O => \N__5727\,
            I => \N__5716\
        );

    \I__839\ : InMux
    port map (
            O => \N__5724\,
            I => \N__5713\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__5719\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_0\
        );

    \I__837\ : Odrv4
    port map (
            O => \N__5716\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_0\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__5713\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_0\
        );

    \I__835\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5703\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__5703\,
            I => \U712_CHIP_RAM.m93_i_a2_4\
        );

    \I__833\ : IoInMux
    port map (
            O => \N__5700\,
            I => \N__5697\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__5697\,
            I => \N__5694\
        );

    \I__831\ : Span12Mux_s7_h
    port map (
            O => \N__5694\,
            I => \N__5691\
        );

    \I__830\ : Span12Mux_h
    port map (
            O => \N__5691\,
            I => \N__5688\
        );

    \I__829\ : Odrv12
    port map (
            O => \N__5688\,
            I => \CMA_c_8\
        );

    \I__828\ : InMux
    port map (
            O => \N__5685\,
            I => \N__5682\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__5682\,
            I => \N__5679\
        );

    \I__826\ : Odrv4
    port map (
            O => \N__5679\,
            I => \U712_CHIP_RAM.CMA_5_i_0_9\
        );

    \I__825\ : InMux
    port map (
            O => \N__5676\,
            I => \N__5673\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__5673\,
            I => \N__5670\
        );

    \I__823\ : Span4Mux_v
    port map (
            O => \N__5670\,
            I => \N__5667\
        );

    \I__822\ : Span4Mux_v
    port map (
            O => \N__5667\,
            I => \N__5664\
        );

    \I__821\ : Span4Mux_v
    port map (
            O => \N__5664\,
            I => \N__5661\
        );

    \I__820\ : Sp12to4
    port map (
            O => \N__5661\,
            I => \N__5658\
        );

    \I__819\ : Odrv12
    port map (
            O => \N__5658\,
            I => \A_c_19\
        );

    \I__818\ : IoInMux
    port map (
            O => \N__5655\,
            I => \N__5652\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__5652\,
            I => \N__5649\
        );

    \I__816\ : Span12Mux_s7_h
    port map (
            O => \N__5649\,
            I => \N__5646\
        );

    \I__815\ : Span12Mux_h
    port map (
            O => \N__5646\,
            I => \N__5643\
        );

    \I__814\ : Odrv12
    port map (
            O => \N__5643\,
            I => \CMA_c_9\
        );

    \I__813\ : InMux
    port map (
            O => \N__5640\,
            I => \N__5637\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5637\,
            I => \U712_CHIP_RAM.m123_i_2\
        );

    \I__811\ : CascadeMux
    port map (
            O => \N__5634\,
            I => \N__5630\
        );

    \I__810\ : InMux
    port map (
            O => \N__5633\,
            I => \N__5626\
        );

    \I__809\ : InMux
    port map (
            O => \N__5630\,
            I => \N__5623\
        );

    \I__808\ : InMux
    port map (
            O => \N__5629\,
            I => \N__5620\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__5626\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__5623\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__5620\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__804\ : InMux
    port map (
            O => \N__5613\,
            I => \N__5610\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5610\,
            I => \U712_CHIP_RAM.N_190\
        );

    \I__802\ : InMux
    port map (
            O => \N__5607\,
            I => \N__5604\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__5604\,
            I => \N__5600\
        );

    \I__800\ : InMux
    port map (
            O => \N__5603\,
            I => \N__5597\
        );

    \I__799\ : Odrv4
    port map (
            O => \N__5600\,
            I => \U712_CHIP_RAM.N_476\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__5597\,
            I => \U712_CHIP_RAM.N_476\
        );

    \I__797\ : InMux
    port map (
            O => \N__5592\,
            I => \N__5589\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__5589\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1\
        );

    \I__795\ : InMux
    port map (
            O => \N__5586\,
            I => \N__5583\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__5583\,
            I => \U712_CHIP_RAM.N_344\
        );

    \I__793\ : CascadeMux
    port map (
            O => \N__5580\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1_cascade_\
        );

    \I__792\ : InMux
    port map (
            O => \N__5577\,
            I => \N__5573\
        );

    \I__791\ : InMux
    port map (
            O => \N__5576\,
            I => \N__5568\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__5573\,
            I => \N__5565\
        );

    \I__789\ : InMux
    port map (
            O => \N__5572\,
            I => \N__5562\
        );

    \I__788\ : InMux
    port map (
            O => \N__5571\,
            I => \N__5559\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5568\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__786\ : Odrv4
    port map (
            O => \N__5565\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__5562\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__5559\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__5550\,
            I => \N__5539\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__5549\,
            I => \N__5536\
        );

    \I__781\ : InMux
    port map (
            O => \N__5548\,
            I => \N__5533\
        );

    \I__780\ : InMux
    port map (
            O => \N__5547\,
            I => \N__5528\
        );

    \I__779\ : InMux
    port map (
            O => \N__5546\,
            I => \N__5528\
        );

    \I__778\ : InMux
    port map (
            O => \N__5545\,
            I => \N__5525\
        );

    \I__777\ : CascadeMux
    port map (
            O => \N__5544\,
            I => \N__5520\
        );

    \I__776\ : InMux
    port map (
            O => \N__5543\,
            I => \N__5517\
        );

    \I__775\ : InMux
    port map (
            O => \N__5542\,
            I => \N__5510\
        );

    \I__774\ : InMux
    port map (
            O => \N__5539\,
            I => \N__5510\
        );

    \I__773\ : InMux
    port map (
            O => \N__5536\,
            I => \N__5510\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__5533\,
            I => \N__5507\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__5528\,
            I => \N__5504\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__5525\,
            I => \N__5498\
        );

    \I__769\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5495\
        );

    \I__768\ : InMux
    port map (
            O => \N__5523\,
            I => \N__5492\
        );

    \I__767\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5489\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__5517\,
            I => \N__5484\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__5510\,
            I => \N__5484\
        );

    \I__764\ : Span4Mux_v
    port map (
            O => \N__5507\,
            I => \N__5479\
        );

    \I__763\ : Span4Mux_v
    port map (
            O => \N__5504\,
            I => \N__5479\
        );

    \I__762\ : InMux
    port map (
            O => \N__5503\,
            I => \N__5474\
        );

    \I__761\ : InMux
    port map (
            O => \N__5502\,
            I => \N__5474\
        );

    \I__760\ : InMux
    port map (
            O => \N__5501\,
            I => \N__5471\
        );

    \I__759\ : Span4Mux_h
    port map (
            O => \N__5498\,
            I => \N__5468\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5495\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__5492\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__5489\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__755\ : Odrv4
    port map (
            O => \N__5484\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__754\ : Odrv4
    port map (
            O => \N__5479\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__5474\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__5471\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__751\ : Odrv4
    port map (
            O => \N__5468\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__750\ : InMux
    port map (
            O => \N__5451\,
            I => \N__5447\
        );

    \I__749\ : InMux
    port map (
            O => \N__5450\,
            I => \N__5437\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__5447\,
            I => \N__5434\
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__5446\,
            I => \N__5429\
        );

    \I__746\ : InMux
    port map (
            O => \N__5445\,
            I => \N__5425\
        );

    \I__745\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5422\
        );

    \I__744\ : InMux
    port map (
            O => \N__5443\,
            I => \N__5410\
        );

    \I__743\ : InMux
    port map (
            O => \N__5442\,
            I => \N__5410\
        );

    \I__742\ : InMux
    port map (
            O => \N__5441\,
            I => \N__5410\
        );

    \I__741\ : InMux
    port map (
            O => \N__5440\,
            I => \N__5410\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__5437\,
            I => \N__5407\
        );

    \I__739\ : Span4Mux_v
    port map (
            O => \N__5434\,
            I => \N__5404\
        );

    \I__738\ : InMux
    port map (
            O => \N__5433\,
            I => \N__5401\
        );

    \I__737\ : InMux
    port map (
            O => \N__5432\,
            I => \N__5398\
        );

    \I__736\ : InMux
    port map (
            O => \N__5429\,
            I => \N__5395\
        );

    \I__735\ : InMux
    port map (
            O => \N__5428\,
            I => \N__5392\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__5425\,
            I => \N__5387\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__5422\,
            I => \N__5387\
        );

    \I__732\ : InMux
    port map (
            O => \N__5421\,
            I => \N__5382\
        );

    \I__731\ : InMux
    port map (
            O => \N__5420\,
            I => \N__5382\
        );

    \I__730\ : InMux
    port map (
            O => \N__5419\,
            I => \N__5379\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__5410\,
            I => \N__5374\
        );

    \I__728\ : Span4Mux_h
    port map (
            O => \N__5407\,
            I => \N__5374\
        );

    \I__727\ : Odrv4
    port map (
            O => \N__5404\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5401\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__5398\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__5395\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__5392\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__722\ : Odrv4
    port map (
            O => \N__5387\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__5382\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__5379\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__719\ : Odrv4
    port map (
            O => \N__5374\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__718\ : InMux
    port map (
            O => \N__5355\,
            I => \N__5349\
        );

    \I__717\ : InMux
    port map (
            O => \N__5354\,
            I => \N__5343\
        );

    \I__716\ : InMux
    port map (
            O => \N__5353\,
            I => \N__5343\
        );

    \I__715\ : InMux
    port map (
            O => \N__5352\,
            I => \N__5340\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__5349\,
            I => \N__5336\
        );

    \I__713\ : InMux
    port map (
            O => \N__5348\,
            I => \N__5333\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__5343\,
            I => \N__5328\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__5340\,
            I => \N__5328\
        );

    \I__710\ : InMux
    port map (
            O => \N__5339\,
            I => \N__5325\
        );

    \I__709\ : Odrv4
    port map (
            O => \N__5336\,
            I => \U712_CHIP_RAM.N_307\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__5333\,
            I => \U712_CHIP_RAM.N_307\
        );

    \I__707\ : Odrv4
    port map (
            O => \N__5328\,
            I => \U712_CHIP_RAM.N_307\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__5325\,
            I => \U712_CHIP_RAM.N_307\
        );

    \I__705\ : CascadeMux
    port map (
            O => \N__5316\,
            I => \U712_CHIP_RAM.N_551_cascade_\
        );

    \I__704\ : CascadeMux
    port map (
            O => \N__5313\,
            I => \N__5310\
        );

    \I__703\ : InMux
    port map (
            O => \N__5310\,
            I => \N__5307\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5307\,
            I => \N__5302\
        );

    \I__701\ : InMux
    port map (
            O => \N__5306\,
            I => \N__5299\
        );

    \I__700\ : InMux
    port map (
            O => \N__5305\,
            I => \N__5296\
        );

    \I__699\ : Odrv4
    port map (
            O => \N__5302\,
            I => \U712_CHIP_RAM.N_304\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__5299\,
            I => \U712_CHIP_RAM.N_304\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__5296\,
            I => \U712_CHIP_RAM.N_304\
        );

    \I__696\ : CascadeMux
    port map (
            O => \N__5289\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_1_1_cascade_\
        );

    \I__695\ : InMux
    port map (
            O => \N__5286\,
            I => \N__5283\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__5283\,
            I => \U712_CHIP_RAM.N_378\
        );

    \I__693\ : InMux
    port map (
            O => \N__5280\,
            I => \N__5271\
        );

    \I__692\ : InMux
    port map (
            O => \N__5279\,
            I => \N__5271\
        );

    \I__691\ : InMux
    port map (
            O => \N__5278\,
            I => \N__5271\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__5271\,
            I => \N__5267\
        );

    \I__689\ : InMux
    port map (
            O => \N__5270\,
            I => \N__5263\
        );

    \I__688\ : Span4Mux_h
    port map (
            O => \N__5267\,
            I => \N__5260\
        );

    \I__687\ : InMux
    port map (
            O => \N__5266\,
            I => \N__5257\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__5263\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__685\ : Odrv4
    port map (
            O => \N__5260\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__5257\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__683\ : CascadeMux
    port map (
            O => \N__5250\,
            I => \N__5247\
        );

    \I__682\ : InMux
    port map (
            O => \N__5247\,
            I => \N__5242\
        );

    \I__681\ : InMux
    port map (
            O => \N__5246\,
            I => \N__5237\
        );

    \I__680\ : InMux
    port map (
            O => \N__5245\,
            I => \N__5237\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__5242\,
            I => \N__5231\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__5237\,
            I => \N__5231\
        );

    \I__677\ : InMux
    port map (
            O => \N__5236\,
            I => \N__5227\
        );

    \I__676\ : Span4Mux_h
    port map (
            O => \N__5231\,
            I => \N__5224\
        );

    \I__675\ : InMux
    port map (
            O => \N__5230\,
            I => \N__5221\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__5227\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__673\ : Odrv4
    port map (
            O => \N__5224\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__5221\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__671\ : InMux
    port map (
            O => \N__5214\,
            I => \N__5205\
        );

    \I__670\ : InMux
    port map (
            O => \N__5213\,
            I => \N__5205\
        );

    \I__669\ : InMux
    port map (
            O => \N__5212\,
            I => \N__5205\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__5205\,
            I => \U712_CHIP_RAM.SDRAM_CMDs_0_4\
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__5202\,
            I => \U712_CHIP_RAM.N_396_cascade_\
        );

    \I__666\ : InMux
    port map (
            O => \N__5199\,
            I => \N__5196\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__5196\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_0_2\
        );

    \I__664\ : InMux
    port map (
            O => \N__5193\,
            I => \N__5190\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__5190\,
            I => \U712_CHIP_RAM.N_397\
        );

    \I__662\ : InMux
    port map (
            O => \N__5187\,
            I => \N__5184\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__5184\,
            I => \N__5181\
        );

    \I__660\ : Span4Mux_h
    port map (
            O => \N__5181\,
            I => \N__5178\
        );

    \I__659\ : Odrv4
    port map (
            O => \N__5178\,
            I => \U712_CHIP_RAM.N_555\
        );

    \I__658\ : InMux
    port map (
            O => \N__5175\,
            I => \N__5172\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__5172\,
            I => \N__5169\
        );

    \I__656\ : Span4Mux_h
    port map (
            O => \N__5169\,
            I => \N__5166\
        );

    \I__655\ : Odrv4
    port map (
            O => \N__5166\,
            I => \U712_CHIP_RAM.N_449\
        );

    \I__654\ : CascadeMux
    port map (
            O => \N__5163\,
            I => \N__5160\
        );

    \I__653\ : InMux
    port map (
            O => \N__5160\,
            I => \N__5154\
        );

    \I__652\ : InMux
    port map (
            O => \N__5159\,
            I => \N__5154\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__5154\,
            I => \N__5151\
        );

    \I__650\ : Span4Mux_h
    port map (
            O => \N__5151\,
            I => \N__5148\
        );

    \I__649\ : Odrv4
    port map (
            O => \N__5148\,
            I => \U712_CHIP_RAM.SDRAM_CMDs_0_1\
        );

    \I__648\ : InMux
    port map (
            O => \N__5145\,
            I => \N__5142\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__5142\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_1_3\
        );

    \I__646\ : CEMux
    port map (
            O => \N__5139\,
            I => \N__5136\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__5136\,
            I => \N__5133\
        );

    \I__644\ : Span4Mux_v
    port map (
            O => \N__5133\,
            I => \N__5130\
        );

    \I__643\ : Odrv4
    port map (
            O => \N__5130\,
            I => \U712_CHIP_RAM.N_194_0\
        );

    \I__642\ : InMux
    port map (
            O => \N__5127\,
            I => \N__5124\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__5124\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa\
        );

    \I__640\ : CascadeMux
    port map (
            O => \N__5121\,
            I => \N__5117\
        );

    \I__639\ : InMux
    port map (
            O => \N__5120\,
            I => \N__5105\
        );

    \I__638\ : InMux
    port map (
            O => \N__5117\,
            I => \N__5105\
        );

    \I__637\ : InMux
    port map (
            O => \N__5116\,
            I => \N__5099\
        );

    \I__636\ : InMux
    port map (
            O => \N__5115\,
            I => \N__5099\
        );

    \I__635\ : InMux
    port map (
            O => \N__5114\,
            I => \N__5094\
        );

    \I__634\ : InMux
    port map (
            O => \N__5113\,
            I => \N__5094\
        );

    \I__633\ : InMux
    port map (
            O => \N__5112\,
            I => \N__5091\
        );

    \I__632\ : InMux
    port map (
            O => \N__5111\,
            I => \N__5080\
        );

    \I__631\ : InMux
    port map (
            O => \N__5110\,
            I => \N__5080\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__5105\,
            I => \N__5077\
        );

    \I__629\ : InMux
    port map (
            O => \N__5104\,
            I => \N__5074\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__5099\,
            I => \N__5069\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__5094\,
            I => \N__5069\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__5091\,
            I => \N__5066\
        );

    \I__625\ : InMux
    port map (
            O => \N__5090\,
            I => \N__5061\
        );

    \I__624\ : InMux
    port map (
            O => \N__5089\,
            I => \N__5061\
        );

    \I__623\ : InMux
    port map (
            O => \N__5088\,
            I => \N__5054\
        );

    \I__622\ : InMux
    port map (
            O => \N__5087\,
            I => \N__5054\
        );

    \I__621\ : InMux
    port map (
            O => \N__5086\,
            I => \N__5054\
        );

    \I__620\ : InMux
    port map (
            O => \N__5085\,
            I => \N__5051\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__5080\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__618\ : Odrv4
    port map (
            O => \N__5077\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__5074\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__616\ : Odrv4
    port map (
            O => \N__5069\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__615\ : Odrv4
    port map (
            O => \N__5066\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__5061\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__5054\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__5051\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__611\ : InMux
    port map (
            O => \N__5034\,
            I => \N__5031\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__5031\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__609\ : IoInMux
    port map (
            O => \N__5028\,
            I => \N__5025\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__5025\,
            I => \N__5022\
        );

    \I__607\ : IoSpan4Mux
    port map (
            O => \N__5022\,
            I => \N__5019\
        );

    \I__606\ : Sp12to4
    port map (
            O => \N__5019\,
            I => \N__5016\
        );

    \I__605\ : Span12Mux_s7_h
    port map (
            O => \N__5016\,
            I => \N__5013\
        );

    \I__604\ : Span12Mux_h
    port map (
            O => \N__5013\,
            I => \N__5010\
        );

    \I__603\ : Odrv12
    port map (
            O => \N__5010\,
            I => \CMA_c_6\
        );

    \I__602\ : InMux
    port map (
            O => \N__5007\,
            I => \N__5004\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__5004\,
            I => \N__5001\
        );

    \I__600\ : Sp12to4
    port map (
            O => \N__5001\,
            I => \N__4998\
        );

    \I__599\ : Span12Mux_v
    port map (
            O => \N__4998\,
            I => \N__4995\
        );

    \I__598\ : Span12Mux_h
    port map (
            O => \N__4995\,
            I => \N__4992\
        );

    \I__597\ : Odrv12
    port map (
            O => \N__4992\,
            I => \A_c_12\
        );

    \I__596\ : InMux
    port map (
            O => \N__4989\,
            I => \N__4986\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__4986\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\
        );

    \I__594\ : CascadeMux
    port map (
            O => \N__4983\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\
        );

    \I__593\ : InMux
    port map (
            O => \N__4980\,
            I => \N__4977\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__4977\,
            I => \N__4974\
        );

    \I__591\ : Sp12to4
    port map (
            O => \N__4974\,
            I => \N__4971\
        );

    \I__590\ : Span12Mux_v
    port map (
            O => \N__4971\,
            I => \N__4968\
        );

    \I__589\ : Span12Mux_h
    port map (
            O => \N__4968\,
            I => \N__4965\
        );

    \I__588\ : Odrv12
    port map (
            O => \N__4965\,
            I => \A_c_16\
        );

    \I__587\ : InMux
    port map (
            O => \N__4962\,
            I => \N__4959\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__4959\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\
        );

    \I__585\ : IoInMux
    port map (
            O => \N__4956\,
            I => \N__4953\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__4953\,
            I => \N__4950\
        );

    \I__583\ : Span4Mux_s1_v
    port map (
            O => \N__4950\,
            I => \N__4947\
        );

    \I__582\ : Span4Mux_v
    port map (
            O => \N__4947\,
            I => \N__4944\
        );

    \I__581\ : Span4Mux_v
    port map (
            O => \N__4944\,
            I => \N__4941\
        );

    \I__580\ : Odrv4
    port map (
            O => \N__4941\,
            I => \VBENn_c\
        );

    \I__579\ : InMux
    port map (
            O => \N__4938\,
            I => \N__4935\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__4935\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_6\
        );

    \I__577\ : InMux
    port map (
            O => \N__4932\,
            I => \N__4928\
        );

    \I__576\ : InMux
    port map (
            O => \N__4931\,
            I => \N__4925\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__4928\,
            I => \U712_CHIP_RAM.N_194\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__4925\,
            I => \U712_CHIP_RAM.N_194\
        );

    \I__573\ : CascadeMux
    port map (
            O => \N__4920\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_5_cascade_\
        );

    \I__572\ : InMux
    port map (
            O => \N__4917\,
            I => \N__4914\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__4914\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_1\
        );

    \I__570\ : InMux
    port map (
            O => \N__4911\,
            I => \N__4908\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__4908\,
            I => \N__4903\
        );

    \I__568\ : CascadeMux
    port map (
            O => \N__4907\,
            I => \N__4900\
        );

    \I__567\ : InMux
    port map (
            O => \N__4906\,
            I => \N__4897\
        );

    \I__566\ : Span4Mux_h
    port map (
            O => \N__4903\,
            I => \N__4894\
        );

    \I__565\ : InMux
    port map (
            O => \N__4900\,
            I => \N__4891\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__4897\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__563\ : Odrv4
    port map (
            O => \N__4894\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__4891\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__561\ : InMux
    port map (
            O => \N__4884\,
            I => \N__4881\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__4881\,
            I => \N__4877\
        );

    \I__559\ : InMux
    port map (
            O => \N__4880\,
            I => \N__4873\
        );

    \I__558\ : Span4Mux_h
    port map (
            O => \N__4877\,
            I => \N__4870\
        );

    \I__557\ : InMux
    port map (
            O => \N__4876\,
            I => \N__4867\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__4873\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__555\ : Odrv4
    port map (
            O => \N__4870\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__4867\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__553\ : CascadeMux
    port map (
            O => \N__4860\,
            I => \N__4855\
        );

    \I__552\ : InMux
    port map (
            O => \N__4859\,
            I => \N__4852\
        );

    \I__551\ : InMux
    port map (
            O => \N__4858\,
            I => \N__4849\
        );

    \I__550\ : InMux
    port map (
            O => \N__4855\,
            I => \N__4846\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4852\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_1\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__4849\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_1\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4846\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_1\
        );

    \I__546\ : InMux
    port map (
            O => \N__4839\,
            I => \N__4835\
        );

    \I__545\ : InMux
    port map (
            O => \N__4838\,
            I => \N__4832\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__4835\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_2\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4832\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_2\
        );

    \I__542\ : InMux
    port map (
            O => \N__4827\,
            I => \U712_CHIP_RAM.un3_DBR_COUNT_cry_1\
        );

    \I__541\ : InMux
    port map (
            O => \N__4824\,
            I => \N__4820\
        );

    \I__540\ : InMux
    port map (
            O => \N__4823\,
            I => \N__4817\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__4820\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_3\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__4817\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_3\
        );

    \I__537\ : InMux
    port map (
            O => \N__4812\,
            I => \U712_CHIP_RAM.un3_DBR_COUNT_cry_2\
        );

    \I__536\ : InMux
    port map (
            O => \N__4809\,
            I => \N__4805\
        );

    \I__535\ : InMux
    port map (
            O => \N__4808\,
            I => \N__4802\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__4805\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_4\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__4802\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_4\
        );

    \I__532\ : InMux
    port map (
            O => \N__4797\,
            I => \U712_CHIP_RAM.un3_DBR_COUNT_cry_3\
        );

    \I__531\ : InMux
    port map (
            O => \N__4794\,
            I => \N__4790\
        );

    \I__530\ : InMux
    port map (
            O => \N__4793\,
            I => \N__4787\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__4790\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_5\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__4787\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_5\
        );

    \I__527\ : InMux
    port map (
            O => \N__4782\,
            I => \U712_CHIP_RAM.un3_DBR_COUNT_cry_4\
        );

    \I__526\ : InMux
    port map (
            O => \N__4779\,
            I => \U712_CHIP_RAM.un3_DBR_COUNT_cry_5\
        );

    \I__525\ : InMux
    port map (
            O => \N__4776\,
            I => \U712_CHIP_RAM.un3_DBR_COUNT_cry_6\
        );

    \I__524\ : InMux
    port map (
            O => \N__4773\,
            I => \N__4769\
        );

    \I__523\ : InMux
    port map (
            O => \N__4772\,
            I => \N__4766\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__4769\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_7\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4766\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_7\
        );

    \I__520\ : InMux
    port map (
            O => \N__4761\,
            I => \N__4757\
        );

    \I__519\ : InMux
    port map (
            O => \N__4760\,
            I => \N__4754\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__4757\,
            I => \N__4751\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__4754\,
            I => \N__4748\
        );

    \I__516\ : Span4Mux_v
    port map (
            O => \N__4751\,
            I => \N__4745\
        );

    \I__515\ : Span4Mux_v
    port map (
            O => \N__4748\,
            I => \N__4742\
        );

    \I__514\ : Sp12to4
    port map (
            O => \N__4745\,
            I => \N__4737\
        );

    \I__513\ : Sp12to4
    port map (
            O => \N__4742\,
            I => \N__4737\
        );

    \I__512\ : Span12Mux_h
    port map (
            O => \N__4737\,
            I => \N__4734\
        );

    \I__511\ : Span12Mux_v
    port map (
            O => \N__4734\,
            I => \N__4731\
        );

    \I__510\ : Odrv12
    port map (
            O => \N__4731\,
            I => \DBRn_c\
        );

    \I__509\ : CascadeMux
    port map (
            O => \N__4728\,
            I => \U712_CHIP_RAM.N_307_cascade_\
        );

    \I__508\ : CascadeMux
    port map (
            O => \N__4725\,
            I => \U712_CHIP_RAM.N_467_cascade_\
        );

    \I__507\ : CascadeMux
    port map (
            O => \N__4722\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\
        );

    \I__506\ : InMux
    port map (
            O => \N__4719\,
            I => \N__4716\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4716\,
            I => \N__4713\
        );

    \I__504\ : Span4Mux_h
    port map (
            O => \N__4713\,
            I => \N__4710\
        );

    \I__503\ : Odrv4
    port map (
            O => \N__4710\,
            I => \U712_CHIP_RAM.N_440\
        );

    \I__502\ : CascadeMux
    port map (
            O => \N__4707\,
            I => \U712_CHIP_RAM.N_304_cascade_\
        );

    \I__501\ : CascadeMux
    port map (
            O => \N__4704\,
            I => \U712_CHIP_RAM.N_312_cascade_\
        );

    \I__500\ : CascadeMux
    port map (
            O => \N__4701\,
            I => \N__4698\
        );

    \I__499\ : InMux
    port map (
            O => \N__4698\,
            I => \N__4695\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__4695\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__497\ : InMux
    port map (
            O => \N__4692\,
            I => \N__4679\
        );

    \I__496\ : InMux
    port map (
            O => \N__4691\,
            I => \N__4679\
        );

    \I__495\ : InMux
    port map (
            O => \N__4690\,
            I => \N__4679\
        );

    \I__494\ : InMux
    port map (
            O => \N__4689\,
            I => \N__4676\
        );

    \I__493\ : InMux
    port map (
            O => \N__4688\,
            I => \N__4669\
        );

    \I__492\ : InMux
    port map (
            O => \N__4687\,
            I => \N__4669\
        );

    \I__491\ : InMux
    port map (
            O => \N__4686\,
            I => \N__4669\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__4679\,
            I => \U712_CHIP_RAM.N_39\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4676\,
            I => \U712_CHIP_RAM.N_39\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__4669\,
            I => \U712_CHIP_RAM.N_39\
        );

    \I__487\ : InMux
    port map (
            O => \N__4662\,
            I => \N__4659\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__4659\,
            I => \N__4655\
        );

    \I__485\ : InMux
    port map (
            O => \N__4658\,
            I => \N__4652\
        );

    \I__484\ : Sp12to4
    port map (
            O => \N__4655\,
            I => \N__4649\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__4652\,
            I => \U712_CHIP_RAM.N_326\
        );

    \I__482\ : Odrv12
    port map (
            O => \N__4649\,
            I => \U712_CHIP_RAM.N_326\
        );

    \I__481\ : CascadeMux
    port map (
            O => \N__4644\,
            I => \U712_CHIP_RAM.N_39_cascade_\
        );

    \I__480\ : CEMux
    port map (
            O => \N__4641\,
            I => \N__4638\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4638\,
            I => \N__4634\
        );

    \I__478\ : CEMux
    port map (
            O => \N__4637\,
            I => \N__4631\
        );

    \I__477\ : Sp12to4
    port map (
            O => \N__4634\,
            I => \N__4626\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__4631\,
            I => \N__4626\
        );

    \I__475\ : Odrv12
    port map (
            O => \N__4626\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__474\ : CascadeMux
    port map (
            O => \N__4623\,
            I => \N__4620\
        );

    \I__473\ : InMux
    port map (
            O => \N__4620\,
            I => \N__4616\
        );

    \I__472\ : InMux
    port map (
            O => \N__4619\,
            I => \N__4613\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__4616\,
            I => \U712_CHIP_RAM.N_20_0\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4613\,
            I => \U712_CHIP_RAM.N_20_0\
        );

    \I__469\ : InMux
    port map (
            O => \N__4608\,
            I => \N__4605\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__4605\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_0_a3_0_a2_0\
        );

    \I__467\ : InMux
    port map (
            O => \N__4602\,
            I => \N__4599\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__4599\,
            I => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\
        );

    \I__465\ : InMux
    port map (
            O => \N__4596\,
            I => \N__4593\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__4593\,
            I => \U712_CHIP_RAM.m101_i_1\
        );

    \I__463\ : CascadeMux
    port map (
            O => \N__4590\,
            I => \U712_CHIP_RAM.N_305_cascade_\
        );

    \I__462\ : InMux
    port map (
            O => \N__4587\,
            I => \N__4584\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__4584\,
            I => \U712_CHIP_RAM.N_376\
        );

    \I__460\ : CascadeMux
    port map (
            O => \N__4581\,
            I => \U712_CHIP_RAM.m101_i_0_cascade_\
        );

    \I__459\ : InMux
    port map (
            O => \N__4578\,
            I => \N__4575\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__4575\,
            I => \U712_CHIP_RAM.m101_i_2\
        );

    \I__457\ : InMux
    port map (
            O => \N__4572\,
            I => \N__4569\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__4569\,
            I => \N__4566\
        );

    \I__455\ : Span12Mux_v
    port map (
            O => \N__4566\,
            I => \N__4563\
        );

    \I__454\ : Odrv12
    port map (
            O => \N__4563\,
            I => \A_c_5\
        );

    \I__453\ : InMux
    port map (
            O => \N__4560\,
            I => \N__4557\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__4557\,
            I => \N__4554\
        );

    \I__451\ : Span4Mux_h
    port map (
            O => \N__4554\,
            I => \N__4551\
        );

    \I__450\ : Sp12to4
    port map (
            O => \N__4551\,
            I => \N__4548\
        );

    \I__449\ : Span12Mux_v
    port map (
            O => \N__4548\,
            I => \N__4545\
        );

    \I__448\ : Odrv12
    port map (
            O => \N__4545\,
            I => \A_c_18\
        );

    \I__447\ : CascadeMux
    port map (
            O => \N__4542\,
            I => \U712_CHIP_RAM.N_436_cascade_\
        );

    \I__446\ : CascadeMux
    port map (
            O => \N__4539\,
            I => \U712_CHIP_RAM.N_194_cascade_\
        );

    \I__445\ : InMux
    port map (
            O => \N__4536\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__444\ : InMux
    port map (
            O => \N__4533\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__443\ : InMux
    port map (
            O => \N__4530\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__442\ : InMux
    port map (
            O => \N__4527\,
            I => \N__4524\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__4524\,
            I => \N__4521\
        );

    \I__440\ : Span4Mux_v
    port map (
            O => \N__4521\,
            I => \N__4518\
        );

    \I__439\ : Sp12to4
    port map (
            O => \N__4518\,
            I => \N__4515\
        );

    \I__438\ : Odrv12
    port map (
            O => \N__4515\,
            I => \A_c_8\
        );

    \I__437\ : InMux
    port map (
            O => \N__4512\,
            I => \N__4509\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__4509\,
            I => \N__4506\
        );

    \I__435\ : Span12Mux_h
    port map (
            O => \N__4506\,
            I => \N__4503\
        );

    \I__434\ : Span12Mux_v
    port map (
            O => \N__4503\,
            I => \N__4500\
        );

    \I__433\ : Odrv12
    port map (
            O => \N__4500\,
            I => \A_c_2\
        );

    \I__432\ : InMux
    port map (
            O => \N__4497\,
            I => \N__4494\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__4494\,
            I => \N__4491\
        );

    \I__430\ : Span4Mux_h
    port map (
            O => \N__4491\,
            I => \N__4488\
        );

    \I__429\ : Sp12to4
    port map (
            O => \N__4488\,
            I => \N__4485\
        );

    \I__428\ : Span12Mux_v
    port map (
            O => \N__4485\,
            I => \N__4482\
        );

    \I__427\ : Odrv12
    port map (
            O => \N__4482\,
            I => \A_c_3\
        );

    \I__426\ : InMux
    port map (
            O => \N__4479\,
            I => \N__4476\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__4476\,
            I => \N__4473\
        );

    \I__424\ : Span4Mux_v
    port map (
            O => \N__4473\,
            I => \N__4470\
        );

    \I__423\ : Span4Mux_v
    port map (
            O => \N__4470\,
            I => \N__4467\
        );

    \I__422\ : Sp12to4
    port map (
            O => \N__4467\,
            I => \N__4464\
        );

    \I__421\ : Odrv12
    port map (
            O => \N__4464\,
            I => \A_c_4\
        );

    \I__420\ : InMux
    port map (
            O => \N__4461\,
            I => \N__4458\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__4458\,
            I => \N__4455\
        );

    \I__418\ : Span4Mux_v
    port map (
            O => \N__4455\,
            I => \N__4452\
        );

    \I__417\ : Sp12to4
    port map (
            O => \N__4452\,
            I => \N__4449\
        );

    \I__416\ : Odrv12
    port map (
            O => \N__4449\,
            I => \A_c_7\
        );

    \I__415\ : IoInMux
    port map (
            O => \N__4446\,
            I => \N__4443\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__4443\,
            I => \N__4440\
        );

    \I__413\ : IoSpan4Mux
    port map (
            O => \N__4440\,
            I => \N__4437\
        );

    \I__412\ : Sp12to4
    port map (
            O => \N__4437\,
            I => \N__4434\
        );

    \I__411\ : Span12Mux_s9_h
    port map (
            O => \N__4434\,
            I => \N__4431\
        );

    \I__410\ : Span12Mux_h
    port map (
            O => \N__4431\,
            I => \N__4427\
        );

    \I__409\ : InMux
    port map (
            O => \N__4430\,
            I => \N__4424\
        );

    \I__408\ : Odrv12
    port map (
            O => \N__4427\,
            I => \CLK_EN_c\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__4424\,
            I => \CLK_EN_c\
        );

    \I__406\ : CascadeMux
    port map (
            O => \N__4419\,
            I => \U712_CHIP_RAM.m77_0_a2_0_2_cascade_\
        );

    \I__405\ : InMux
    port map (
            O => \N__4416\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__404\ : InMux
    port map (
            O => \N__4413\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__403\ : InMux
    port map (
            O => \N__4410\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__402\ : InMux
    port map (
            O => \N__4407\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__401\ : IoInMux
    port map (
            O => \N__4404\,
            I => \N__4401\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__4401\,
            I => \N__4398\
        );

    \I__399\ : Span4Mux_s3_v
    port map (
            O => \N__4398\,
            I => \N__4395\
        );

    \I__398\ : Span4Mux_h
    port map (
            O => \N__4395\,
            I => \N__4392\
        );

    \I__397\ : Odrv4
    port map (
            O => \N__4392\,
            I => \CLK80_PLL_i_i\
        );

    \I__396\ : InMux
    port map (
            O => \N__4389\,
            I => \N__4386\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__4386\,
            I => \N__4383\
        );

    \I__394\ : Span12Mux_h
    port map (
            O => \N__4383\,
            I => \N__4380\
        );

    \I__393\ : Span12Mux_v
    port map (
            O => \N__4380\,
            I => \N__4377\
        );

    \I__392\ : Odrv12
    port map (
            O => \N__4377\,
            I => \REGSPACEn_c\
        );

    \I__391\ : CascadeMux
    port map (
            O => \N__4374\,
            I => \U712_CHIP_RAM.N_555_cascade_\
        );

    \I__390\ : CascadeMux
    port map (
            O => \N__4371\,
            I => \U712_CHIP_RAM.N_390_cascade_\
        );

    \I__389\ : InMux
    port map (
            O => \N__4368\,
            I => \N__4365\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__4365\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_2_0\
        );

    \I__387\ : CascadeMux
    port map (
            O => \N__4362\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_2_3_cascade_\
        );

    \I__386\ : InMux
    port map (
            O => \N__4359\,
            I => \N__4356\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__4356\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_2_2\
        );

    \I__384\ : IoInMux
    port map (
            O => \N__4353\,
            I => \N__4350\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__4350\,
            I => \N__4347\
        );

    \I__382\ : Odrv12
    port map (
            O => \N__4347\,
            I => \DBRn_c_i_0\
        );

    \I__381\ : IoInMux
    port map (
            O => \N__4344\,
            I => \N__4341\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__4341\,
            I => \N__4338\
        );

    \I__379\ : Span4Mux_s0_v
    port map (
            O => \N__4338\,
            I => \N__4335\
        );

    \I__378\ : Span4Mux_v
    port map (
            O => \N__4335\,
            I => \N__4332\
        );

    \I__377\ : Sp12to4
    port map (
            O => \N__4332\,
            I => \N__4329\
        );

    \I__376\ : Span12Mux_h
    port map (
            O => \N__4329\,
            I => \N__4326\
        );

    \I__375\ : Span12Mux_v
    port map (
            O => \N__4326\,
            I => \N__4323\
        );

    \I__374\ : Odrv12
    port map (
            O => \N__4323\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            I => \N__7492\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__7491\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            I => \N__7486\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            I => \N__7489\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__7493\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            I => \N__7487\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            I => \N__7490\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__7494\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_10_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_10_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_7_0_\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8468\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__9195\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4353\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8169\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9828\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8615\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_3_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9993\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6486\,
            in2 => \_gnd_net_\,
            in3 => \N__4389\,
            lcout => \U712_REG_SM.N_402\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_3_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100100010"
        )
    port map (
            in0 => \N__5114\,
            in1 => \N__6199\,
            in2 => \N__5550\,
            in3 => \N__6081\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIMT791_1_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6196\,
            in1 => \N__5441\,
            in2 => \_gnd_net_\,
            in3 => \N__5113\,
            lcout => \U712_CHIP_RAM.N_555\,
            ltout => \U712_CHIP_RAM.N_555_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__5542\,
            in1 => \_gnd_net_\,
            in2 => \N__4374\,
            in3 => \N__5633\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_390_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101111"
        )
    port map (
            in0 => \N__5355\,
            in1 => \_gnd_net_\,
            in2 => \N__4371\,
            in3 => \N__4368\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMDsr_2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101111001000"
        )
    port map (
            in0 => \N__4359\,
            in1 => \N__4932\,
            in2 => \N__4362\,
            in3 => \N__7904\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9953\,
            ce => 'H',
            sr => \N__9799\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__6200\,
            in1 => \_gnd_net_\,
            in2 => \N__6097\,
            in3 => \N__5443\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__5440\,
            in1 => \N__6197\,
            in2 => \N__5549\,
            in3 => \N__6077\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDs_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_2_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__6198\,
            in1 => \_gnd_net_\,
            in2 => \N__6096\,
            in3 => \N__5442\,
            lcout => \U712_CHIP_RAM.N_449\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011111100000100"
        )
    port map (
            in0 => \N__5354\,
            in1 => \N__4608\,
            in2 => \N__4623\,
            in3 => \N__4430\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9959\,
            ce => 'H',
            sr => \N__9794\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6240\,
            in1 => \N__5433\,
            in2 => \N__6089\,
            in3 => \N__10946\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m77_0_a2_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__5353\,
            in1 => \N__4619\,
            in2 => \N__4419\,
            in3 => \N__5523\,
            lcout => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__7440\,
            in1 => \N__5104\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.LATCH_CLK_6\,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4690\,
            in1 => \N__5432\,
            in2 => \_gnd_net_\,
            in3 => \N__4416\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__9966\,
            ce => \N__4641\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6088\,
            in2 => \_gnd_net_\,
            in3 => \N__4413\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4691\,
            in1 => \N__5524\,
            in2 => \_gnd_net_\,
            in3 => \N__4410\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__9966\,
            ce => \N__4641\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4686\,
            in1 => \N__5270\,
            in2 => \_gnd_net_\,
            in3 => \N__4407\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__9966\,
            ce => \N__4641\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4692\,
            in1 => \N__4880\,
            in2 => \_gnd_net_\,
            in3 => \N__4536\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__9966\,
            ce => \N__4641\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4687\,
            in1 => \N__5236\,
            in2 => \_gnd_net_\,
            in3 => \N__4533\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__9966\,
            ce => \N__4641\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__4906\,
            in1 => \N__4688\,
            in2 => \_gnd_net_\,
            in3 => \N__4530\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9966\,
            ce => \N__4641\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4527\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9972\,
            ce => \N__7551\,
            sr => \N__9784\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4512\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9977\,
            ce => \N__7559\,
            sr => \N__9774\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4497\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9977\,
            ce => \N__7559\,
            sr => \N__9774\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4479\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9977\,
            ce => \N__7559\,
            sr => \N__9774\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4461\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9977\,
            ce => \N__7559\,
            sr => \N__9774\
        );

    \U712_CHIP_RAM.DBR_COUNT_1_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5730\,
            in2 => \_gnd_net_\,
            in3 => \N__4859\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9982\,
            ce => 'H',
            sr => \N__6363\
        );

    \U712_CHIP_RAM.DBR_COUNT_0_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5731\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9982\,
            ce => 'H',
            sr => \N__6363\
        );

    \DBRn_ibuf_RNIBAB_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4761\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4572\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9943\,
            ce => \N__7558\,
            sr => \N__9800\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4560\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9943\,
            ce => \N__7558\,
            sr => \N__9800\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__6596\,
            in1 => \N__8334\,
            in2 => \_gnd_net_\,
            in3 => \N__6627\,
            lcout => \U712_CHIP_RAM.CMA_5_i_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101111010"
        )
    port map (
            in0 => \N__6201\,
            in1 => \N__5445\,
            in2 => \N__6094\,
            in3 => \N__5115\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9183\,
            in3 => \N__6070\,
            lcout => \U712_CHIP_RAM.DBENn_7_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNICN5A2_2_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6069\,
            in1 => \N__6258\,
            in2 => \_gnd_net_\,
            in3 => \N__5629\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_436_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITD0EA_0_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__4578\,
            in1 => \N__4587\,
            in2 => \N__4542\,
            in3 => \N__4596\,
            lcout => \U712_CHIP_RAM.N_194\,
            ltout => \U712_CHIP_RAM.N_194_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIJNSTA_0_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4539\,
            in3 => \N__9827\,
            lcout => \U712_CHIP_RAM.N_194_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIDTSL_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5577\,
            in1 => \N__10944\,
            in2 => \_gnd_net_\,
            in3 => \N__5444\,
            lcout => \U712_CHIP_RAM.N_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6202\,
            in1 => \N__5543\,
            in2 => \N__6095\,
            in3 => \N__5116\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_0_a3_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__10409\,
            in1 => \N__4602\,
            in2 => \N__8712\,
            in3 => \N__5613\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9954\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__6167\,
            in1 => \N__10410\,
            in2 => \_gnd_net_\,
            in3 => \N__5127\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9954\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI3M1M2_1_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__5421\,
            in1 => \N__6165\,
            in2 => \_gnd_net_\,
            in3 => \N__5352\,
            lcout => \U712_CHIP_RAM.m101_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5420\,
            in2 => \_gnd_net_\,
            in3 => \N__5086\,
            lcout => \U712_CHIP_RAM.N_305\,
            ltout => \U712_CHIP_RAM.N_305_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNI7MCB2_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001011"
        )
    port map (
            in0 => \N__6022\,
            in1 => \N__5871\,
            in2 => \N__4590\,
            in3 => \N__5503\,
            lcout => \U712_CHIP_RAM.N_376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_3_1_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100111001101"
        )
    port map (
            in0 => \N__6166\,
            in1 => \N__5088\,
            in2 => \N__5446\,
            in3 => \N__6024\,
            lcout => \U712_CHIP_RAM.N_378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIGB4P1_3_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__6021\,
            in1 => \N__6163\,
            in2 => \N__10418\,
            in3 => \N__5502\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m101_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI7AC23_0_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110101"
        )
    port map (
            in0 => \N__6164\,
            in1 => \N__6023\,
            in2 => \N__4581\,
            in3 => \N__5087\,
            lcout => \U712_CHIP_RAM.m101_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001111"
        )
    port map (
            in0 => \N__5428\,
            in1 => \N__5306\,
            in2 => \N__5544\,
            in3 => \N__6026\,
            lcout => \U712_CHIP_RAM.m123_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5571\,
            in2 => \_gnd_net_\,
            in3 => \N__5089\,
            lcout => \U712_CHIP_RAM.N_304\,
            ltout => \U712_CHIP_RAM.N_304_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNID3LR1_0_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__5090\,
            in1 => \N__6221\,
            in2 => \N__4707\,
            in3 => \N__6025\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_312_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIBB455_0_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011111111"
        )
    port map (
            in0 => \N__5941\,
            in1 => \_gnd_net_\,
            in2 => \N__4704\,
            in3 => \N__10408\,
            lcout => \U712_CHIP_RAM.N_326\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__10407\,
            in1 => \N__5592\,
            in2 => \N__4701\,
            in3 => \N__4689\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9960\,
            ce => \N__4637\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIA8V79_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011111010"
        )
    port map (
            in0 => \N__4662\,
            in1 => \N__6222\,
            in2 => \N__6995\,
            in3 => \N__6027\,
            lcout => \U712_CHIP_RAM.N_39\,
            ltout => \U712_CHIP_RAM.N_39_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__4658\,
            in1 => \N__5034\,
            in2 => \N__4644\,
            in3 => \N__4719\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9960\,
            ce => \N__4637\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__6254\,
            in1 => \N__10393\,
            in2 => \N__5872\,
            in3 => \N__5603\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5230\,
            in1 => \N__4876\,
            in2 => \N__4907\,
            in3 => \N__5266\,
            lcout => \U712_CHIP_RAM.N_307\,
            ltout => \U712_CHIP_RAM.N_307_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5501\,
            in1 => \N__5419\,
            in2 => \N__4728\,
            in3 => \N__5085\,
            lcout => \U712_CHIP_RAM.N_467\,
            ltout => \U712_CHIP_RAM.N_467_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__6212\,
            in1 => \_gnd_net_\,
            in2 => \N__4725\,
            in3 => \N__6028\,
            lcout => \U712_CHIP_RAM.N_476\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU7TF5_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6029\,
            in1 => \N__5816\,
            in2 => \N__6987\,
            in3 => \N__6213\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKHPV5_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4722\,
            in3 => \N__9825\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010000000"
        )
    port map (
            in0 => \N__6030\,
            in1 => \N__6214\,
            in2 => \N__6988\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_440\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6215\,
            in1 => \N__5864\,
            in2 => \N__6093\,
            in3 => \N__6979\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9967\,
            ce => \N__6267\,
            sr => \N__9775\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_2_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4838\,
            in1 => \N__4772\,
            in2 => \N__4860\,
            in3 => \N__4823\,
            lcout => \U712_CHIP_RAM.m93_i_a2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4793\,
            in1 => \N__4808\,
            in2 => \_gnd_net_\,
            in3 => \N__6378\,
            lcout => \U712_CHIP_RAM.m93_i_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_0_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5572\,
            in2 => \_gnd_net_\,
            in3 => \N__5112\,
            lcout => \U712_CHIP_RAM.N_321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000000000"
        )
    port map (
            in0 => \N__7441\,
            in1 => \N__6330\,
            in2 => \N__5876\,
            in3 => \N__10384\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9973\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.un3_DBR_COUNT_cry_1_c_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4858\,
            in2 => \N__5732\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \U712_CHIP_RAM.un3_DBR_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBR_COUNT_2_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4839\,
            in2 => \_gnd_net_\,
            in3 => \N__4827\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un3_DBR_COUNT_cry_1\,
            carryout => \U712_CHIP_RAM.un3_DBR_COUNT_cry_2\,
            clk => \N__9978\,
            ce => 'H',
            sr => \N__6362\
        );

    \U712_CHIP_RAM.DBR_COUNT_3_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4824\,
            in2 => \_gnd_net_\,
            in3 => \N__4812\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un3_DBR_COUNT_cry_2\,
            carryout => \U712_CHIP_RAM.un3_DBR_COUNT_cry_3\,
            clk => \N__9978\,
            ce => 'H',
            sr => \N__6362\
        );

    \U712_CHIP_RAM.DBR_COUNT_4_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4809\,
            in2 => \_gnd_net_\,
            in3 => \N__4797\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un3_DBR_COUNT_cry_3\,
            carryout => \U712_CHIP_RAM.un3_DBR_COUNT_cry_4\,
            clk => \N__9978\,
            ce => 'H',
            sr => \N__6362\
        );

    \U712_CHIP_RAM.DBR_COUNT_5_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4794\,
            in2 => \_gnd_net_\,
            in3 => \N__4782\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un3_DBR_COUNT_cry_4\,
            carryout => \U712_CHIP_RAM.un3_DBR_COUNT_cry_5\,
            clk => \N__9978\,
            ce => 'H',
            sr => \N__6362\
        );

    \U712_CHIP_RAM.DBR_COUNT_6_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5757\,
            in2 => \_gnd_net_\,
            in3 => \N__4779\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un3_DBR_COUNT_cry_5\,
            carryout => \U712_CHIP_RAM.un3_DBR_COUNT_cry_6\,
            clk => \N__9978\,
            ce => 'H',
            sr => \N__6362\
        );

    \U712_CHIP_RAM.DBR_COUNT_7_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4773\,
            in2 => \_gnd_net_\,
            in3 => \N__4776\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9978\,
            ce => 'H',
            sr => \N__6362\
        );

    \DBR_SYNC_0_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4760\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9987\,
            ce => 'H',
            sr => \N__9755\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5007\,
            in1 => \N__4989\,
            in2 => \_gnd_net_\,
            in3 => \N__8332\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8333\,
            in1 => \N__10947\,
            in2 => \N__4983\,
            in3 => \N__9123\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4980\,
            in1 => \N__4962\,
            in2 => \_gnd_net_\,
            in3 => \N__8331\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_0_a2_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__10948\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11897\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111101110"
        )
    port map (
            in0 => \N__4917\,
            in1 => \N__5213\,
            in2 => \N__5313\,
            in3 => \N__6220\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMDsr_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101111001000"
        )
    port map (
            in0 => \N__4938\,
            in1 => \N__4931\,
            in2 => \N__4920\,
            in3 => \N__6631\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9944\,
            ce => 'H',
            sr => \N__9791\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__5546\,
            in1 => \N__5245\,
            in2 => \_gnd_net_\,
            in3 => \N__5278\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6ORT_7_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4911\,
            in2 => \_gnd_net_\,
            in3 => \N__4884\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDs_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_2_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011110"
        )
    port map (
            in0 => \N__6098\,
            in1 => \N__5246\,
            in2 => \N__5121\,
            in3 => \N__5279\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMDsr_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_2_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__5212\,
            in1 => \N__5547\,
            in2 => \N__5289\,
            in3 => \N__5120\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_1_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5286\,
            in1 => \N__5280\,
            in2 => \N__5250\,
            in3 => \N__5214\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_1_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000100"
        )
    port map (
            in0 => \N__6062\,
            in1 => \N__6209\,
            in2 => \N__6315\,
            in3 => \N__5451\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_396_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_1_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5159\,
            in1 => \N__5193\,
            in2 => \N__5202\,
            in3 => \N__5199\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9947\,
            ce => \N__5139\,
            sr => \N__9785\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_1_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__6060\,
            in1 => \N__5548\,
            in2 => \N__6223\,
            in3 => \N__5877\,
            lcout => \U712_CHIP_RAM.N_397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_2_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5187\,
            in1 => \N__5175\,
            in2 => \N__5163\,
            in3 => \N__5145\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9947\,
            ce => \N__5139\,
            sr => \N__9785\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6061\,
            in1 => \N__5946\,
            in2 => \N__6224\,
            in3 => \N__5111\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7364\,
            in2 => \_gnd_net_\,
            in3 => \N__5110\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__7787\,
            in1 => \N__9099\,
            in2 => \N__7757\,
            in3 => \N__7053\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9955\,
            ce => \N__7654\,
            sr => \N__9776\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__7788\,
            in1 => \N__9090\,
            in2 => \N__7758\,
            in3 => \N__6681\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9955\,
            ce => \N__7654\,
            sr => \N__9776\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__5685\,
            in1 => \N__5676\,
            in2 => \N__10945\,
            in3 => \N__9234\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9955\,
            ce => \N__7654\,
            sr => \N__9776\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__5640\,
            in1 => \N__6216\,
            in2 => \N__5634\,
            in3 => \N__5348\,
            lcout => \U712_CHIP_RAM.N_190\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__5859\,
            in1 => \N__6932\,
            in2 => \_gnd_net_\,
            in3 => \N__11258\,
            lcout => \U712_CHIP_RAM.N_344\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIB0JV5_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__5607\,
            in1 => \N__5817\,
            in2 => \_gnd_net_\,
            in3 => \N__5860\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__10385\,
            in1 => \N__5586\,
            in2 => \N__5580\,
            in3 => \N__5576\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9961\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_3_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__5545\,
            in1 => \N__5450\,
            in2 => \_gnd_net_\,
            in3 => \N__5339\,
            lcout => \U712_CHIP_RAM.N_551\,
            ltout => \U712_CHIP_RAM.N_551_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOBA64_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6050\,
            in1 => \N__6211\,
            in2 => \N__5316\,
            in3 => \N__5305\,
            lcout => \U712_CHIP_RAM.N_435\,
            ltout => \U712_CHIP_RAM.N_435_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI41RO8_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6273\,
            in3 => \N__6883\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9824\,
            in1 => \_gnd_net_\,
            in2 => \N__6270\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6210\,
            in1 => \N__5858\,
            in2 => \N__6986\,
            in3 => \N__6049\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000101"
        )
    port map (
            in0 => \N__7192\,
            in1 => \_gnd_net_\,
            in2 => \N__6311\,
            in3 => \N__6376\,
            lcout => \U712_CHIP_RAM.N_325\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6239\,
            in1 => \N__6225\,
            in2 => \N__6099\,
            in3 => \N__5945\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__10404\,
            in1 => \N__5888\,
            in2 => \N__5925\,
            in3 => \N__5922\,
            lcout => \RAMENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9968\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6377\,
            in1 => \N__6307\,
            in2 => \N__7200\,
            in3 => \N__5857\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5792\,
            in1 => \N__5766\,
            in2 => \_gnd_net_\,
            in3 => \N__8358\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__5756\,
            in1 => \N__5745\,
            in2 => \N__5739\,
            in3 => \N__5706\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_428_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__10405\,
            in1 => \N__8997\,
            in2 => \N__6381\,
            in3 => \N__6291\,
            lcout => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9968\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_3_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10381\,
            in2 => \_gnd_net_\,
            in3 => \N__9021\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9974\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__10380\,
            in1 => \N__8996\,
            in2 => \_gnd_net_\,
            in3 => \N__6287\,
            lcout => \U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_4_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6339\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10382\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9974\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__6345\,
            in1 => \N__6338\,
            in2 => \_gnd_net_\,
            in3 => \N__6286\,
            lcout => \U712_CHIP_RAM.N_430\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__7136\,
            in1 => \N__7151\,
            in2 => \N__7122\,
            in3 => \N__7166\,
            lcout => \U712_CHIP_RAM.REFRESH5lt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7523\,
            in2 => \_gnd_net_\,
            in3 => \N__7103\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.REFRESH5lto7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001010"
        )
    port map (
            in0 => \N__10383\,
            in1 => \N__7505\,
            in2 => \N__6324\,
            in3 => \N__6321\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9974\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10253\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6516\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9979\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNIFFA4_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7415\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7448\,
            lcout => \U712_CHIP_RAM.m50_i_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__11122\,
            in1 => \N__10252\,
            in2 => \_gnd_net_\,
            in3 => \N__11055\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9979\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_1_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6510\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9983\,
            ce => 'H',
            sr => \N__9754\
        );

    \U712_CHIP_RAM.m37_i_o2_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010111011"
        )
    port map (
            in0 => \N__11688\,
            in1 => \N__11497\,
            in2 => \N__11601\,
            in3 => \N__11358\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_335_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNIVU9S_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__11051\,
            in1 => \N__11747\,
            in2 => \N__6504\,
            in3 => \N__10952\,
            lcout => \N_202_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6482\,
            in2 => \_gnd_net_\,
            in3 => \N__6459\,
            lcout => \U712_CHIP_RAM.N_419\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.N_165_i_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__11127\,
            in1 => \N__11044\,
            in2 => \_gnd_net_\,
            in3 => \N__11174\,
            lcout => \N_165_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WEn_LC_10_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6633\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9937\,
            ce => 'H',
            sr => \N__9801\
        );

    \U712_CHIP_RAM.RASn_LC_10_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6597\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9938\,
            ce => 'H',
            sr => \N__9795\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_10_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__7798\,
            in1 => \N__7830\,
            in2 => \N__7754\,
            in3 => \N__6675\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9940\,
            ce => \N__7650\,
            sr => \N__9792\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110001111"
        )
    port map (
            in0 => \N__10949\,
            in1 => \N__7719\,
            in2 => \N__8330\,
            in3 => \N__8202\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6648\,
            in1 => \N__10950\,
            in2 => \_gnd_net_\,
            in3 => \N__9111\,
            lcout => \U712_CHIP_RAM.N_361\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIE8IL_0_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6626\,
            in2 => \_gnd_net_\,
            in3 => \N__6589\,
            lcout => \U712_CHIP_RAM.N_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIUI4B1_0_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6587\,
            in1 => \N__8284\,
            in2 => \N__6632\,
            in3 => \N__7905\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => \U712_CHIP_RAM.REFRESH_RST_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIB72G2_3_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__8285\,
            in1 => \N__7906\,
            in2 => \N__6600\,
            in3 => \N__6588\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_CMA25_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI1HUV2_3_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6567\,
            in3 => \N__9826\,
            lcout => \U712_CHIP_RAM.un1_CMA25_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8286\,
            in1 => \N__6564\,
            in2 => \_gnd_net_\,
            in3 => \N__6531\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__8211\,
            in1 => \N__10951\,
            in2 => \N__6519\,
            in3 => \N__8290\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__7721\,
            in1 => \N__6843\,
            in2 => \N__8368\,
            in3 => \N__7221\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9945\,
            ce => \N__7656\,
            sr => \N__9777\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100000101"
        )
    port map (
            in0 => \N__7720\,
            in1 => \N__10909\,
            in2 => \N__8367\,
            in3 => \N__8198\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6797\,
            in1 => \N__6777\,
            in2 => \_gnd_net_\,
            in3 => \N__8353\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8354\,
            in1 => \N__10910\,
            in2 => \N__6765\,
            in3 => \N__8748\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6762\,
            in2 => \N__6756\,
            in3 => \N__6753\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9945\,
            ce => \N__7656\,
            sr => \N__9777\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__10888\,
            in1 => \N__6729\,
            in2 => \N__8338\,
            in3 => \N__9447\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6720\,
            in1 => \N__7569\,
            in2 => \_gnd_net_\,
            in3 => \N__8304\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__7031\,
            in1 => \N__8313\,
            in2 => \_gnd_net_\,
            in3 => \N__6702\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8315\,
            in1 => \N__10889\,
            in2 => \N__6684\,
            in3 => \N__8595\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011000000"
        )
    port map (
            in0 => \N__6925\,
            in1 => \N__11155\,
            in2 => \N__10406\,
            in3 => \N__6885\,
            lcout => \DMA_WRITE_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7089\,
            in1 => \N__7068\,
            in2 => \_gnd_net_\,
            in3 => \N__8306\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__10887\,
            in1 => \N__8314\,
            in2 => \N__7056\,
            in3 => \N__8736\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNII0RI_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10886\,
            in2 => \_gnd_net_\,
            in3 => \N__8305\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__7020\,
            in1 => \N__7047\,
            in2 => \N__10743\,
            in3 => \N__7032\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9956\,
            ce => 'H',
            sr => \N__9762\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__10896\,
            in1 => \N__7019\,
            in2 => \_gnd_net_\,
            in3 => \N__7008\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9956\,
            ce => 'H',
            sr => \N__9762\
        );

    \U712_CHIP_RAM.DBENn_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100111011101110"
        )
    port map (
            in0 => \N__7002\,
            in1 => \N__7404\,
            in2 => \N__6996\,
            in3 => \N__6945\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9956\,
            ce => 'H',
            sr => \N__9762\
        );

    \U712_CHIP_RAM.DBDIR_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__6854\,
            in1 => \N__6933\,
            in2 => \_gnd_net_\,
            in3 => \N__6884\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9956\,
            ce => 'H',
            sr => \N__9762\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110011110100"
        )
    port map (
            in0 => \N__8648\,
            in1 => \N__7245\,
            in2 => \N__7965\,
            in3 => \N__8574\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9956\,
            ce => 'H',
            sr => \N__9762\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7230\,
            in1 => \N__10891\,
            in2 => \_gnd_net_\,
            in3 => \N__9030\,
            lcout => \U712_CHIP_RAM.N_367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000010100000"
        )
    port map (
            in0 => \N__7212\,
            in1 => \N__10892\,
            in2 => \N__10417\,
            in3 => \N__7196\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9962\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7176\,
            in2 => \_gnd_net_\,
            in3 => \N__7170\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_10_10_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__7488\,
            ce => 'H',
            sr => \N__7461\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7167\,
            in2 => \_gnd_net_\,
            in3 => \N__7155\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__7488\,
            ce => 'H',
            sr => \N__7461\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7152\,
            in2 => \_gnd_net_\,
            in3 => \N__7140\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__7488\,
            ce => 'H',
            sr => \N__7461\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7137\,
            in2 => \_gnd_net_\,
            in3 => \N__7125\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__7488\,
            ce => 'H',
            sr => \N__7461\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7121\,
            in2 => \_gnd_net_\,
            in3 => \N__7107\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__7488\,
            ce => 'H',
            sr => \N__7461\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7104\,
            in2 => \_gnd_net_\,
            in3 => \N__7092\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__7488\,
            ce => 'H',
            sr => \N__7461\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7524\,
            in2 => \_gnd_net_\,
            in3 => \N__7512\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__7488\,
            ce => 'H',
            sr => \N__7461\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7506\,
            in2 => \_gnd_net_\,
            in3 => \N__7509\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7488\,
            ce => 'H',
            sr => \N__7461\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__7452\,
            in1 => \N__7414\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.START_RST_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__7376\,
            in1 => \N__8086\,
            in2 => \_gnd_net_\,
            in3 => \N__8785\,
            lcout => \U712_REG_SM.START_RSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9980\,
            ce => 'H',
            sr => \N__9750\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000010100000"
        )
    port map (
            in0 => \N__7386\,
            in1 => \N__7377\,
            in2 => \N__10419\,
            in3 => \N__8109\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9984\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_11_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CRCSn_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7913\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9939\,
            ce => 'H',
            sr => \N__9786\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__7799\,
            in1 => \N__9297\,
            in2 => \N__7753\,
            in3 => \N__7314\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9941\,
            ce => \N__7643\,
            sr => \N__9778\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__7914\,
            in1 => \N__8365\,
            in2 => \_gnd_net_\,
            in3 => \N__7736\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9941\,
            ce => \N__7643\,
            sr => \N__9778\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__10932\,
            in1 => \N__7857\,
            in2 => \N__8370\,
            in3 => \N__8178\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__7740\,
            in1 => \N__7800\,
            in2 => \N__7845\,
            in3 => \N__9504\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9941\,
            ce => \N__7643\,
            sr => \N__9778\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9163\,
            in1 => \N__10741\,
            in2 => \_gnd_net_\,
            in3 => \N__9603\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9222\,
            ce => \N__10494\,
            sr => \N__9766\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__7786\,
            in1 => \N__8184\,
            in2 => \N__7755\,
            in3 => \N__7596\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9946\,
            ce => \N__7655\,
            sr => \N__9763\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__7789\,
            in1 => \N__9081\,
            in2 => \N__7756\,
            in3 => \N__7677\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9946\,
            ce => \N__7655\,
            sr => \N__9763\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__10890\,
            in1 => \N__7602\,
            in2 => \N__8369\,
            in3 => \N__10515\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7590\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9949\,
            ce => \N__7563\,
            sr => \N__9759\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001000100010"
        )
    port map (
            in0 => \N__7985\,
            in1 => \N__8641\,
            in2 => \N__7932\,
            in3 => \N__8727\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9957\,
            ce => 'H',
            sr => \N__9756\
        );

    \U712_CYCLE_TERM.TACK_EN_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011111111"
        )
    port map (
            in0 => \N__7989\,
            in1 => \N__8004\,
            in2 => \_gnd_net_\,
            in3 => \N__8721\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9957\,
            ce => 'H',
            sr => \N__9756\
        );

    \U712_REG_SM.REG_TACK_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__8066\,
            in1 => \N__8688\,
            in2 => \N__7923\,
            in3 => \N__7971\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9957\,
            ce => 'H',
            sr => \N__9756\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__10396\,
            in1 => \_gnd_net_\,
            in2 => \N__7961\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__8883\,
            in1 => \N__8836\,
            in2 => \_gnd_net_\,
            in3 => \N__10097\,
            lcout => \U712_REG_SM.N_373\,
            ltout => \U712_REG_SM.N_373_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8132\,
            in2 => \N__7974\,
            in3 => \N__8912\,
            lcout => \U712_REG_SM.N_130\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10395\,
            in2 => \_gnd_net_\,
            in3 => \N__7941\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__10394\,
            in1 => \N__8573\,
            in2 => \_gnd_net_\,
            in3 => \N__8649\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7954\,
            in2 => \_gnd_net_\,
            in3 => \N__7940\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__8913\,
            in1 => \N__8837\,
            in2 => \_gnd_net_\,
            in3 => \N__10098\,
            lcout => \U712_REG_SM.N_406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_0_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8153\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9969\,
            ce => 'H',
            sr => \N__9751\
        );

    \U712_REG_SM.WRITE_CYCLE_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__11234\,
            in1 => \N__8133\,
            in2 => \_gnd_net_\,
            in3 => \N__8088\,
            lcout => \U712_REG_SM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9969\,
            ce => 'H',
            sr => \N__9751\
        );

    \U712_REG_SM.C3_SYNC_1_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8121\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9969\,
            ce => 'H',
            sr => \N__9751\
        );

    \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8949\,
            in2 => \_gnd_net_\,
            in3 => \N__8777\,
            lcout => \U712_REG_SM.N_328\,
            ltout => \U712_REG_SM.N_328_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8108\,
            in1 => \N__8914\,
            in2 => \N__8115\,
            in3 => \N__8882\,
            lcout => \U712_REG_SM.N_412\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8844\,
            in2 => \_gnd_net_\,
            in3 => \N__10101\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_331_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__8778\,
            in1 => \N__10400\,
            in2 => \N__8112\,
            in3 => \N__8087\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9975\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_RNO_0_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001100010"
        )
    port map (
            in0 => \N__8846\,
            in1 => \N__8393\,
            in2 => \N__8786\,
            in3 => \N__8107\,
            lcout => \U712_REG_SM.REGENn_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8847\,
            in1 => \N__8106\,
            in2 => \N__10104\,
            in3 => \N__8414\,
            lcout => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__8928\,
            in1 => \N__8922\,
            in2 => \N__8067\,
            in3 => \N__8475\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9981\,
            ce => 'H',
            sr => \N__9745\
        );

    \U712_REG_SM.C1_SYNC_0_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8469\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9985\,
            ce => 'H',
            sr => \N__9744\
        );

    \U712_REG_SM.C1_SYNC_1_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8433\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9985\,
            ce => 'H',
            sr => \N__9744\
        );

    \U712_REG_SM.REGENn_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100011011000100"
        )
    port map (
            in0 => \N__8427\,
            in1 => \N__8389\,
            in2 => \N__10113\,
            in3 => \N__8418\,
            lcout => \REGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9988\,
            ce => 'H',
            sr => \N__9743\
        );

    \U712_CHIP_RAM.CASn_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8366\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9936\,
            ce => 'H',
            sr => \N__9773\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9544\,
            in1 => \N__10733\,
            in2 => \_gnd_net_\,
            in3 => \N__9350\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__10499\,
            sr => \N__9765\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9552\,
            in1 => \N__10729\,
            in2 => \_gnd_net_\,
            in3 => \N__9351\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9221\,
            ce => \N__10497\,
            sr => \N__9761\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__9171\,
            in1 => \_gnd_net_\,
            in2 => \N__10742\,
            in3 => \N__10797\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9221\,
            ce => \N__10497\,
            sr => \N__9761\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9602\,
            in1 => \N__10721\,
            in2 => \_gnd_net_\,
            in3 => \N__9154\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__10495\,
            sr => \N__9758\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9551\,
            in1 => \N__10720\,
            in2 => \_gnd_net_\,
            in3 => \N__9601\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__10495\,
            sr => \N__9758\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9069\,
            in1 => \N__10722\,
            in2 => \_gnd_net_\,
            in3 => \N__9495\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__10495\,
            sr => \N__9758\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__8685\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8713\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__8714\,
            in1 => \N__8686\,
            in2 => \_gnd_net_\,
            in3 => \N__8665\,
            lcout => \U712_CYCLE_TERM.N_332\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011111"
        )
    port map (
            in0 => \N__8715\,
            in1 => \N__8687\,
            in2 => \N__8670\,
            in3 => \N__8640\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_455_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__8666\,
            in1 => \N__10318\,
            in2 => \N__8652\,
            in3 => \N__8568\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__8619\,
            in1 => \N__10736\,
            in2 => \N__8594\,
            in3 => \N__9282\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            ce => 'H',
            sr => \N__9753\
        );

    \pll_RNI8MQ3_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8569\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000100"
        )
    port map (
            in0 => \N__9003\,
            in1 => \N__10232\,
            in2 => \N__8853\,
            in3 => \N__10103\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9958\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011011000"
        )
    port map (
            in0 => \N__10231\,
            in1 => \N__8961\,
            in2 => \N__11884\,
            in3 => \N__9012\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9958\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8993\,
            in2 => \_gnd_net_\,
            in3 => \N__8843\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_330_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000100010"
        )
    port map (
            in0 => \N__10325\,
            in1 => \N__8934\,
            in2 => \N__9006\,
            in3 => \N__10102\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9965\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__8911\,
            in1 => \N__8841\,
            in2 => \N__8955\,
            in3 => \N__8994\,
            lcout => \U712_REG_SM.N_413\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_0_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10100\,
            in1 => \N__8995\,
            in2 => \N__8852\,
            in3 => \N__8953\,
            lcout => \U712_REG_SM.N_410\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000101"
        )
    port map (
            in0 => \N__8954\,
            in1 => \N__8842\,
            in2 => \N__8787\,
            in3 => \N__10099\,
            lcout => \U712_REG_SM.STATE_COUNTc_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__8881\,
            in1 => \N__10065\,
            in2 => \_gnd_net_\,
            in3 => \N__8848\,
            lcout => \U712_REG_SM.N_308\,
            ltout => \U712_REG_SM.N_308_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__8877\,
            in1 => \N__8921\,
            in2 => \N__8886\,
            in3 => \N__10326\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9971\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIVCF31_4_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011011111"
        )
    port map (
            in0 => \N__8876\,
            in1 => \N__8845\,
            in2 => \N__10096\,
            in3 => \N__8776\,
            lcout => \U712_REG_SM.un1_REGENn_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10327\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9349\,
            in1 => \N__10735\,
            in2 => \_gnd_net_\,
            in3 => \N__9396\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10503\,
            sr => \N__9779\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9170\,
            in1 => \N__10734\,
            in2 => \_gnd_net_\,
            in3 => \N__10796\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            ce => \N__10500\,
            sr => \N__9767\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10557\,
            in1 => \N__10715\,
            in2 => \_gnd_net_\,
            in3 => \N__10795\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9218\,
            ce => \N__10498\,
            sr => \N__9764\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10558\,
            in1 => \N__10716\,
            in2 => \_gnd_net_\,
            in3 => \N__9068\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9218\,
            ce => \N__10498\,
            sr => \N__9764\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__9494\,
            in1 => \_gnd_net_\,
            in2 => \N__10737\,
            in3 => \N__9288\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9218\,
            ce => \N__10498\,
            sr => \N__9764\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9493\,
            in1 => \N__10702\,
            in2 => \_gnd_net_\,
            in3 => \N__9067\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9217\,
            ce => \N__10496\,
            sr => \N__9760\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10560\,
            in1 => \N__10701\,
            in2 => \_gnd_net_\,
            in3 => \N__9066\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__10493\,
            sr => \N__9757\
        );

    \U712_CHIP_RAM.RAS_SYNC_2_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10317\,
            in2 => \_gnd_net_\,
            in3 => \N__10179\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9964\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_RNO_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9823\,
            in2 => \_gnd_net_\,
            in3 => \N__10127\,
            lcout => \U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9589\,
            in1 => \N__10714\,
            in2 => \_gnd_net_\,
            in3 => \N__9543\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9220\,
            ce => \N__10505\,
            sr => \N__9787\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9287\,
            in1 => \N__10642\,
            in2 => \_gnd_net_\,
            in3 => \N__9483\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__10501\,
            sr => \N__9768\
        );

    \U712_REG_SM.ASn_ess_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10116\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9986\,
            ce => \N__9414\,
            sr => \N__9749\
        );

    \U712_REG_SM.UDSn_RNO_0_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__11467\,
            in1 => \N__11602\,
            in2 => \N__11400\,
            in3 => \N__11250\,
            lcout => \U712_REG_SM.N_459\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.N_336_i_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001011001000"
        )
    port map (
            in0 => \N__11689\,
            in1 => \N__11466\,
            in2 => \N__11617\,
            in3 => \N__11343\,
            lcout => \N_336_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9392\,
            in1 => \N__9339\,
            in2 => \_gnd_net_\,
            in3 => \N__10713\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9219\,
            ce => \N__10506\,
            sr => \N__9793\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10665\,
            in1 => \N__10445\,
            in2 => \_gnd_net_\,
            in3 => \N__9286\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9216\,
            ce => \N__10504\,
            sr => \N__9780\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10785\,
            in1 => \N__10712\,
            in2 => \_gnd_net_\,
            in3 => \N__10559\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__10502\,
            sr => \N__9769\
        );

    \U712_CHIP_RAM.RAS_SYNC_0_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__10350\,
            in1 => \N__10458\,
            in2 => \_gnd_net_\,
            in3 => \N__10446\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9970\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_1_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10300\,
            in2 => \_gnd_net_\,
            in3 => \N__10185\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9976\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111000001110"
        )
    port map (
            in0 => \N__10114\,
            in1 => \N__9636\,
            in2 => \N__10137\,
            in3 => \N__10154\,
            lcout => \LDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9989\,
            ce => 'H',
            sr => \N__9752\
        );

    \U712_REG_SM.UDSn_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111001111100010"
        )
    port map (
            in0 => \N__10143\,
            in1 => \N__10136\,
            in2 => \N__10010\,
            in3 => \N__10115\,
            lcout => \UDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9989\,
            ce => 'H',
            sr => \N__9752\
        );

    \U712_REG_SM.LDSn_RNO_0_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__11603\,
            in1 => \N__11515\,
            in2 => \N__11259\,
            in3 => \N__11397\,
            lcout => \U712_REG_SM.N_404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.N_335_i_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101110000"
        )
    port map (
            in0 => \N__11690\,
            in1 => \N__11607\,
            in2 => \N__11380\,
            in3 => \N__11498\,
            lcout => \N_335_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.N_337_i_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111010000"
        )
    port map (
            in0 => \N__11691\,
            in1 => \N__11608\,
            in2 => \N__11381\,
            in3 => \N__11499\,
            lcout => \N_337_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_177_i_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111011101"
        )
    port map (
            in0 => \N__11804\,
            in1 => \N__11043\,
            in2 => \N__11820\,
            in3 => \N__10965\,
            lcout => \N_177_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m40_i_o2_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010101001111"
        )
    port map (
            in0 => \N__11705\,
            in1 => \N__11612\,
            in2 => \N__11379\,
            in3 => \N__11517\,
            lcout => \N_334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_175_i_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__11123\,
            in1 => \N__11808\,
            in2 => \N__11766\,
            in3 => \N__10966\,
            lcout => \N_175_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m58_i_o2_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110100110111"
        )
    port map (
            in0 => \N__11616\,
            in1 => \N__11399\,
            in2 => \N__11706\,
            in3 => \N__11482\,
            lcout => \N_336\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m34_i_o2_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111001011101"
        )
    port map (
            in0 => \N__11481\,
            in1 => \N__11701\,
            in2 => \N__11619\,
            in3 => \N__11398\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_337_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNI8LI41_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100010011"
        )
    port map (
            in0 => \N__10973\,
            in1 => \N__11754\,
            in2 => \N__11730\,
            in3 => \N__11110\,
            lcout => \N_200_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.N_334_i_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110100000"
        )
    port map (
            in0 => \N__11692\,
            in1 => \N__11618\,
            in2 => \N__11516\,
            in3 => \N__11368\,
            lcout => \N_334_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001111111"
        )
    port map (
            in0 => \N__11120\,
            in1 => \N__11257\,
            in2 => \N__11020\,
            in3 => \N__11175\,
            lcout => \N_379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.N_167_i_LC_24_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__11121\,
            in1 => \N__11013\,
            in2 => \N__10977\,
            in3 => \N__11898\,
            lcout => \N_167_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

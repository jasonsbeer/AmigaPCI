// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Feb 19 2025 16:48:39

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    CMA,
    SIZ,
    DRA,
    A,
    RAMENn,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    RAMSPACEn,
    WEn,
    REGENn,
    LLBEn,
    DBRn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    output [10:0] CMA;
    input [1:0] SIZ;
    input [9:0] DRA;
    input [20:0] A;
    output RAMENn;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    output LLBEn;
    input DBRn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__11973;
    wire N__11972;
    wire N__11971;
    wire N__11964;
    wire N__11963;
    wire N__11962;
    wire N__11955;
    wire N__11954;
    wire N__11953;
    wire N__11946;
    wire N__11945;
    wire N__11944;
    wire N__11937;
    wire N__11936;
    wire N__11935;
    wire N__11928;
    wire N__11927;
    wire N__11926;
    wire N__11919;
    wire N__11918;
    wire N__11917;
    wire N__11910;
    wire N__11909;
    wire N__11908;
    wire N__11901;
    wire N__11900;
    wire N__11899;
    wire N__11892;
    wire N__11891;
    wire N__11890;
    wire N__11883;
    wire N__11882;
    wire N__11881;
    wire N__11874;
    wire N__11873;
    wire N__11872;
    wire N__11865;
    wire N__11864;
    wire N__11863;
    wire N__11856;
    wire N__11855;
    wire N__11854;
    wire N__11847;
    wire N__11846;
    wire N__11845;
    wire N__11838;
    wire N__11837;
    wire N__11836;
    wire N__11829;
    wire N__11828;
    wire N__11827;
    wire N__11820;
    wire N__11819;
    wire N__11818;
    wire N__11811;
    wire N__11810;
    wire N__11809;
    wire N__11802;
    wire N__11801;
    wire N__11800;
    wire N__11793;
    wire N__11792;
    wire N__11791;
    wire N__11784;
    wire N__11783;
    wire N__11782;
    wire N__11775;
    wire N__11774;
    wire N__11773;
    wire N__11766;
    wire N__11765;
    wire N__11764;
    wire N__11757;
    wire N__11756;
    wire N__11755;
    wire N__11748;
    wire N__11747;
    wire N__11746;
    wire N__11739;
    wire N__11738;
    wire N__11737;
    wire N__11730;
    wire N__11729;
    wire N__11728;
    wire N__11721;
    wire N__11720;
    wire N__11719;
    wire N__11712;
    wire N__11711;
    wire N__11710;
    wire N__11703;
    wire N__11702;
    wire N__11701;
    wire N__11694;
    wire N__11693;
    wire N__11692;
    wire N__11685;
    wire N__11684;
    wire N__11683;
    wire N__11676;
    wire N__11675;
    wire N__11674;
    wire N__11667;
    wire N__11666;
    wire N__11665;
    wire N__11658;
    wire N__11657;
    wire N__11656;
    wire N__11649;
    wire N__11648;
    wire N__11647;
    wire N__11640;
    wire N__11639;
    wire N__11638;
    wire N__11631;
    wire N__11630;
    wire N__11629;
    wire N__11622;
    wire N__11621;
    wire N__11620;
    wire N__11613;
    wire N__11612;
    wire N__11611;
    wire N__11604;
    wire N__11603;
    wire N__11602;
    wire N__11595;
    wire N__11594;
    wire N__11593;
    wire N__11586;
    wire N__11585;
    wire N__11584;
    wire N__11577;
    wire N__11576;
    wire N__11575;
    wire N__11568;
    wire N__11567;
    wire N__11566;
    wire N__11559;
    wire N__11558;
    wire N__11557;
    wire N__11550;
    wire N__11549;
    wire N__11548;
    wire N__11541;
    wire N__11540;
    wire N__11539;
    wire N__11532;
    wire N__11531;
    wire N__11530;
    wire N__11523;
    wire N__11522;
    wire N__11521;
    wire N__11514;
    wire N__11513;
    wire N__11512;
    wire N__11505;
    wire N__11504;
    wire N__11503;
    wire N__11496;
    wire N__11495;
    wire N__11494;
    wire N__11487;
    wire N__11486;
    wire N__11485;
    wire N__11478;
    wire N__11477;
    wire N__11476;
    wire N__11469;
    wire N__11468;
    wire N__11467;
    wire N__11460;
    wire N__11459;
    wire N__11458;
    wire N__11451;
    wire N__11450;
    wire N__11449;
    wire N__11442;
    wire N__11441;
    wire N__11440;
    wire N__11433;
    wire N__11432;
    wire N__11431;
    wire N__11424;
    wire N__11423;
    wire N__11422;
    wire N__11415;
    wire N__11414;
    wire N__11413;
    wire N__11406;
    wire N__11405;
    wire N__11404;
    wire N__11397;
    wire N__11396;
    wire N__11395;
    wire N__11388;
    wire N__11387;
    wire N__11386;
    wire N__11379;
    wire N__11378;
    wire N__11377;
    wire N__11370;
    wire N__11369;
    wire N__11368;
    wire N__11361;
    wire N__11360;
    wire N__11359;
    wire N__11352;
    wire N__11351;
    wire N__11350;
    wire N__11343;
    wire N__11342;
    wire N__11341;
    wire N__11334;
    wire N__11333;
    wire N__11332;
    wire N__11325;
    wire N__11324;
    wire N__11323;
    wire N__11316;
    wire N__11315;
    wire N__11314;
    wire N__11307;
    wire N__11306;
    wire N__11305;
    wire N__11298;
    wire N__11297;
    wire N__11296;
    wire N__11289;
    wire N__11288;
    wire N__11287;
    wire N__11280;
    wire N__11279;
    wire N__11278;
    wire N__11271;
    wire N__11270;
    wire N__11269;
    wire N__11262;
    wire N__11261;
    wire N__11260;
    wire N__11253;
    wire N__11252;
    wire N__11251;
    wire N__11244;
    wire N__11243;
    wire N__11242;
    wire N__11235;
    wire N__11234;
    wire N__11233;
    wire N__11226;
    wire N__11225;
    wire N__11224;
    wire N__11217;
    wire N__11216;
    wire N__11215;
    wire N__11208;
    wire N__11207;
    wire N__11206;
    wire N__11199;
    wire N__11198;
    wire N__11197;
    wire N__11190;
    wire N__11189;
    wire N__11188;
    wire N__11181;
    wire N__11180;
    wire N__11179;
    wire N__11172;
    wire N__11171;
    wire N__11170;
    wire N__11153;
    wire N__11152;
    wire N__11149;
    wire N__11146;
    wire N__11145;
    wire N__11142;
    wire N__11139;
    wire N__11136;
    wire N__11133;
    wire N__11128;
    wire N__11127;
    wire N__11124;
    wire N__11121;
    wire N__11118;
    wire N__11115;
    wire N__11112;
    wire N__11109;
    wire N__11106;
    wire N__11103;
    wire N__11100;
    wire N__11097;
    wire N__11094;
    wire N__11091;
    wire N__11084;
    wire N__11081;
    wire N__11078;
    wire N__11075;
    wire N__11072;
    wire N__11071;
    wire N__11070;
    wire N__11069;
    wire N__11066;
    wire N__11063;
    wire N__11062;
    wire N__11061;
    wire N__11060;
    wire N__11059;
    wire N__11056;
    wire N__11055;
    wire N__11054;
    wire N__11053;
    wire N__11050;
    wire N__11049;
    wire N__11048;
    wire N__11043;
    wire N__11038;
    wire N__11033;
    wire N__11032;
    wire N__11025;
    wire N__11022;
    wire N__11017;
    wire N__11016;
    wire N__11013;
    wire N__11012;
    wire N__11007;
    wire N__11004;
    wire N__11003;
    wire N__11002;
    wire N__11001;
    wire N__11000;
    wire N__10997;
    wire N__10996;
    wire N__10993;
    wire N__10988;
    wire N__10985;
    wire N__10982;
    wire N__10979;
    wire N__10974;
    wire N__10969;
    wire N__10964;
    wire N__10959;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10937;
    wire N__10934;
    wire N__10931;
    wire N__10928;
    wire N__10925;
    wire N__10922;
    wire N__10919;
    wire N__10914;
    wire N__10911;
    wire N__10908;
    wire N__10901;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10888;
    wire N__10887;
    wire N__10886;
    wire N__10885;
    wire N__10884;
    wire N__10883;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10861;
    wire N__10860;
    wire N__10859;
    wire N__10858;
    wire N__10857;
    wire N__10856;
    wire N__10855;
    wire N__10854;
    wire N__10853;
    wire N__10832;
    wire N__10829;
    wire N__10826;
    wire N__10825;
    wire N__10824;
    wire N__10823;
    wire N__10822;
    wire N__10817;
    wire N__10814;
    wire N__10811;
    wire N__10808;
    wire N__10807;
    wire N__10806;
    wire N__10805;
    wire N__10804;
    wire N__10803;
    wire N__10802;
    wire N__10801;
    wire N__10800;
    wire N__10797;
    wire N__10796;
    wire N__10795;
    wire N__10794;
    wire N__10793;
    wire N__10790;
    wire N__10789;
    wire N__10788;
    wire N__10787;
    wire N__10786;
    wire N__10785;
    wire N__10784;
    wire N__10783;
    wire N__10782;
    wire N__10781;
    wire N__10780;
    wire N__10779;
    wire N__10778;
    wire N__10777;
    wire N__10776;
    wire N__10775;
    wire N__10772;
    wire N__10771;
    wire N__10770;
    wire N__10769;
    wire N__10768;
    wire N__10767;
    wire N__10766;
    wire N__10763;
    wire N__10762;
    wire N__10761;
    wire N__10760;
    wire N__10759;
    wire N__10758;
    wire N__10757;
    wire N__10670;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10655;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10637;
    wire N__10634;
    wire N__10631;
    wire N__10628;
    wire N__10625;
    wire N__10622;
    wire N__10619;
    wire N__10616;
    wire N__10613;
    wire N__10610;
    wire N__10609;
    wire N__10608;
    wire N__10607;
    wire N__10604;
    wire N__10599;
    wire N__10596;
    wire N__10589;
    wire N__10586;
    wire N__10583;
    wire N__10580;
    wire N__10577;
    wire N__10576;
    wire N__10575;
    wire N__10572;
    wire N__10569;
    wire N__10568;
    wire N__10565;
    wire N__10560;
    wire N__10557;
    wire N__10554;
    wire N__10551;
    wire N__10548;
    wire N__10545;
    wire N__10542;
    wire N__10539;
    wire N__10536;
    wire N__10533;
    wire N__10530;
    wire N__10527;
    wire N__10520;
    wire N__10519;
    wire N__10514;
    wire N__10511;
    wire N__10508;
    wire N__10505;
    wire N__10502;
    wire N__10501;
    wire N__10500;
    wire N__10499;
    wire N__10496;
    wire N__10491;
    wire N__10488;
    wire N__10485;
    wire N__10480;
    wire N__10475;
    wire N__10472;
    wire N__10469;
    wire N__10466;
    wire N__10465;
    wire N__10464;
    wire N__10461;
    wire N__10458;
    wire N__10455;
    wire N__10454;
    wire N__10449;
    wire N__10446;
    wire N__10443;
    wire N__10440;
    wire N__10437;
    wire N__10434;
    wire N__10431;
    wire N__10428;
    wire N__10425;
    wire N__10422;
    wire N__10419;
    wire N__10416;
    wire N__10413;
    wire N__10408;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10376;
    wire N__10375;
    wire N__10372;
    wire N__10369;
    wire N__10366;
    wire N__10361;
    wire N__10358;
    wire N__10357;
    wire N__10354;
    wire N__10351;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10327;
    wire N__10326;
    wire N__10323;
    wire N__10322;
    wire N__10317;
    wire N__10314;
    wire N__10311;
    wire N__10308;
    wire N__10307;
    wire N__10306;
    wire N__10301;
    wire N__10298;
    wire N__10295;
    wire N__10292;
    wire N__10291;
    wire N__10288;
    wire N__10285;
    wire N__10280;
    wire N__10277;
    wire N__10276;
    wire N__10273;
    wire N__10268;
    wire N__10265;
    wire N__10262;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10246;
    wire N__10245;
    wire N__10244;
    wire N__10243;
    wire N__10242;
    wire N__10241;
    wire N__10240;
    wire N__10237;
    wire N__10236;
    wire N__10233;
    wire N__10230;
    wire N__10227;
    wire N__10222;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10202;
    wire N__10193;
    wire N__10190;
    wire N__10185;
    wire N__10182;
    wire N__10179;
    wire N__10176;
    wire N__10173;
    wire N__10170;
    wire N__10167;
    wire N__10160;
    wire N__10157;
    wire N__10156;
    wire N__10155;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10147;
    wire N__10144;
    wire N__10143;
    wire N__10140;
    wire N__10139;
    wire N__10134;
    wire N__10131;
    wire N__10128;
    wire N__10123;
    wire N__10122;
    wire N__10121;
    wire N__10118;
    wire N__10115;
    wire N__10110;
    wire N__10107;
    wire N__10102;
    wire N__10099;
    wire N__10096;
    wire N__10089;
    wire N__10086;
    wire N__10081;
    wire N__10078;
    wire N__10075;
    wire N__10072;
    wire N__10069;
    wire N__10064;
    wire N__10061;
    wire N__10060;
    wire N__10059;
    wire N__10056;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10048;
    wire N__10045;
    wire N__10042;
    wire N__10039;
    wire N__10036;
    wire N__10035;
    wire N__10032;
    wire N__10027;
    wire N__10024;
    wire N__10021;
    wire N__10018;
    wire N__10015;
    wire N__10012;
    wire N__10009;
    wire N__10006;
    wire N__10001;
    wire N__9998;
    wire N__9991;
    wire N__9988;
    wire N__9985;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9967;
    wire N__9964;
    wire N__9963;
    wire N__9960;
    wire N__9959;
    wire N__9958;
    wire N__9955;
    wire N__9952;
    wire N__9949;
    wire N__9944;
    wire N__9939;
    wire N__9934;
    wire N__9933;
    wire N__9930;
    wire N__9927;
    wire N__9924;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9895;
    wire N__9894;
    wire N__9893;
    wire N__9890;
    wire N__9889;
    wire N__9886;
    wire N__9883;
    wire N__9880;
    wire N__9877;
    wire N__9872;
    wire N__9869;
    wire N__9866;
    wire N__9861;
    wire N__9860;
    wire N__9855;
    wire N__9852;
    wire N__9849;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9830;
    wire N__9827;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9817;
    wire N__9816;
    wire N__9815;
    wire N__9814;
    wire N__9813;
    wire N__9812;
    wire N__9811;
    wire N__9810;
    wire N__9809;
    wire N__9808;
    wire N__9807;
    wire N__9806;
    wire N__9805;
    wire N__9804;
    wire N__9803;
    wire N__9802;
    wire N__9801;
    wire N__9800;
    wire N__9797;
    wire N__9796;
    wire N__9795;
    wire N__9794;
    wire N__9793;
    wire N__9792;
    wire N__9791;
    wire N__9790;
    wire N__9789;
    wire N__9788;
    wire N__9787;
    wire N__9786;
    wire N__9785;
    wire N__9784;
    wire N__9783;
    wire N__9782;
    wire N__9713;
    wire N__9710;
    wire N__9709;
    wire N__9708;
    wire N__9707;
    wire N__9706;
    wire N__9705;
    wire N__9704;
    wire N__9703;
    wire N__9700;
    wire N__9699;
    wire N__9696;
    wire N__9695;
    wire N__9694;
    wire N__9691;
    wire N__9690;
    wire N__9689;
    wire N__9686;
    wire N__9683;
    wire N__9682;
    wire N__9681;
    wire N__9678;
    wire N__9675;
    wire N__9674;
    wire N__9673;
    wire N__9670;
    wire N__9665;
    wire N__9662;
    wire N__9661;
    wire N__9658;
    wire N__9657;
    wire N__9656;
    wire N__9653;
    wire N__9646;
    wire N__9645;
    wire N__9644;
    wire N__9639;
    wire N__9638;
    wire N__9637;
    wire N__9634;
    wire N__9631;
    wire N__9626;
    wire N__9621;
    wire N__9618;
    wire N__9613;
    wire N__9608;
    wire N__9603;
    wire N__9598;
    wire N__9595;
    wire N__9592;
    wire N__9589;
    wire N__9586;
    wire N__9581;
    wire N__9578;
    wire N__9573;
    wire N__9568;
    wire N__9561;
    wire N__9556;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9532;
    wire N__9531;
    wire N__9528;
    wire N__9527;
    wire N__9526;
    wire N__9525;
    wire N__9524;
    wire N__9523;
    wire N__9522;
    wire N__9521;
    wire N__9520;
    wire N__9519;
    wire N__9516;
    wire N__9513;
    wire N__9512;
    wire N__9509;
    wire N__9506;
    wire N__9503;
    wire N__9502;
    wire N__9499;
    wire N__9498;
    wire N__9495;
    wire N__9494;
    wire N__9493;
    wire N__9492;
    wire N__9489;
    wire N__9484;
    wire N__9479;
    wire N__9476;
    wire N__9471;
    wire N__9468;
    wire N__9465;
    wire N__9464;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9448;
    wire N__9443;
    wire N__9442;
    wire N__9437;
    wire N__9432;
    wire N__9427;
    wire N__9424;
    wire N__9421;
    wire N__9420;
    wire N__9419;
    wire N__9418;
    wire N__9417;
    wire N__9406;
    wire N__9403;
    wire N__9400;
    wire N__9397;
    wire N__9394;
    wire N__9389;
    wire N__9382;
    wire N__9379;
    wire N__9374;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9347;
    wire N__9344;
    wire N__9341;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9326;
    wire N__9323;
    wire N__9322;
    wire N__9321;
    wire N__9316;
    wire N__9313;
    wire N__9310;
    wire N__9307;
    wire N__9306;
    wire N__9303;
    wire N__9300;
    wire N__9297;
    wire N__9294;
    wire N__9291;
    wire N__9288;
    wire N__9281;
    wire N__9278;
    wire N__9275;
    wire N__9274;
    wire N__9271;
    wire N__9268;
    wire N__9267;
    wire N__9262;
    wire N__9259;
    wire N__9258;
    wire N__9255;
    wire N__9252;
    wire N__9249;
    wire N__9246;
    wire N__9241;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9223;
    wire N__9220;
    wire N__9217;
    wire N__9216;
    wire N__9211;
    wire N__9208;
    wire N__9207;
    wire N__9204;
    wire N__9201;
    wire N__9198;
    wire N__9193;
    wire N__9190;
    wire N__9187;
    wire N__9184;
    wire N__9179;
    wire N__9176;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9140;
    wire N__9137;
    wire N__9134;
    wire N__9131;
    wire N__9130;
    wire N__9129;
    wire N__9128;
    wire N__9127;
    wire N__9124;
    wire N__9121;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9074;
    wire N__9071;
    wire N__9068;
    wire N__9065;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9040;
    wire N__9039;
    wire N__9036;
    wire N__9033;
    wire N__9030;
    wire N__9027;
    wire N__9026;
    wire N__9019;
    wire N__9016;
    wire N__9011;
    wire N__9008;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8996;
    wire N__8993;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8960;
    wire N__8957;
    wire N__8956;
    wire N__8953;
    wire N__8950;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8921;
    wire N__8918;
    wire N__8915;
    wire N__8912;
    wire N__8909;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8894;
    wire N__8891;
    wire N__8888;
    wire N__8885;
    wire N__8882;
    wire N__8879;
    wire N__8876;
    wire N__8875;
    wire N__8872;
    wire N__8871;
    wire N__8868;
    wire N__8865;
    wire N__8862;
    wire N__8861;
    wire N__8856;
    wire N__8853;
    wire N__8850;
    wire N__8847;
    wire N__8844;
    wire N__8841;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8798;
    wire N__8795;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8783;
    wire N__8782;
    wire N__8781;
    wire N__8778;
    wire N__8775;
    wire N__8772;
    wire N__8771;
    wire N__8770;
    wire N__8767;
    wire N__8766;
    wire N__8763;
    wire N__8760;
    wire N__8759;
    wire N__8758;
    wire N__8757;
    wire N__8752;
    wire N__8749;
    wire N__8746;
    wire N__8743;
    wire N__8740;
    wire N__8733;
    wire N__8720;
    wire N__8719;
    wire N__8718;
    wire N__8717;
    wire N__8716;
    wire N__8715;
    wire N__8712;
    wire N__8707;
    wire N__8704;
    wire N__8699;
    wire N__8690;
    wire N__8687;
    wire N__8684;
    wire N__8681;
    wire N__8678;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8602;
    wire N__8601;
    wire N__8598;
    wire N__8595;
    wire N__8590;
    wire N__8587;
    wire N__8582;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8524;
    wire N__8519;
    wire N__8516;
    wire N__8513;
    wire N__8510;
    wire N__8507;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8482;
    wire N__8481;
    wire N__8478;
    wire N__8475;
    wire N__8474;
    wire N__8467;
    wire N__8464;
    wire N__8461;
    wire N__8458;
    wire N__8455;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8440;
    wire N__8437;
    wire N__8434;
    wire N__8431;
    wire N__8428;
    wire N__8425;
    wire N__8422;
    wire N__8419;
    wire N__8416;
    wire N__8415;
    wire N__8410;
    wire N__8407;
    wire N__8404;
    wire N__8401;
    wire N__8396;
    wire N__8393;
    wire N__8392;
    wire N__8391;
    wire N__8390;
    wire N__8389;
    wire N__8388;
    wire N__8387;
    wire N__8386;
    wire N__8383;
    wire N__8376;
    wire N__8375;
    wire N__8374;
    wire N__8373;
    wire N__8372;
    wire N__8365;
    wire N__8364;
    wire N__8363;
    wire N__8362;
    wire N__8361;
    wire N__8360;
    wire N__8359;
    wire N__8356;
    wire N__8353;
    wire N__8350;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8329;
    wire N__8326;
    wire N__8321;
    wire N__8318;
    wire N__8315;
    wire N__8308;
    wire N__8305;
    wire N__8296;
    wire N__8295;
    wire N__8292;
    wire N__8287;
    wire N__8282;
    wire N__8279;
    wire N__8270;
    wire N__8267;
    wire N__8264;
    wire N__8261;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8251;
    wire N__8250;
    wire N__8245;
    wire N__8242;
    wire N__8241;
    wire N__8236;
    wire N__8233;
    wire N__8232;
    wire N__8229;
    wire N__8226;
    wire N__8223;
    wire N__8216;
    wire N__8215;
    wire N__8212;
    wire N__8209;
    wire N__8206;
    wire N__8203;
    wire N__8198;
    wire N__8195;
    wire N__8192;
    wire N__8191;
    wire N__8190;
    wire N__8189;
    wire N__8184;
    wire N__8181;
    wire N__8178;
    wire N__8173;
    wire N__8172;
    wire N__8171;
    wire N__8168;
    wire N__8165;
    wire N__8160;
    wire N__8157;
    wire N__8154;
    wire N__8151;
    wire N__8148;
    wire N__8145;
    wire N__8142;
    wire N__8139;
    wire N__8134;
    wire N__8131;
    wire N__8126;
    wire N__8125;
    wire N__8124;
    wire N__8121;
    wire N__8118;
    wire N__8115;
    wire N__8112;
    wire N__8109;
    wire N__8106;
    wire N__8103;
    wire N__8100;
    wire N__8097;
    wire N__8094;
    wire N__8091;
    wire N__8088;
    wire N__8085;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8069;
    wire N__8066;
    wire N__8063;
    wire N__8060;
    wire N__8057;
    wire N__8054;
    wire N__8051;
    wire N__8048;
    wire N__8045;
    wire N__8042;
    wire N__8039;
    wire N__8036;
    wire N__8033;
    wire N__8030;
    wire N__8027;
    wire N__8024;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8012;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8000;
    wire N__7997;
    wire N__7994;
    wire N__7991;
    wire N__7988;
    wire N__7985;
    wire N__7982;
    wire N__7979;
    wire N__7976;
    wire N__7973;
    wire N__7972;
    wire N__7971;
    wire N__7970;
    wire N__7969;
    wire N__7968;
    wire N__7967;
    wire N__7966;
    wire N__7965;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7951;
    wire N__7950;
    wire N__7949;
    wire N__7946;
    wire N__7945;
    wire N__7942;
    wire N__7937;
    wire N__7934;
    wire N__7929;
    wire N__7924;
    wire N__7923;
    wire N__7922;
    wire N__7921;
    wire N__7918;
    wire N__7915;
    wire N__7910;
    wire N__7907;
    wire N__7904;
    wire N__7899;
    wire N__7896;
    wire N__7893;
    wire N__7890;
    wire N__7871;
    wire N__7870;
    wire N__7869;
    wire N__7868;
    wire N__7867;
    wire N__7864;
    wire N__7861;
    wire N__7858;
    wire N__7855;
    wire N__7852;
    wire N__7851;
    wire N__7850;
    wire N__7849;
    wire N__7848;
    wire N__7847;
    wire N__7846;
    wire N__7841;
    wire N__7836;
    wire N__7833;
    wire N__7832;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7819;
    wire N__7816;
    wire N__7815;
    wire N__7814;
    wire N__7813;
    wire N__7812;
    wire N__7811;
    wire N__7810;
    wire N__7809;
    wire N__7808;
    wire N__7805;
    wire N__7802;
    wire N__7797;
    wire N__7794;
    wire N__7787;
    wire N__7778;
    wire N__7775;
    wire N__7762;
    wire N__7745;
    wire N__7742;
    wire N__7741;
    wire N__7740;
    wire N__7737;
    wire N__7734;
    wire N__7731;
    wire N__7726;
    wire N__7723;
    wire N__7720;
    wire N__7715;
    wire N__7712;
    wire N__7709;
    wire N__7706;
    wire N__7703;
    wire N__7700;
    wire N__7697;
    wire N__7696;
    wire N__7691;
    wire N__7688;
    wire N__7685;
    wire N__7682;
    wire N__7679;
    wire N__7676;
    wire N__7673;
    wire N__7670;
    wire N__7667;
    wire N__7664;
    wire N__7661;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7639;
    wire N__7634;
    wire N__7631;
    wire N__7628;
    wire N__7625;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7613;
    wire N__7612;
    wire N__7611;
    wire N__7610;
    wire N__7609;
    wire N__7606;
    wire N__7605;
    wire N__7596;
    wire N__7593;
    wire N__7590;
    wire N__7589;
    wire N__7588;
    wire N__7585;
    wire N__7580;
    wire N__7575;
    wire N__7568;
    wire N__7567;
    wire N__7566;
    wire N__7563;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7550;
    wire N__7547;
    wire N__7546;
    wire N__7545;
    wire N__7542;
    wire N__7537;
    wire N__7534;
    wire N__7531;
    wire N__7528;
    wire N__7525;
    wire N__7522;
    wire N__7521;
    wire N__7518;
    wire N__7513;
    wire N__7512;
    wire N__7511;
    wire N__7510;
    wire N__7507;
    wire N__7504;
    wire N__7501;
    wire N__7496;
    wire N__7491;
    wire N__7488;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7468;
    wire N__7465;
    wire N__7462;
    wire N__7457;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7444;
    wire N__7443;
    wire N__7440;
    wire N__7439;
    wire N__7438;
    wire N__7437;
    wire N__7436;
    wire N__7435;
    wire N__7434;
    wire N__7433;
    wire N__7432;
    wire N__7429;
    wire N__7428;
    wire N__7427;
    wire N__7426;
    wire N__7423;
    wire N__7420;
    wire N__7417;
    wire N__7416;
    wire N__7415;
    wire N__7414;
    wire N__7413;
    wire N__7410;
    wire N__7403;
    wire N__7396;
    wire N__7395;
    wire N__7392;
    wire N__7387;
    wire N__7386;
    wire N__7385;
    wire N__7382;
    wire N__7381;
    wire N__7380;
    wire N__7379;
    wire N__7378;
    wire N__7375;
    wire N__7372;
    wire N__7369;
    wire N__7360;
    wire N__7353;
    wire N__7350;
    wire N__7345;
    wire N__7340;
    wire N__7337;
    wire N__7334;
    wire N__7327;
    wire N__7304;
    wire N__7303;
    wire N__7298;
    wire N__7295;
    wire N__7294;
    wire N__7291;
    wire N__7288;
    wire N__7287;
    wire N__7286;
    wire N__7285;
    wire N__7284;
    wire N__7279;
    wire N__7276;
    wire N__7273;
    wire N__7270;
    wire N__7269;
    wire N__7268;
    wire N__7265;
    wire N__7256;
    wire N__7251;
    wire N__7248;
    wire N__7247;
    wire N__7246;
    wire N__7245;
    wire N__7242;
    wire N__7239;
    wire N__7236;
    wire N__7229;
    wire N__7220;
    wire N__7219;
    wire N__7218;
    wire N__7217;
    wire N__7214;
    wire N__7211;
    wire N__7210;
    wire N__7209;
    wire N__7206;
    wire N__7203;
    wire N__7202;
    wire N__7199;
    wire N__7196;
    wire N__7195;
    wire N__7194;
    wire N__7193;
    wire N__7188;
    wire N__7183;
    wire N__7180;
    wire N__7175;
    wire N__7168;
    wire N__7161;
    wire N__7154;
    wire N__7151;
    wire N__7150;
    wire N__7147;
    wire N__7146;
    wire N__7145;
    wire N__7144;
    wire N__7143;
    wire N__7142;
    wire N__7139;
    wire N__7138;
    wire N__7135;
    wire N__7132;
    wire N__7127;
    wire N__7126;
    wire N__7125;
    wire N__7122;
    wire N__7121;
    wire N__7118;
    wire N__7115;
    wire N__7114;
    wire N__7113;
    wire N__7112;
    wire N__7109;
    wire N__7102;
    wire N__7099;
    wire N__7098;
    wire N__7097;
    wire N__7094;
    wire N__7091;
    wire N__7086;
    wire N__7083;
    wire N__7080;
    wire N__7079;
    wire N__7076;
    wire N__7073;
    wire N__7072;
    wire N__7071;
    wire N__7070;
    wire N__7069;
    wire N__7066;
    wire N__7063;
    wire N__7060;
    wire N__7055;
    wire N__7044;
    wire N__7037;
    wire N__7034;
    wire N__7031;
    wire N__7026;
    wire N__7007;
    wire N__7004;
    wire N__7001;
    wire N__7000;
    wire N__6997;
    wire N__6994;
    wire N__6989;
    wire N__6988;
    wire N__6985;
    wire N__6982;
    wire N__6977;
    wire N__6976;
    wire N__6973;
    wire N__6970;
    wire N__6967;
    wire N__6962;
    wire N__6961;
    wire N__6958;
    wire N__6955;
    wire N__6950;
    wire N__6949;
    wire N__6946;
    wire N__6943;
    wire N__6938;
    wire N__6937;
    wire N__6934;
    wire N__6931;
    wire N__6926;
    wire N__6925;
    wire N__6922;
    wire N__6919;
    wire N__6916;
    wire N__6911;
    wire N__6908;
    wire N__6905;
    wire N__6902;
    wire N__6901;
    wire N__6898;
    wire N__6895;
    wire N__6892;
    wire N__6887;
    wire N__6884;
    wire N__6881;
    wire N__6880;
    wire N__6877;
    wire N__6874;
    wire N__6871;
    wire N__6870;
    wire N__6869;
    wire N__6866;
    wire N__6863;
    wire N__6860;
    wire N__6857;
    wire N__6848;
    wire N__6847;
    wire N__6846;
    wire N__6845;
    wire N__6844;
    wire N__6843;
    wire N__6842;
    wire N__6835;
    wire N__6828;
    wire N__6825;
    wire N__6820;
    wire N__6815;
    wire N__6812;
    wire N__6811;
    wire N__6808;
    wire N__6805;
    wire N__6802;
    wire N__6797;
    wire N__6796;
    wire N__6793;
    wire N__6790;
    wire N__6787;
    wire N__6784;
    wire N__6779;
    wire N__6776;
    wire N__6773;
    wire N__6770;
    wire N__6767;
    wire N__6764;
    wire N__6761;
    wire N__6758;
    wire N__6755;
    wire N__6754;
    wire N__6751;
    wire N__6748;
    wire N__6747;
    wire N__6744;
    wire N__6741;
    wire N__6738;
    wire N__6735;
    wire N__6734;
    wire N__6733;
    wire N__6732;
    wire N__6731;
    wire N__6730;
    wire N__6729;
    wire N__6726;
    wire N__6723;
    wire N__6704;
    wire N__6701;
    wire N__6698;
    wire N__6695;
    wire N__6692;
    wire N__6689;
    wire N__6686;
    wire N__6683;
    wire N__6680;
    wire N__6677;
    wire N__6674;
    wire N__6671;
    wire N__6668;
    wire N__6665;
    wire N__6662;
    wire N__6659;
    wire N__6656;
    wire N__6653;
    wire N__6650;
    wire N__6649;
    wire N__6646;
    wire N__6643;
    wire N__6638;
    wire N__6635;
    wire N__6634;
    wire N__6631;
    wire N__6628;
    wire N__6623;
    wire N__6620;
    wire N__6619;
    wire N__6616;
    wire N__6613;
    wire N__6608;
    wire N__6605;
    wire N__6602;
    wire N__6599;
    wire N__6596;
    wire N__6593;
    wire N__6590;
    wire N__6587;
    wire N__6584;
    wire N__6581;
    wire N__6578;
    wire N__6575;
    wire N__6572;
    wire N__6571;
    wire N__6566;
    wire N__6563;
    wire N__6562;
    wire N__6559;
    wire N__6556;
    wire N__6555;
    wire N__6554;
    wire N__6551;
    wire N__6548;
    wire N__6545;
    wire N__6542;
    wire N__6539;
    wire N__6536;
    wire N__6533;
    wire N__6530;
    wire N__6525;
    wire N__6522;
    wire N__6519;
    wire N__6516;
    wire N__6513;
    wire N__6510;
    wire N__6505;
    wire N__6500;
    wire N__6497;
    wire N__6494;
    wire N__6491;
    wire N__6488;
    wire N__6485;
    wire N__6482;
    wire N__6479;
    wire N__6476;
    wire N__6473;
    wire N__6470;
    wire N__6467;
    wire N__6464;
    wire N__6461;
    wire N__6458;
    wire N__6455;
    wire N__6452;
    wire N__6449;
    wire N__6446;
    wire N__6443;
    wire N__6440;
    wire N__6437;
    wire N__6434;
    wire N__6431;
    wire N__6428;
    wire N__6425;
    wire N__6422;
    wire N__6419;
    wire N__6416;
    wire N__6413;
    wire N__6410;
    wire N__6407;
    wire N__6404;
    wire N__6401;
    wire N__6398;
    wire N__6395;
    wire N__6392;
    wire N__6389;
    wire N__6386;
    wire N__6383;
    wire N__6380;
    wire N__6377;
    wire N__6376;
    wire N__6375;
    wire N__6374;
    wire N__6371;
    wire N__6368;
    wire N__6365;
    wire N__6364;
    wire N__6361;
    wire N__6358;
    wire N__6357;
    wire N__6356;
    wire N__6355;
    wire N__6354;
    wire N__6351;
    wire N__6348;
    wire N__6345;
    wire N__6340;
    wire N__6337;
    wire N__6330;
    wire N__6317;
    wire N__6314;
    wire N__6311;
    wire N__6308;
    wire N__6305;
    wire N__6302;
    wire N__6299;
    wire N__6296;
    wire N__6293;
    wire N__6290;
    wire N__6287;
    wire N__6284;
    wire N__6281;
    wire N__6278;
    wire N__6275;
    wire N__6272;
    wire N__6269;
    wire N__6266;
    wire N__6263;
    wire N__6260;
    wire N__6257;
    wire N__6254;
    wire N__6251;
    wire N__6248;
    wire N__6245;
    wire N__6242;
    wire N__6239;
    wire N__6236;
    wire N__6233;
    wire N__6230;
    wire N__6229;
    wire N__6228;
    wire N__6225;
    wire N__6224;
    wire N__6223;
    wire N__6220;
    wire N__6217;
    wire N__6214;
    wire N__6205;
    wire N__6202;
    wire N__6199;
    wire N__6198;
    wire N__6195;
    wire N__6192;
    wire N__6189;
    wire N__6182;
    wire N__6179;
    wire N__6176;
    wire N__6173;
    wire N__6170;
    wire N__6167;
    wire N__6164;
    wire N__6161;
    wire N__6158;
    wire N__6155;
    wire N__6152;
    wire N__6151;
    wire N__6148;
    wire N__6147;
    wire N__6146;
    wire N__6141;
    wire N__6136;
    wire N__6133;
    wire N__6130;
    wire N__6127;
    wire N__6122;
    wire N__6119;
    wire N__6116;
    wire N__6113;
    wire N__6110;
    wire N__6107;
    wire N__6104;
    wire N__6101;
    wire N__6098;
    wire N__6095;
    wire N__6092;
    wire N__6089;
    wire N__6088;
    wire N__6087;
    wire N__6084;
    wire N__6083;
    wire N__6082;
    wire N__6081;
    wire N__6078;
    wire N__6075;
    wire N__6074;
    wire N__6073;
    wire N__6070;
    wire N__6069;
    wire N__6068;
    wire N__6067;
    wire N__6066;
    wire N__6059;
    wire N__6056;
    wire N__6053;
    wire N__6050;
    wire N__6047;
    wire N__6044;
    wire N__6039;
    wire N__6034;
    wire N__6017;
    wire N__6014;
    wire N__6011;
    wire N__6008;
    wire N__6005;
    wire N__6004;
    wire N__6003;
    wire N__6000;
    wire N__5997;
    wire N__5994;
    wire N__5993;
    wire N__5992;
    wire N__5991;
    wire N__5988;
    wire N__5983;
    wire N__5980;
    wire N__5977;
    wire N__5974;
    wire N__5971;
    wire N__5966;
    wire N__5957;
    wire N__5954;
    wire N__5953;
    wire N__5950;
    wire N__5949;
    wire N__5948;
    wire N__5945;
    wire N__5942;
    wire N__5939;
    wire N__5936;
    wire N__5929;
    wire N__5924;
    wire N__5921;
    wire N__5920;
    wire N__5919;
    wire N__5916;
    wire N__5915;
    wire N__5914;
    wire N__5911;
    wire N__5908;
    wire N__5905;
    wire N__5902;
    wire N__5899;
    wire N__5892;
    wire N__5885;
    wire N__5884;
    wire N__5883;
    wire N__5880;
    wire N__5877;
    wire N__5874;
    wire N__5873;
    wire N__5872;
    wire N__5871;
    wire N__5870;
    wire N__5869;
    wire N__5866;
    wire N__5863;
    wire N__5860;
    wire N__5857;
    wire N__5854;
    wire N__5851;
    wire N__5846;
    wire N__5843;
    wire N__5836;
    wire N__5825;
    wire N__5822;
    wire N__5819;
    wire N__5816;
    wire N__5815;
    wire N__5812;
    wire N__5809;
    wire N__5804;
    wire N__5801;
    wire N__5798;
    wire N__5795;
    wire N__5794;
    wire N__5793;
    wire N__5792;
    wire N__5791;
    wire N__5790;
    wire N__5787;
    wire N__5782;
    wire N__5777;
    wire N__5774;
    wire N__5771;
    wire N__5766;
    wire N__5759;
    wire N__5756;
    wire N__5755;
    wire N__5752;
    wire N__5749;
    wire N__5748;
    wire N__5747;
    wire N__5744;
    wire N__5741;
    wire N__5738;
    wire N__5735;
    wire N__5732;
    wire N__5723;
    wire N__5722;
    wire N__5719;
    wire N__5716;
    wire N__5713;
    wire N__5712;
    wire N__5707;
    wire N__5704;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5681;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5671;
    wire N__5670;
    wire N__5669;
    wire N__5666;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5654;
    wire N__5651;
    wire N__5648;
    wire N__5647;
    wire N__5644;
    wire N__5641;
    wire N__5636;
    wire N__5633;
    wire N__5624;
    wire N__5621;
    wire N__5620;
    wire N__5619;
    wire N__5618;
    wire N__5617;
    wire N__5614;
    wire N__5611;
    wire N__5608;
    wire N__5605;
    wire N__5602;
    wire N__5599;
    wire N__5596;
    wire N__5585;
    wire N__5584;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5572;
    wire N__5569;
    wire N__5568;
    wire N__5567;
    wire N__5564;
    wire N__5563;
    wire N__5560;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5544;
    wire N__5537;
    wire N__5534;
    wire N__5531;
    wire N__5528;
    wire N__5525;
    wire N__5522;
    wire N__5521;
    wire N__5520;
    wire N__5517;
    wire N__5512;
    wire N__5507;
    wire N__5504;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5489;
    wire N__5486;
    wire N__5483;
    wire N__5480;
    wire N__5477;
    wire N__5474;
    wire N__5471;
    wire N__5468;
    wire N__5465;
    wire N__5462;
    wire N__5459;
    wire N__5456;
    wire N__5455;
    wire N__5454;
    wire N__5449;
    wire N__5448;
    wire N__5447;
    wire N__5446;
    wire N__5445;
    wire N__5444;
    wire N__5443;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5433;
    wire N__5430;
    wire N__5427;
    wire N__5424;
    wire N__5417;
    wire N__5414;
    wire N__5411;
    wire N__5396;
    wire N__5393;
    wire N__5390;
    wire N__5387;
    wire N__5384;
    wire N__5381;
    wire N__5378;
    wire N__5375;
    wire N__5372;
    wire N__5369;
    wire N__5366;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5354;
    wire N__5353;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5339;
    wire N__5338;
    wire N__5333;
    wire N__5330;
    wire N__5327;
    wire N__5326;
    wire N__5325;
    wire N__5322;
    wire N__5319;
    wire N__5316;
    wire N__5309;
    wire N__5306;
    wire N__5305;
    wire N__5302;
    wire N__5299;
    wire N__5294;
    wire N__5291;
    wire N__5290;
    wire N__5289;
    wire N__5286;
    wire N__5283;
    wire N__5280;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5246;
    wire N__5243;
    wire N__5240;
    wire N__5237;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5222;
    wire N__5219;
    wire N__5216;
    wire N__5213;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5198;
    wire N__5195;
    wire N__5192;
    wire N__5189;
    wire N__5186;
    wire N__5183;
    wire N__5180;
    wire N__5177;
    wire N__5174;
    wire N__5171;
    wire N__5168;
    wire N__5165;
    wire N__5162;
    wire N__5159;
    wire N__5156;
    wire N__5153;
    wire N__5150;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5135;
    wire N__5132;
    wire N__5129;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5117;
    wire N__5114;
    wire N__5111;
    wire N__5108;
    wire N__5105;
    wire N__5102;
    wire N__5099;
    wire N__5096;
    wire N__5095;
    wire N__5094;
    wire N__5093;
    wire N__5092;
    wire N__5091;
    wire N__5090;
    wire N__5087;
    wire N__5084;
    wire N__5081;
    wire N__5076;
    wire N__5071;
    wire N__5060;
    wire N__5057;
    wire N__5054;
    wire N__5051;
    wire N__5048;
    wire N__5045;
    wire N__5042;
    wire N__5041;
    wire N__5038;
    wire N__5035;
    wire N__5032;
    wire N__5029;
    wire N__5024;
    wire N__5021;
    wire N__5020;
    wire N__5017;
    wire N__5012;
    wire N__5009;
    wire N__5006;
    wire N__5003;
    wire N__5002;
    wire N__4999;
    wire N__4998;
    wire N__4995;
    wire N__4992;
    wire N__4989;
    wire N__4982;
    wire N__4979;
    wire N__4978;
    wire N__4977;
    wire N__4974;
    wire N__4971;
    wire N__4968;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4943;
    wire N__4942;
    wire N__4939;
    wire N__4936;
    wire N__4931;
    wire N__4930;
    wire N__4927;
    wire N__4924;
    wire N__4919;
    wire N__4918;
    wire N__4917;
    wire N__4916;
    wire N__4907;
    wire N__4904;
    wire N__4903;
    wire N__4902;
    wire N__4897;
    wire N__4894;
    wire N__4889;
    wire N__4886;
    wire N__4883;
    wire N__4880;
    wire N__4877;
    wire N__4876;
    wire N__4873;
    wire N__4870;
    wire N__4865;
    wire N__4862;
    wire N__4859;
    wire N__4856;
    wire N__4853;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4841;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4813;
    wire N__4810;
    wire N__4807;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4793;
    wire N__4792;
    wire N__4789;
    wire N__4786;
    wire N__4781;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4747;
    wire N__4744;
    wire N__4741;
    wire N__4738;
    wire N__4735;
    wire N__4732;
    wire N__4729;
    wire N__4726;
    wire N__4723;
    wire N__4718;
    wire N__4715;
    wire N__4712;
    wire N__4709;
    wire N__4706;
    wire N__4703;
    wire N__4700;
    wire N__4699;
    wire N__4696;
    wire N__4693;
    wire N__4688;
    wire N__4687;
    wire N__4684;
    wire N__4681;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4667;
    wire N__4664;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4652;
    wire N__4649;
    wire N__4648;
    wire N__4645;
    wire N__4642;
    wire N__4637;
    wire N__4636;
    wire N__4633;
    wire N__4630;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4591;
    wire N__4588;
    wire N__4585;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4562;
    wire N__4559;
    wire N__4556;
    wire N__4553;
    wire N__4552;
    wire N__4549;
    wire N__4546;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4525;
    wire N__4522;
    wire N__4519;
    wire N__4516;
    wire N__4513;
    wire N__4510;
    wire N__4507;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4484;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4471;
    wire N__4468;
    wire N__4465;
    wire N__4460;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4450;
    wire N__4447;
    wire N__4446;
    wire N__4443;
    wire N__4442;
    wire N__4441;
    wire N__4440;
    wire N__4437;
    wire N__4434;
    wire N__4431;
    wire N__4424;
    wire N__4415;
    wire N__4414;
    wire N__4413;
    wire N__4412;
    wire N__4409;
    wire N__4408;
    wire N__4407;
    wire N__4400;
    wire N__4397;
    wire N__4394;
    wire N__4391;
    wire N__4388;
    wire N__4385;
    wire N__4376;
    wire N__4373;
    wire N__4370;
    wire N__4369;
    wire N__4366;
    wire N__4363;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4343;
    wire N__4340;
    wire N__4337;
    wire N__4336;
    wire N__4333;
    wire N__4330;
    wire N__4329;
    wire N__4326;
    wire N__4323;
    wire N__4320;
    wire N__4317;
    wire N__4312;
    wire N__4309;
    wire N__4306;
    wire N__4301;
    wire N__4298;
    wire N__4295;
    wire N__4292;
    wire N__4289;
    wire N__4288;
    wire N__4285;
    wire N__4282;
    wire N__4279;
    wire N__4278;
    wire N__4275;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4263;
    wire N__4260;
    wire N__4257;
    wire N__4250;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4240;
    wire N__4235;
    wire N__4232;
    wire N__4229;
    wire N__4226;
    wire N__4223;
    wire N__4220;
    wire N__4217;
    wire N__4214;
    wire N__4213;
    wire N__4210;
    wire N__4207;
    wire N__4202;
    wire N__4199;
    wire N__4196;
    wire N__4193;
    wire N__4190;
    wire N__4187;
    wire N__4186;
    wire N__4185;
    wire N__4184;
    wire N__4181;
    wire N__4180;
    wire N__4177;
    wire N__4174;
    wire N__4171;
    wire N__4166;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4148;
    wire N__4145;
    wire N__4142;
    wire N__4139;
    wire N__4136;
    wire N__4133;
    wire N__4130;
    wire N__4127;
    wire N__4124;
    wire N__4123;
    wire N__4120;
    wire N__4117;
    wire N__4114;
    wire N__4111;
    wire N__4108;
    wire N__4105;
    wire N__4102;
    wire N__4099;
    wire N__4096;
    wire N__4093;
    wire N__4088;
    wire N__4087;
    wire N__4082;
    wire N__4079;
    wire N__4078;
    wire N__4075;
    wire N__4072;
    wire N__4067;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4052;
    wire N__4049;
    wire N__4046;
    wire N__4043;
    wire N__4040;
    wire N__4037;
    wire N__4034;
    wire N__4031;
    wire N__4028;
    wire N__4025;
    wire N__4022;
    wire N__4019;
    wire N__4018;
    wire N__4017;
    wire N__4014;
    wire N__4009;
    wire N__4004;
    wire N__4001;
    wire N__3998;
    wire N__3995;
    wire N__3992;
    wire N__3989;
    wire N__3986;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire N_1062_i;
    wire CLK80_PLL_i_i;
    wire REGSPACEn_c;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.N_348 ;
    wire DBRn_c_i_cascade_;
    wire DBRn_c_i_0;
    wire C1_c;
    wire \U712_REG_SM.REG_CYCLE_START_RNITO6SZ0Z1 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_0 ;
    wire \U712_REG_SM.N_319 ;
    wire ASn_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_cascade_ ;
    wire DBRn_c_i;
    wire \INVU712_CHIP_RAM.DMA_A20C_net ;
    wire \U712_REG_SM.C1_SYNC_RNIAS4F1Z0Z_1 ;
    wire \U712_REG_SM.N_346_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_2 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_1 ;
    wire \U712_REG_SM.STATE_COUNT_srsts_i_i_0_o2_0_1_3_cascade_ ;
    wire \U712_REG_SM.N_342 ;
    wire \U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0_0 ;
    wire \U712_REG_SM.N_106 ;
    wire \U712_REG_SM.N_379 ;
    wire DBRn_c;
    wire REGENn_c;
    wire VBENn_c;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0 ;
    wire \U712_CHIP_RAM.N_409 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0_1 ;
    wire \U712_CHIP_RAM.N_489_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_0_cascade_ ;
    wire \U712_CHIP_RAM.N_361_cascade_ ;
    wire A_c_20;
    wire \U712_CHIP_RAM.DMA_AZ0Z20 ;
    wire \U712_CHIP_RAM.N_416_cascade_ ;
    wire \U712_CHIP_RAM.BANK0_RNOZ0Z_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_i_i_0 ;
    wire BANK0_c;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3_cascade_ ;
    wire \U712_CHIP_RAM.N_410_cascade_ ;
    wire C3_c;
    wire \U712_REG_SM.STATE_COUNT_RNI4BRHZ0Z_3 ;
    wire \U712_REG_SM.N_400 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_12_0 ;
    wire LATCH_CLK_c;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_2 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ;
    wire DBR_SYNCZ0Z_0;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire TACK_OUTn;
    wire TACK_EN_i_ess;
    wire A_c_18;
    wire A_c_16;
    wire \U712_CHIP_RAM.N_489 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0 ;
    wire TSn_c;
    wire RAMSPACEn_c;
    wire AWEn_c;
    wire DBDIR_c;
    wire CONSTANT_ONE_NET;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_cascade_ ;
    wire \U712_CHIP_RAM.N_304 ;
    wire \U712_CHIP_RAM.N_62_cascade_ ;
    wire \U712_CHIP_RAM.N_452 ;
    wire \U712_CHIP_RAM.N_452_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_11_cascade_ ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.N_288_cascade_ ;
    wire \U712_CHIP_RAM.N_372_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1_1_cascade_ ;
    wire \U712_CHIP_RAM.N_366_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_15_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_0_0 ;
    wire A_c_5;
    wire A_c_12;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ;
    wire \U712_CHIP_RAM.N_448 ;
    wire \U712_CHIP_RAM.N_345_cascade_ ;
    wire A_c_2;
    wire A_c_9;
    wire \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_i_0_cascade_ ;
    wire \U712_CHIP_RAM.N_11_2 ;
    wire REG_TACK;
    wire CPU_TACKm;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.TACK_EN6_0_cascade_ ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CYCLE_TERM.N_316_i_0_en ;
    wire \U712_CYCLE_TERM.N_316_i_0_en_0 ;
    wire \U712_BYTE_ENABLE.N_282_i ;
    wire A_c_4;
    wire A_c_11;
    wire \U712_CHIP_RAM.N_371_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_a2_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_0_0_0 ;
    wire \U712_CHIP_RAM.N_371_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_ ;
    wire \U712_CHIP_RAM.N_288 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0 ;
    wire \U712_CHIP_RAM.N_329 ;
    wire \U712_CHIP_RAM.N_414_cascade_ ;
    wire \U712_CHIP_RAM.N_86 ;
    wire DBR_SYNCZ0Z_1;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_373 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER15 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_1 ;
    wire \U712_CHIP_RAM.N_286_cascade_ ;
    wire \U712_CHIP_RAM.N_486 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a2_1 ;
    wire \U712_CHIP_RAM.N_287_cascade_ ;
    wire \U712_CHIP_RAM.N_436 ;
    wire \U712_CHIP_RAM.N_283 ;
    wire \U712_CHIP_RAM.N_347 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_i_0_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_129_i_0_0 ;
    wire \U712_CHIP_RAM.N_286 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.C1_SYNC_RNIAS4F1_0Z0Z_1_cascade_ ;
    wire \U712_REG_SM.ASn_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a2_0_1 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_REG_SM.C1_SYNC_RNIAS4F1_0Z0Z_1 ;
    wire \U712_REG_SM.N_104 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNO_6Z0Z_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1 ;
    wire \U712_CHIP_RAM.N_287 ;
    wire \U712_CHIP_RAM.N_388 ;
    wire \U712_CHIP_RAM.N_370 ;
    wire \U712_BYTE_ENABLE.un1_CUUBEn_i_0_aZ0Z2 ;
    wire N_38_i;
    wire \U712_BYTE_ENABLE.N_426_cascade_ ;
    wire N_47_i;
    wire \U712_BYTE_ENABLE.un1_CLMBEn_i_0_aZ0Z2 ;
    wire DBENn_c;
    wire N_46_i;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2Z0Z_0 ;
    wire \U712_BYTE_ENABLE.N_431 ;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2Z0Z_0_cascade_ ;
    wire N_45_i;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2Z0Z_0 ;
    wire RnW_c;
    wire N_344;
    wire DMA_LATCH_EN_c;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_ ;
    wire CMA_c_7;
    wire A_c_8;
    wire A_c_15;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_ ;
    wire CMA_c_6;
    wire bfn_11_6_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.N_62 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.N_434_i ;
    wire bfn_11_7_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire C1_c_g;
    wire DMA_CYCLEm;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_201_i_i_a2_3_1 ;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire WRITE_CYCLEm;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.N_306_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_i_0 ;
    wire \U712_CHIP_RAM.REFRESH5lto1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH5lto2 ;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.un3_DMA_CYCLE_START ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ;
    wire CMA_c_2;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ;
    wire \U712_CHIP_RAM.CMA_5_0_8_cascade_ ;
    wire A_c_14;
    wire A_c_7;
    wire \U712_CHIP_RAM.N_463_cascade_ ;
    wire \U712_CHIP_RAM.un1_CMA28_0_i ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRTZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ;
    wire CLK40_PLL_i;
    wire CLK40_PLL_i_i;
    wire RESETn_c;
    wire RESETn_c_i;
    wire CASLn_c;
    wire CASUn_c;
    wire REG_CYCLEm;
    wire DRDENn_c;
    wire CRCSn_c;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire CMA_c_3;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CMA_c_10;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.CMA_5_sn_N_5_mux ;
    wire \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9 ;
    wire CMA_c_4;
    wire A_c_19;
    wire CMA_c_9;
    wire A_c_17;
    wire \U712_CHIP_RAM.CMA_5_0_8 ;
    wire CMA_c_8;
    wire A_c_3;
    wire A_c_10;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_0 ;
    wire A_c_13;
    wire A_c_6;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \INVU712_CHIP_RAM.DMA_A1_nesrC_net ;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire CASn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire WEn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire RASn_c;
    wire CLK80_PLL;
    wire CPU_CYCLEm;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire DRA_c_6;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire N_357_i;
    wire N_42;
    wire N_231;
    wire DRA_c_2;
    wire DRA_c_1;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire DRA_c_3;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire N_358_i;
    wire DS_ENm;
    wire N_40;
    wire A_c_1;
    wire A_c_0;
    wire SIZ_c_0;
    wire SIZ_c_1;
    wire LLBEn_c;
    wire DRA_c_9;
    wire RAS0n_c;
    wire AGNUS_REV_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire _gnd_net_;
    wire C3_c_g;
    wire DBRn_c_i_0_g;
    wire RESETn_c_i_g;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL_i),
            .REFERENCECLK(N__4004),
            .RESETB(N__5051),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__11973),
            .DIN(N__11972),
            .DOUT(N__11971),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__11973),
            .PADOUT(N__11972),
            .PADIN(N__11971),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6233),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__11964),
            .DIN(N__11963),
            .DOUT(N__11962),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__11964),
            .PADOUT(N__11963),
            .PADIN(N__11962),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__11955),
            .DIN(N__11954),
            .DOUT(N__11953),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__11955),
            .PADOUT(N__11954),
            .PADIN(N__11953),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8921),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__11946),
            .DIN(N__11945),
            .DOUT(N__11944),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__11946),
            .PADOUT(N__11945),
            .PADIN(N__11944),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6500),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__11937),
            .DIN(N__11936),
            .DOUT(N__11935),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__11937),
            .PADOUT(N__11936),
            .PADIN(N__11935),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__11928),
            .DIN(N__11927),
            .DOUT(N__11926),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__11928),
            .PADOUT(N__11927),
            .PADIN(N__11926),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__11919),
            .DIN(N__11918),
            .DOUT(N__11917),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__11919),
            .PADOUT(N__11918),
            .PADIN(N__11917),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__11910),
            .DIN(N__11909),
            .DOUT(N__11908),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__11910),
            .PADOUT(N__11909),
            .PADIN(N__11908),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__11901),
            .DIN(N__11900),
            .DOUT(N__11899),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__11901),
            .PADOUT(N__11900),
            .PADIN(N__11899),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__11892),
            .DIN(N__11891),
            .DOUT(N__11890),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__11892),
            .PADOUT(N__11891),
            .PADIN(N__11890),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__11883),
            .DIN(N__11882),
            .DOUT(N__11881),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__11883),
            .PADOUT(N__11882),
            .PADIN(N__11881),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6446),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__11874),
            .DIN(N__11873),
            .DOUT(N__11872),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__11874),
            .PADOUT(N__11873),
            .PADIN(N__11872),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10664),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__11865),
            .DIN(N__11864),
            .DOUT(N__11863),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__11865),
            .PADOUT(N__11864),
            .PADIN(N__11863),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__11856),
            .DIN(N__11855),
            .DOUT(N__11854),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__11856),
            .PADOUT(N__11855),
            .PADIN(N__11854),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__11847),
            .DIN(N__11846),
            .DOUT(N__11845),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__11847),
            .PADOUT(N__11846),
            .PADIN(N__11845),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__11838),
            .DIN(N__11837),
            .DOUT(N__11836),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__11838),
            .PADOUT(N__11837),
            .PADIN(N__11836),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4250),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__11829),
            .DIN(N__11828),
            .DOUT(N__11827),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__11829),
            .PADOUT(N__11828),
            .PADIN(N__11827),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__11820),
            .DIN(N__11819),
            .DOUT(N__11818),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__11820),
            .PADOUT(N__11819),
            .PADIN(N__11818),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__11811),
            .DIN(N__11810),
            .DOUT(N__11809),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__11811),
            .PADOUT(N__11810),
            .PADIN(N__11809),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8894),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__11802),
            .DIN(N__11801),
            .DOUT(N__11800),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__11802),
            .PADOUT(N__11801),
            .PADIN(N__11800),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__11793),
            .DIN(N__11792),
            .DOUT(N__11791),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__11793),
            .PADOUT(N__11792),
            .PADIN(N__11791),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8057),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__11784),
            .DIN(N__11783),
            .DOUT(N__11782),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__11784),
            .PADOUT(N__11783),
            .PADIN(N__11782),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__11775),
            .DIN(N__11774),
            .DOUT(N__11773),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__11775),
            .PADOUT(N__11774),
            .PADIN(N__11773),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9980),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__11766),
            .DIN(N__11765),
            .DOUT(N__11764),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__11766),
            .PADOUT(N__11765),
            .PADIN(N__11764),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__11757),
            .DIN(N__11756),
            .DOUT(N__11755),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__11757),
            .PADOUT(N__11756),
            .PADIN(N__11755),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__11748),
            .DIN(N__11747),
            .DOUT(N__11746),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__11748),
            .PADOUT(N__11747),
            .PADIN(N__11746),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__11739),
            .DIN(N__11738),
            .DOUT(N__11737),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__11739),
            .PADOUT(N__11738),
            .PADIN(N__11737),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__11730),
            .DIN(N__11729),
            .DOUT(N__11728),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__11730),
            .PADOUT(N__11729),
            .PADIN(N__11728),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__11721),
            .DIN(N__11720),
            .DOUT(N__11719),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__11721),
            .PADOUT(N__11720),
            .PADIN(N__11719),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6476),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__11712),
            .DIN(N__11711),
            .DOUT(N__11710),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__11712),
            .PADOUT(N__11711),
            .PADIN(N__11710),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__11703),
            .DIN(N__11702),
            .DOUT(N__11701),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__11703),
            .PADOUT(N__11702),
            .PADIN(N__11701),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__11694),
            .DIN(N__11693),
            .DOUT(N__11692),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__11694),
            .PADOUT(N__11693),
            .PADIN(N__11692),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__11685),
            .DIN(N__11684),
            .DOUT(N__11683),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__11685),
            .PADOUT(N__11684),
            .PADIN(N__11683),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__11676),
            .DIN(N__11675),
            .DOUT(N__11674),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__11676),
            .PADOUT(N__11675),
            .PADIN(N__11674),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__11667),
            .DIN(N__11666),
            .DOUT(N__11665),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__11667),
            .PADOUT(N__11666),
            .PADIN(N__11665),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9842),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__11658),
            .DIN(N__11657),
            .DOUT(N__11656),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__11658),
            .PADOUT(N__11657),
            .PADIN(N__11656),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__11649),
            .DIN(N__11648),
            .DOUT(N__11647),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__11649),
            .PADOUT(N__11648),
            .PADIN(N__11647),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4568),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__11640),
            .DIN(N__11639),
            .DOUT(N__11638),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__11640),
            .PADOUT(N__11639),
            .PADIN(N__11638),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8440),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__11631),
            .DIN(N__11630),
            .DOUT(N__11629),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__11631),
            .PADOUT(N__11630),
            .PADIN(N__11629),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4055),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__11622),
            .DIN(N__11621),
            .DOUT(N__11620),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__11622),
            .PADOUT(N__11621),
            .PADIN(N__11620),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__11613),
            .DIN(N__11612),
            .DOUT(N__11611),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__11613),
            .PADOUT(N__11612),
            .PADIN(N__11611),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4232),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__11604),
            .DIN(N__11603),
            .DOUT(N__11602),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__11604),
            .PADOUT(N__11603),
            .PADIN(N__11602),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8024),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuft_iopad (
            .OE(N__11595),
            .DIN(N__11594),
            .DOUT(N__11593),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO RAMENn_obuft_preio (
            .PADOEN(N__11595),
            .PADOUT(N__11594),
            .PADIN(N__11593),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__11586),
            .DIN(N__11585),
            .DOUT(N__11584),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__11586),
            .PADOUT(N__11585),
            .PADIN(N__11584),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__11577),
            .DIN(N__11576),
            .DOUT(N__11575),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__11577),
            .PADOUT(N__11576),
            .PADIN(N__11575),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__11568),
            .DIN(N__11567),
            .DOUT(N__11566),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__11568),
            .PADOUT(N__11567),
            .PADIN(N__11566),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__11559),
            .DIN(N__11558),
            .DOUT(N__11557),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__11559),
            .PADOUT(N__11558),
            .PADIN(N__11557),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__11550),
            .DIN(N__11549),
            .DOUT(N__11548),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__11550),
            .PADOUT(N__11549),
            .PADIN(N__11548),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8834),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__11541),
            .DIN(N__11540),
            .DOUT(N__11539),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__11541),
            .PADOUT(N__11540),
            .PADIN(N__11539),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__11532),
            .DIN(N__11531),
            .DOUT(N__11530),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__11532),
            .PADOUT(N__11531),
            .PADIN(N__11530),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8415),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__11523),
            .DIN(N__11522),
            .DOUT(N__11521),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__11523),
            .PADOUT(N__11522),
            .PADIN(N__11521),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8690),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__11514),
            .DIN(N__11513),
            .DOUT(N__11512),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__11514),
            .PADOUT(N__11513),
            .PADIN(N__11512),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8078),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__11505),
            .DIN(N__11504),
            .DOUT(N__11503),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__11505),
            .PADOUT(N__11504),
            .PADIN(N__11503),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6587),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__11496),
            .DIN(N__11495),
            .DOUT(N__11494),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__11496),
            .PADOUT(N__11495),
            .PADIN(N__11494),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8648),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__11487),
            .DIN(N__11486),
            .DOUT(N__11485),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__11487),
            .PADOUT(N__11486),
            .PADIN(N__11485),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4295),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__11478),
            .DIN(N__11477),
            .DOUT(N__11476),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__11478),
            .PADOUT(N__11477),
            .PADIN(N__11476),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__11469),
            .DIN(N__11468),
            .DOUT(N__11467),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__11469),
            .PADOUT(N__11468),
            .PADIN(N__11467),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__11460),
            .DIN(N__11459),
            .DOUT(N__11458),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__11460),
            .PADOUT(N__11459),
            .PADIN(N__11458),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6182),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__11451),
            .DIN(N__11450),
            .DOUT(N__11449),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__11451),
            .PADOUT(N__11450),
            .PADIN(N__11449),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9917),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__11442),
            .DIN(N__11441),
            .DOUT(N__11440),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__11442),
            .PADOUT(N__11441),
            .PADIN(N__11440),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4712),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__11433),
            .DIN(N__11432),
            .DOUT(N__11431),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__11433),
            .PADOUT(N__11432),
            .PADIN(N__11431),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6266),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__11424),
            .DIN(N__11423),
            .DOUT(N__11422),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__11424),
            .PADOUT(N__11423),
            .PADIN(N__11422),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__11415),
            .DIN(N__11414),
            .DOUT(N__11413),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__11415),
            .PADOUT(N__11414),
            .PADIN(N__11413),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__11406),
            .DIN(N__11405),
            .DOUT(N__11404),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__11406),
            .PADOUT(N__11405),
            .PADIN(N__11404),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__11397),
            .DIN(N__11396),
            .DOUT(N__11395),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__11397),
            .PADOUT(N__11396),
            .PADIN(N__11395),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__11388),
            .DIN(N__11387),
            .DOUT(N__11386),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__11388),
            .PADOUT(N__11387),
            .PADIN(N__11386),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9155),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__11379),
            .DIN(N__11378),
            .DOUT(N__11377),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__11379),
            .PADOUT(N__11378),
            .PADIN(N__11377),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10391),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__11370),
            .DIN(N__11369),
            .DOUT(N__11368),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__11370),
            .PADOUT(N__11369),
            .PADIN(N__11368),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__11361),
            .DIN(N__11360),
            .DOUT(N__11359),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__11361),
            .PADOUT(N__11360),
            .PADIN(N__11359),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6293),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__11352),
            .DIN(N__11351),
            .DOUT(N__11350),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__11352),
            .PADOUT(N__11351),
            .PADIN(N__11350),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4067),
            .DIN0(),
            .DOUT0(N__4889),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__11343),
            .DIN(N__11342),
            .DOUT(N__11341),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__11343),
            .PADOUT(N__11342),
            .PADIN(N__11341),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7676),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__11334),
            .DIN(N__11333),
            .DOUT(N__11332),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__11334),
            .PADOUT(N__11333),
            .PADIN(N__11332),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__11325),
            .DIN(N__11324),
            .DOUT(N__11323),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__11325),
            .PADOUT(N__11324),
            .PADIN(N__11323),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__11316),
            .DIN(N__11315),
            .DOUT(N__11314),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__11316),
            .PADOUT(N__11315),
            .PADIN(N__11314),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8582),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__11307),
            .DIN(N__11306),
            .DOUT(N__11305),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__11307),
            .PADOUT(N__11306),
            .PADIN(N__11305),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__11298),
            .DIN(N__11297),
            .DOUT(N__11296),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__11298),
            .PADOUT(N__11297),
            .PADIN(N__11296),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__11289),
            .DIN(N__11288),
            .DOUT(N__11287),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__11289),
            .PADOUT(N__11288),
            .PADIN(N__11287),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__11280),
            .DIN(N__11279),
            .DOUT(N__11278),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__11280),
            .PADOUT(N__11279),
            .PADIN(N__11278),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__11271),
            .DIN(N__11270),
            .DOUT(N__11269),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__11271),
            .PADOUT(N__11270),
            .PADIN(N__11269),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8804),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__11262),
            .DIN(N__11261),
            .DOUT(N__11260),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__11262),
            .PADOUT(N__11261),
            .PADIN(N__11260),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10649),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__11253),
            .DIN(N__11252),
            .DOUT(N__11251),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__11253),
            .PADOUT(N__11252),
            .PADIN(N__11251),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10631),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__11244),
            .DIN(N__11243),
            .DOUT(N__11242),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__11244),
            .PADOUT(N__11243),
            .PADIN(N__11242),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4958),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__11235),
            .DIN(N__11234),
            .DOUT(N__11233),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__11235),
            .PADOUT(N__11234),
            .PADIN(N__11233),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__11226),
            .DIN(N__11225),
            .DOUT(N__11224),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__11226),
            .PADOUT(N__11225),
            .PADIN(N__11224),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__11217),
            .DIN(N__11216),
            .DOUT(N__11215),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__11217),
            .PADOUT(N__11216),
            .PADIN(N__11215),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6692),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__11208),
            .DIN(N__11207),
            .DOUT(N__11206),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__11208),
            .PADOUT(N__11207),
            .PADIN(N__11206),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__11199),
            .DIN(N__11198),
            .DOUT(N__11197),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__11199),
            .PADOUT(N__11198),
            .PADIN(N__11197),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__11190),
            .DIN(N__11189),
            .DOUT(N__11188),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__11190),
            .PADOUT(N__11189),
            .PADIN(N__11188),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4664),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__11181),
            .DIN(N__11180),
            .DOUT(N__11179),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__11181),
            .PADOUT(N__11180),
            .PADIN(N__11179),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10346),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__11172),
            .DIN(N__11171),
            .DOUT(N__11170),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__11172),
            .PADOUT(N__11171),
            .PADIN(N__11170),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8441),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2732 (
            .O(N__11153),
            .I(N__11149));
    InMux I__2731 (
            .O(N__11152),
            .I(N__11146));
    LocalMux I__2730 (
            .O(N__11149),
            .I(N__11142));
    LocalMux I__2729 (
            .O(N__11146),
            .I(N__11139));
    InMux I__2728 (
            .O(N__11145),
            .I(N__11136));
    Span4Mux_v I__2727 (
            .O(N__11142),
            .I(N__11133));
    Span4Mux_h I__2726 (
            .O(N__11139),
            .I(N__11128));
    LocalMux I__2725 (
            .O(N__11136),
            .I(N__11128));
    Span4Mux_v I__2724 (
            .O(N__11133),
            .I(N__11124));
    Span4Mux_v I__2723 (
            .O(N__11128),
            .I(N__11121));
    InMux I__2722 (
            .O(N__11127),
            .I(N__11118));
    Sp12to4 I__2721 (
            .O(N__11124),
            .I(N__11115));
    Sp12to4 I__2720 (
            .O(N__11121),
            .I(N__11112));
    LocalMux I__2719 (
            .O(N__11118),
            .I(N__11109));
    Span12Mux_h I__2718 (
            .O(N__11115),
            .I(N__11106));
    Span12Mux_h I__2717 (
            .O(N__11112),
            .I(N__11103));
    Span12Mux_v I__2716 (
            .O(N__11109),
            .I(N__11100));
    Span12Mux_v I__2715 (
            .O(N__11106),
            .I(N__11097));
    Span12Mux_v I__2714 (
            .O(N__11103),
            .I(N__11094));
    Span12Mux_v I__2713 (
            .O(N__11100),
            .I(N__11091));
    Odrv12 I__2712 (
            .O(N__11097),
            .I(DRA_c_9));
    Odrv12 I__2711 (
            .O(N__11094),
            .I(DRA_c_9));
    Odrv12 I__2710 (
            .O(N__11091),
            .I(DRA_c_9));
    InMux I__2709 (
            .O(N__11084),
            .I(N__11081));
    LocalMux I__2708 (
            .O(N__11081),
            .I(N__11078));
    Odrv12 I__2707 (
            .O(N__11078),
            .I(RAS0n_c));
    CascadeMux I__2706 (
            .O(N__11075),
            .I(N__11072));
    InMux I__2705 (
            .O(N__11072),
            .I(N__11066));
    InMux I__2704 (
            .O(N__11071),
            .I(N__11063));
    CascadeMux I__2703 (
            .O(N__11070),
            .I(N__11056));
    CascadeMux I__2702 (
            .O(N__11069),
            .I(N__11050));
    LocalMux I__2701 (
            .O(N__11066),
            .I(N__11043));
    LocalMux I__2700 (
            .O(N__11063),
            .I(N__11043));
    InMux I__2699 (
            .O(N__11062),
            .I(N__11038));
    InMux I__2698 (
            .O(N__11061),
            .I(N__11038));
    InMux I__2697 (
            .O(N__11060),
            .I(N__11033));
    InMux I__2696 (
            .O(N__11059),
            .I(N__11033));
    InMux I__2695 (
            .O(N__11056),
            .I(N__11025));
    InMux I__2694 (
            .O(N__11055),
            .I(N__11025));
    InMux I__2693 (
            .O(N__11054),
            .I(N__11025));
    InMux I__2692 (
            .O(N__11053),
            .I(N__11022));
    InMux I__2691 (
            .O(N__11050),
            .I(N__11017));
    InMux I__2690 (
            .O(N__11049),
            .I(N__11017));
    InMux I__2689 (
            .O(N__11048),
            .I(N__11013));
    Span4Mux_h I__2688 (
            .O(N__11043),
            .I(N__11007));
    LocalMux I__2687 (
            .O(N__11038),
            .I(N__11007));
    LocalMux I__2686 (
            .O(N__11033),
            .I(N__11004));
    CascadeMux I__2685 (
            .O(N__11032),
            .I(N__10997));
    LocalMux I__2684 (
            .O(N__11025),
            .I(N__10993));
    LocalMux I__2683 (
            .O(N__11022),
            .I(N__10988));
    LocalMux I__2682 (
            .O(N__11017),
            .I(N__10988));
    InMux I__2681 (
            .O(N__11016),
            .I(N__10985));
    LocalMux I__2680 (
            .O(N__11013),
            .I(N__10982));
    InMux I__2679 (
            .O(N__11012),
            .I(N__10979));
    Span4Mux_h I__2678 (
            .O(N__11007),
            .I(N__10974));
    Span4Mux_v I__2677 (
            .O(N__11004),
            .I(N__10974));
    InMux I__2676 (
            .O(N__11003),
            .I(N__10969));
    InMux I__2675 (
            .O(N__11002),
            .I(N__10969));
    InMux I__2674 (
            .O(N__11001),
            .I(N__10964));
    InMux I__2673 (
            .O(N__11000),
            .I(N__10964));
    InMux I__2672 (
            .O(N__10997),
            .I(N__10959));
    InMux I__2671 (
            .O(N__10996),
            .I(N__10959));
    Span4Mux_v I__2670 (
            .O(N__10993),
            .I(N__10952));
    Span4Mux_h I__2669 (
            .O(N__10988),
            .I(N__10952));
    LocalMux I__2668 (
            .O(N__10985),
            .I(N__10952));
    Span4Mux_v I__2667 (
            .O(N__10982),
            .I(N__10949));
    LocalMux I__2666 (
            .O(N__10979),
            .I(N__10946));
    Sp12to4 I__2665 (
            .O(N__10974),
            .I(N__10937));
    LocalMux I__2664 (
            .O(N__10969),
            .I(N__10937));
    LocalMux I__2663 (
            .O(N__10964),
            .I(N__10937));
    LocalMux I__2662 (
            .O(N__10959),
            .I(N__10937));
    Sp12to4 I__2661 (
            .O(N__10952),
            .I(N__10934));
    Span4Mux_h I__2660 (
            .O(N__10949),
            .I(N__10931));
    Span12Mux_v I__2659 (
            .O(N__10946),
            .I(N__10928));
    Span12Mux_h I__2658 (
            .O(N__10937),
            .I(N__10925));
    Span12Mux_v I__2657 (
            .O(N__10934),
            .I(N__10922));
    Sp12to4 I__2656 (
            .O(N__10931),
            .I(N__10919));
    Span12Mux_h I__2655 (
            .O(N__10928),
            .I(N__10914));
    Span12Mux_v I__2654 (
            .O(N__10925),
            .I(N__10914));
    Span12Mux_h I__2653 (
            .O(N__10922),
            .I(N__10911));
    Span12Mux_v I__2652 (
            .O(N__10919),
            .I(N__10908));
    Odrv12 I__2651 (
            .O(N__10914),
            .I(AGNUS_REV_c));
    Odrv12 I__2650 (
            .O(N__10911),
            .I(AGNUS_REV_c));
    Odrv12 I__2649 (
            .O(N__10908),
            .I(AGNUS_REV_c));
    InMux I__2648 (
            .O(N__10901),
            .I(N__10898));
    LocalMux I__2647 (
            .O(N__10898),
            .I(N__10895));
    Span12Mux_h I__2646 (
            .O(N__10895),
            .I(N__10892));
    Odrv12 I__2645 (
            .O(N__10892),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    ClkMux I__2644 (
            .O(N__10889),
            .I(N__10868));
    ClkMux I__2643 (
            .O(N__10888),
            .I(N__10868));
    ClkMux I__2642 (
            .O(N__10887),
            .I(N__10868));
    ClkMux I__2641 (
            .O(N__10886),
            .I(N__10868));
    ClkMux I__2640 (
            .O(N__10885),
            .I(N__10868));
    ClkMux I__2639 (
            .O(N__10884),
            .I(N__10868));
    ClkMux I__2638 (
            .O(N__10883),
            .I(N__10868));
    GlobalMux I__2637 (
            .O(N__10868),
            .I(N__10865));
    gio2CtrlBuf I__2636 (
            .O(N__10865),
            .I(C3_c_g));
    CEMux I__2635 (
            .O(N__10862),
            .I(N__10832));
    CEMux I__2634 (
            .O(N__10861),
            .I(N__10832));
    CEMux I__2633 (
            .O(N__10860),
            .I(N__10832));
    CEMux I__2632 (
            .O(N__10859),
            .I(N__10832));
    CEMux I__2631 (
            .O(N__10858),
            .I(N__10832));
    CEMux I__2630 (
            .O(N__10857),
            .I(N__10832));
    CEMux I__2629 (
            .O(N__10856),
            .I(N__10832));
    CEMux I__2628 (
            .O(N__10855),
            .I(N__10832));
    CEMux I__2627 (
            .O(N__10854),
            .I(N__10832));
    CEMux I__2626 (
            .O(N__10853),
            .I(N__10832));
    GlobalMux I__2625 (
            .O(N__10832),
            .I(N__10829));
    gio2CtrlBuf I__2624 (
            .O(N__10829),
            .I(DBRn_c_i_0_g));
    InMux I__2623 (
            .O(N__10826),
            .I(N__10817));
    InMux I__2622 (
            .O(N__10825),
            .I(N__10817));
    InMux I__2621 (
            .O(N__10824),
            .I(N__10814));
    InMux I__2620 (
            .O(N__10823),
            .I(N__10811));
    InMux I__2619 (
            .O(N__10822),
            .I(N__10808));
    LocalMux I__2618 (
            .O(N__10817),
            .I(N__10797));
    LocalMux I__2617 (
            .O(N__10814),
            .I(N__10790));
    LocalMux I__2616 (
            .O(N__10811),
            .I(N__10772));
    LocalMux I__2615 (
            .O(N__10808),
            .I(N__10763));
    SRMux I__2614 (
            .O(N__10807),
            .I(N__10670));
    SRMux I__2613 (
            .O(N__10806),
            .I(N__10670));
    SRMux I__2612 (
            .O(N__10805),
            .I(N__10670));
    SRMux I__2611 (
            .O(N__10804),
            .I(N__10670));
    SRMux I__2610 (
            .O(N__10803),
            .I(N__10670));
    SRMux I__2609 (
            .O(N__10802),
            .I(N__10670));
    SRMux I__2608 (
            .O(N__10801),
            .I(N__10670));
    SRMux I__2607 (
            .O(N__10800),
            .I(N__10670));
    Glb2LocalMux I__2606 (
            .O(N__10797),
            .I(N__10670));
    SRMux I__2605 (
            .O(N__10796),
            .I(N__10670));
    SRMux I__2604 (
            .O(N__10795),
            .I(N__10670));
    SRMux I__2603 (
            .O(N__10794),
            .I(N__10670));
    SRMux I__2602 (
            .O(N__10793),
            .I(N__10670));
    Glb2LocalMux I__2601 (
            .O(N__10790),
            .I(N__10670));
    SRMux I__2600 (
            .O(N__10789),
            .I(N__10670));
    SRMux I__2599 (
            .O(N__10788),
            .I(N__10670));
    SRMux I__2598 (
            .O(N__10787),
            .I(N__10670));
    SRMux I__2597 (
            .O(N__10786),
            .I(N__10670));
    SRMux I__2596 (
            .O(N__10785),
            .I(N__10670));
    SRMux I__2595 (
            .O(N__10784),
            .I(N__10670));
    SRMux I__2594 (
            .O(N__10783),
            .I(N__10670));
    SRMux I__2593 (
            .O(N__10782),
            .I(N__10670));
    SRMux I__2592 (
            .O(N__10781),
            .I(N__10670));
    SRMux I__2591 (
            .O(N__10780),
            .I(N__10670));
    SRMux I__2590 (
            .O(N__10779),
            .I(N__10670));
    SRMux I__2589 (
            .O(N__10778),
            .I(N__10670));
    SRMux I__2588 (
            .O(N__10777),
            .I(N__10670));
    SRMux I__2587 (
            .O(N__10776),
            .I(N__10670));
    SRMux I__2586 (
            .O(N__10775),
            .I(N__10670));
    Glb2LocalMux I__2585 (
            .O(N__10772),
            .I(N__10670));
    SRMux I__2584 (
            .O(N__10771),
            .I(N__10670));
    SRMux I__2583 (
            .O(N__10770),
            .I(N__10670));
    SRMux I__2582 (
            .O(N__10769),
            .I(N__10670));
    SRMux I__2581 (
            .O(N__10768),
            .I(N__10670));
    SRMux I__2580 (
            .O(N__10767),
            .I(N__10670));
    SRMux I__2579 (
            .O(N__10766),
            .I(N__10670));
    Glb2LocalMux I__2578 (
            .O(N__10763),
            .I(N__10670));
    SRMux I__2577 (
            .O(N__10762),
            .I(N__10670));
    SRMux I__2576 (
            .O(N__10761),
            .I(N__10670));
    SRMux I__2575 (
            .O(N__10760),
            .I(N__10670));
    SRMux I__2574 (
            .O(N__10759),
            .I(N__10670));
    SRMux I__2573 (
            .O(N__10758),
            .I(N__10670));
    SRMux I__2572 (
            .O(N__10757),
            .I(N__10670));
    GlobalMux I__2571 (
            .O(N__10670),
            .I(N__10667));
    gio2CtrlBuf I__2570 (
            .O(N__10667),
            .I(RESETn_c_i_g));
    IoInMux I__2569 (
            .O(N__10664),
            .I(N__10661));
    LocalMux I__2568 (
            .O(N__10661),
            .I(N__10658));
    Span4Mux_s0_v I__2567 (
            .O(N__10658),
            .I(N__10655));
    Span4Mux_v I__2566 (
            .O(N__10655),
            .I(N__10652));
    Odrv4 I__2565 (
            .O(N__10652),
            .I(N_357_i));
    IoInMux I__2564 (
            .O(N__10649),
            .I(N__10646));
    LocalMux I__2563 (
            .O(N__10646),
            .I(N__10643));
    Span4Mux_s2_v I__2562 (
            .O(N__10643),
            .I(N__10640));
    Span4Mux_v I__2561 (
            .O(N__10640),
            .I(N__10637));
    Sp12to4 I__2560 (
            .O(N__10637),
            .I(N__10634));
    Odrv12 I__2559 (
            .O(N__10634),
            .I(N_42));
    IoInMux I__2558 (
            .O(N__10631),
            .I(N__10628));
    LocalMux I__2557 (
            .O(N__10628),
            .I(N__10625));
    Span4Mux_s2_v I__2556 (
            .O(N__10625),
            .I(N__10622));
    Span4Mux_h I__2555 (
            .O(N__10622),
            .I(N__10619));
    Span4Mux_v I__2554 (
            .O(N__10619),
            .I(N__10616));
    Odrv4 I__2553 (
            .O(N__10616),
            .I(N_231));
    InMux I__2552 (
            .O(N__10613),
            .I(N__10610));
    LocalMux I__2551 (
            .O(N__10610),
            .I(N__10604));
    InMux I__2550 (
            .O(N__10609),
            .I(N__10599));
    InMux I__2549 (
            .O(N__10608),
            .I(N__10599));
    InMux I__2548 (
            .O(N__10607),
            .I(N__10596));
    Span4Mux_v I__2547 (
            .O(N__10604),
            .I(N__10589));
    LocalMux I__2546 (
            .O(N__10599),
            .I(N__10589));
    LocalMux I__2545 (
            .O(N__10596),
            .I(N__10589));
    Span4Mux_h I__2544 (
            .O(N__10589),
            .I(N__10586));
    Sp12to4 I__2543 (
            .O(N__10586),
            .I(N__10583));
    Span12Mux_v I__2542 (
            .O(N__10583),
            .I(N__10580));
    Odrv12 I__2541 (
            .O(N__10580),
            .I(DRA_c_2));
    InMux I__2540 (
            .O(N__10577),
            .I(N__10572));
    InMux I__2539 (
            .O(N__10576),
            .I(N__10569));
    InMux I__2538 (
            .O(N__10575),
            .I(N__10565));
    LocalMux I__2537 (
            .O(N__10572),
            .I(N__10560));
    LocalMux I__2536 (
            .O(N__10569),
            .I(N__10560));
    InMux I__2535 (
            .O(N__10568),
            .I(N__10557));
    LocalMux I__2534 (
            .O(N__10565),
            .I(N__10554));
    Span4Mux_h I__2533 (
            .O(N__10560),
            .I(N__10551));
    LocalMux I__2532 (
            .O(N__10557),
            .I(N__10548));
    Sp12to4 I__2531 (
            .O(N__10554),
            .I(N__10545));
    Sp12to4 I__2530 (
            .O(N__10551),
            .I(N__10542));
    Span12Mux_h I__2529 (
            .O(N__10548),
            .I(N__10539));
    Span12Mux_v I__2528 (
            .O(N__10545),
            .I(N__10536));
    Span12Mux_v I__2527 (
            .O(N__10542),
            .I(N__10533));
    Span12Mux_v I__2526 (
            .O(N__10539),
            .I(N__10530));
    Span12Mux_h I__2525 (
            .O(N__10536),
            .I(N__10527));
    Odrv12 I__2524 (
            .O(N__10533),
            .I(DRA_c_1));
    Odrv12 I__2523 (
            .O(N__10530),
            .I(DRA_c_1));
    Odrv12 I__2522 (
            .O(N__10527),
            .I(DRA_c_1));
    InMux I__2521 (
            .O(N__10520),
            .I(N__10514));
    InMux I__2520 (
            .O(N__10519),
            .I(N__10514));
    LocalMux I__2519 (
            .O(N__10514),
            .I(N__10511));
    Span4Mux_v I__2518 (
            .O(N__10511),
            .I(N__10508));
    Odrv4 I__2517 (
            .O(N__10508),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__2516 (
            .O(N__10505),
            .I(N__10502));
    LocalMux I__2515 (
            .O(N__10502),
            .I(N__10496));
    InMux I__2514 (
            .O(N__10501),
            .I(N__10491));
    InMux I__2513 (
            .O(N__10500),
            .I(N__10491));
    InMux I__2512 (
            .O(N__10499),
            .I(N__10488));
    Span4Mux_v I__2511 (
            .O(N__10496),
            .I(N__10485));
    LocalMux I__2510 (
            .O(N__10491),
            .I(N__10480));
    LocalMux I__2509 (
            .O(N__10488),
            .I(N__10480));
    Span4Mux_h I__2508 (
            .O(N__10485),
            .I(N__10475));
    Span4Mux_h I__2507 (
            .O(N__10480),
            .I(N__10475));
    Sp12to4 I__2506 (
            .O(N__10475),
            .I(N__10472));
    Span12Mux_v I__2505 (
            .O(N__10472),
            .I(N__10469));
    Odrv12 I__2504 (
            .O(N__10469),
            .I(DRA_c_3));
    InMux I__2503 (
            .O(N__10466),
            .I(N__10461));
    InMux I__2502 (
            .O(N__10465),
            .I(N__10458));
    InMux I__2501 (
            .O(N__10464),
            .I(N__10455));
    LocalMux I__2500 (
            .O(N__10461),
            .I(N__10449));
    LocalMux I__2499 (
            .O(N__10458),
            .I(N__10449));
    LocalMux I__2498 (
            .O(N__10455),
            .I(N__10446));
    InMux I__2497 (
            .O(N__10454),
            .I(N__10443));
    Span4Mux_v I__2496 (
            .O(N__10449),
            .I(N__10440));
    Span4Mux_v I__2495 (
            .O(N__10446),
            .I(N__10437));
    LocalMux I__2494 (
            .O(N__10443),
            .I(N__10434));
    Span4Mux_v I__2493 (
            .O(N__10440),
            .I(N__10431));
    Sp12to4 I__2492 (
            .O(N__10437),
            .I(N__10428));
    Sp12to4 I__2491 (
            .O(N__10434),
            .I(N__10425));
    Sp12to4 I__2490 (
            .O(N__10431),
            .I(N__10422));
    Span12Mux_h I__2489 (
            .O(N__10428),
            .I(N__10419));
    Span12Mux_v I__2488 (
            .O(N__10425),
            .I(N__10416));
    Span12Mux_h I__2487 (
            .O(N__10422),
            .I(N__10413));
    Span12Mux_v I__2486 (
            .O(N__10419),
            .I(N__10408));
    Span12Mux_h I__2485 (
            .O(N__10416),
            .I(N__10408));
    Odrv12 I__2484 (
            .O(N__10413),
            .I(DRA_c_4));
    Odrv12 I__2483 (
            .O(N__10408),
            .I(DRA_c_4));
    InMux I__2482 (
            .O(N__10403),
            .I(N__10400));
    LocalMux I__2481 (
            .O(N__10400),
            .I(N__10397));
    Span4Mux_h I__2480 (
            .O(N__10397),
            .I(N__10394));
    Odrv4 I__2479 (
            .O(N__10394),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    IoInMux I__2478 (
            .O(N__10391),
            .I(N__10388));
    LocalMux I__2477 (
            .O(N__10388),
            .I(N__10385));
    Span4Mux_s0_v I__2476 (
            .O(N__10385),
            .I(N__10382));
    Span4Mux_v I__2475 (
            .O(N__10382),
            .I(N__10379));
    Odrv4 I__2474 (
            .O(N__10379),
            .I(N_358_i));
    InMux I__2473 (
            .O(N__10376),
            .I(N__10372));
    InMux I__2472 (
            .O(N__10375),
            .I(N__10369));
    LocalMux I__2471 (
            .O(N__10372),
            .I(N__10366));
    LocalMux I__2470 (
            .O(N__10369),
            .I(N__10361));
    Span4Mux_h I__2469 (
            .O(N__10366),
            .I(N__10361));
    Sp12to4 I__2468 (
            .O(N__10361),
            .I(N__10358));
    Span12Mux_v I__2467 (
            .O(N__10358),
            .I(N__10354));
    InMux I__2466 (
            .O(N__10357),
            .I(N__10351));
    Odrv12 I__2465 (
            .O(N__10354),
            .I(DS_ENm));
    LocalMux I__2464 (
            .O(N__10351),
            .I(DS_ENm));
    IoInMux I__2463 (
            .O(N__10346),
            .I(N__10343));
    LocalMux I__2462 (
            .O(N__10343),
            .I(N__10340));
    Span4Mux_s2_v I__2461 (
            .O(N__10340),
            .I(N__10337));
    Span4Mux_v I__2460 (
            .O(N__10337),
            .I(N__10334));
    Sp12to4 I__2459 (
            .O(N__10334),
            .I(N__10331));
    Odrv12 I__2458 (
            .O(N__10331),
            .I(N_40));
    InMux I__2457 (
            .O(N__10328),
            .I(N__10323));
    InMux I__2456 (
            .O(N__10327),
            .I(N__10317));
    InMux I__2455 (
            .O(N__10326),
            .I(N__10317));
    LocalMux I__2454 (
            .O(N__10323),
            .I(N__10314));
    InMux I__2453 (
            .O(N__10322),
            .I(N__10311));
    LocalMux I__2452 (
            .O(N__10317),
            .I(N__10308));
    Span4Mux_h I__2451 (
            .O(N__10314),
            .I(N__10301));
    LocalMux I__2450 (
            .O(N__10311),
            .I(N__10301));
    Span4Mux_v I__2449 (
            .O(N__10308),
            .I(N__10298));
    InMux I__2448 (
            .O(N__10307),
            .I(N__10295));
    InMux I__2447 (
            .O(N__10306),
            .I(N__10292));
    Span4Mux_v I__2446 (
            .O(N__10301),
            .I(N__10288));
    Span4Mux_v I__2445 (
            .O(N__10298),
            .I(N__10285));
    LocalMux I__2444 (
            .O(N__10295),
            .I(N__10280));
    LocalMux I__2443 (
            .O(N__10292),
            .I(N__10280));
    InMux I__2442 (
            .O(N__10291),
            .I(N__10277));
    Span4Mux_v I__2441 (
            .O(N__10288),
            .I(N__10273));
    Span4Mux_v I__2440 (
            .O(N__10285),
            .I(N__10268));
    Span4Mux_v I__2439 (
            .O(N__10280),
            .I(N__10268));
    LocalMux I__2438 (
            .O(N__10277),
            .I(N__10265));
    InMux I__2437 (
            .O(N__10276),
            .I(N__10262));
    Sp12to4 I__2436 (
            .O(N__10273),
            .I(N__10253));
    Sp12to4 I__2435 (
            .O(N__10268),
            .I(N__10253));
    Sp12to4 I__2434 (
            .O(N__10265),
            .I(N__10253));
    LocalMux I__2433 (
            .O(N__10262),
            .I(N__10253));
    Span12Mux_h I__2432 (
            .O(N__10253),
            .I(N__10250));
    Odrv12 I__2431 (
            .O(N__10250),
            .I(A_c_1));
    CascadeMux I__2430 (
            .O(N__10247),
            .I(N__10237));
    CascadeMux I__2429 (
            .O(N__10246),
            .I(N__10233));
    InMux I__2428 (
            .O(N__10245),
            .I(N__10230));
    CascadeMux I__2427 (
            .O(N__10244),
            .I(N__10227));
    InMux I__2426 (
            .O(N__10243),
            .I(N__10222));
    InMux I__2425 (
            .O(N__10242),
            .I(N__10222));
    InMux I__2424 (
            .O(N__10241),
            .I(N__10217));
    InMux I__2423 (
            .O(N__10240),
            .I(N__10217));
    InMux I__2422 (
            .O(N__10237),
            .I(N__10214));
    InMux I__2421 (
            .O(N__10236),
            .I(N__10211));
    InMux I__2420 (
            .O(N__10233),
            .I(N__10208));
    LocalMux I__2419 (
            .O(N__10230),
            .I(N__10205));
    InMux I__2418 (
            .O(N__10227),
            .I(N__10202));
    LocalMux I__2417 (
            .O(N__10222),
            .I(N__10193));
    LocalMux I__2416 (
            .O(N__10217),
            .I(N__10193));
    LocalMux I__2415 (
            .O(N__10214),
            .I(N__10193));
    LocalMux I__2414 (
            .O(N__10211),
            .I(N__10193));
    LocalMux I__2413 (
            .O(N__10208),
            .I(N__10190));
    Span4Mux_v I__2412 (
            .O(N__10205),
            .I(N__10185));
    LocalMux I__2411 (
            .O(N__10202),
            .I(N__10185));
    Span4Mux_v I__2410 (
            .O(N__10193),
            .I(N__10182));
    Span4Mux_v I__2409 (
            .O(N__10190),
            .I(N__10179));
    Span4Mux_h I__2408 (
            .O(N__10185),
            .I(N__10176));
    Sp12to4 I__2407 (
            .O(N__10182),
            .I(N__10173));
    Span4Mux_v I__2406 (
            .O(N__10179),
            .I(N__10170));
    Span4Mux_v I__2405 (
            .O(N__10176),
            .I(N__10167));
    Span12Mux_h I__2404 (
            .O(N__10173),
            .I(N__10160));
    Sp12to4 I__2403 (
            .O(N__10170),
            .I(N__10160));
    Sp12to4 I__2402 (
            .O(N__10167),
            .I(N__10160));
    Odrv12 I__2401 (
            .O(N__10160),
            .I(A_c_0));
    InMux I__2400 (
            .O(N__10157),
            .I(N__10151));
    InMux I__2399 (
            .O(N__10156),
            .I(N__10148));
    CascadeMux I__2398 (
            .O(N__10155),
            .I(N__10144));
    CascadeMux I__2397 (
            .O(N__10154),
            .I(N__10140));
    LocalMux I__2396 (
            .O(N__10151),
            .I(N__10134));
    LocalMux I__2395 (
            .O(N__10148),
            .I(N__10134));
    InMux I__2394 (
            .O(N__10147),
            .I(N__10131));
    InMux I__2393 (
            .O(N__10144),
            .I(N__10128));
    InMux I__2392 (
            .O(N__10143),
            .I(N__10123));
    InMux I__2391 (
            .O(N__10140),
            .I(N__10123));
    InMux I__2390 (
            .O(N__10139),
            .I(N__10118));
    Span4Mux_v I__2389 (
            .O(N__10134),
            .I(N__10115));
    LocalMux I__2388 (
            .O(N__10131),
            .I(N__10110));
    LocalMux I__2387 (
            .O(N__10128),
            .I(N__10110));
    LocalMux I__2386 (
            .O(N__10123),
            .I(N__10107));
    InMux I__2385 (
            .O(N__10122),
            .I(N__10102));
    InMux I__2384 (
            .O(N__10121),
            .I(N__10102));
    LocalMux I__2383 (
            .O(N__10118),
            .I(N__10099));
    Span4Mux_v I__2382 (
            .O(N__10115),
            .I(N__10096));
    Span4Mux_v I__2381 (
            .O(N__10110),
            .I(N__10089));
    Span4Mux_h I__2380 (
            .O(N__10107),
            .I(N__10089));
    LocalMux I__2379 (
            .O(N__10102),
            .I(N__10089));
    Span4Mux_v I__2378 (
            .O(N__10099),
            .I(N__10086));
    Span4Mux_v I__2377 (
            .O(N__10096),
            .I(N__10081));
    Span4Mux_h I__2376 (
            .O(N__10089),
            .I(N__10081));
    Span4Mux_v I__2375 (
            .O(N__10086),
            .I(N__10078));
    Span4Mux_v I__2374 (
            .O(N__10081),
            .I(N__10075));
    Span4Mux_v I__2373 (
            .O(N__10078),
            .I(N__10072));
    Span4Mux_h I__2372 (
            .O(N__10075),
            .I(N__10069));
    Sp12to4 I__2371 (
            .O(N__10072),
            .I(N__10064));
    Sp12to4 I__2370 (
            .O(N__10069),
            .I(N__10064));
    Odrv12 I__2369 (
            .O(N__10064),
            .I(SIZ_c_0));
    InMux I__2368 (
            .O(N__10061),
            .I(N__10056));
    InMux I__2367 (
            .O(N__10060),
            .I(N__10052));
    InMux I__2366 (
            .O(N__10059),
            .I(N__10049));
    LocalMux I__2365 (
            .O(N__10056),
            .I(N__10045));
    InMux I__2364 (
            .O(N__10055),
            .I(N__10042));
    LocalMux I__2363 (
            .O(N__10052),
            .I(N__10039));
    LocalMux I__2362 (
            .O(N__10049),
            .I(N__10036));
    CascadeMux I__2361 (
            .O(N__10048),
            .I(N__10032));
    Span4Mux_h I__2360 (
            .O(N__10045),
            .I(N__10027));
    LocalMux I__2359 (
            .O(N__10042),
            .I(N__10027));
    Span4Mux_v I__2358 (
            .O(N__10039),
            .I(N__10024));
    Span4Mux_h I__2357 (
            .O(N__10036),
            .I(N__10021));
    InMux I__2356 (
            .O(N__10035),
            .I(N__10018));
    InMux I__2355 (
            .O(N__10032),
            .I(N__10015));
    Sp12to4 I__2354 (
            .O(N__10027),
            .I(N__10012));
    Span4Mux_v I__2353 (
            .O(N__10024),
            .I(N__10009));
    Span4Mux_v I__2352 (
            .O(N__10021),
            .I(N__10006));
    LocalMux I__2351 (
            .O(N__10018),
            .I(N__10001));
    LocalMux I__2350 (
            .O(N__10015),
            .I(N__10001));
    Span12Mux_v I__2349 (
            .O(N__10012),
            .I(N__9998));
    Sp12to4 I__2348 (
            .O(N__10009),
            .I(N__9991));
    Sp12to4 I__2347 (
            .O(N__10006),
            .I(N__9991));
    Span12Mux_v I__2346 (
            .O(N__10001),
            .I(N__9991));
    Span12Mux_h I__2345 (
            .O(N__9998),
            .I(N__9988));
    Span12Mux_h I__2344 (
            .O(N__9991),
            .I(N__9985));
    Odrv12 I__2343 (
            .O(N__9988),
            .I(SIZ_c_1));
    Odrv12 I__2342 (
            .O(N__9985),
            .I(SIZ_c_1));
    IoInMux I__2341 (
            .O(N__9980),
            .I(N__9977));
    LocalMux I__2340 (
            .O(N__9977),
            .I(N__9974));
    Span4Mux_s3_v I__2339 (
            .O(N__9974),
            .I(N__9971));
    Odrv4 I__2338 (
            .O(N__9971),
            .I(LLBEn_c));
    InMux I__2337 (
            .O(N__9968),
            .I(N__9964));
    InMux I__2336 (
            .O(N__9967),
            .I(N__9960));
    LocalMux I__2335 (
            .O(N__9964),
            .I(N__9955));
    InMux I__2334 (
            .O(N__9963),
            .I(N__9952));
    LocalMux I__2333 (
            .O(N__9960),
            .I(N__9949));
    InMux I__2332 (
            .O(N__9959),
            .I(N__9944));
    InMux I__2331 (
            .O(N__9958),
            .I(N__9944));
    Span4Mux_v I__2330 (
            .O(N__9955),
            .I(N__9939));
    LocalMux I__2329 (
            .O(N__9952),
            .I(N__9939));
    Span4Mux_v I__2328 (
            .O(N__9949),
            .I(N__9934));
    LocalMux I__2327 (
            .O(N__9944),
            .I(N__9934));
    Span4Mux_h I__2326 (
            .O(N__9939),
            .I(N__9930));
    Span4Mux_h I__2325 (
            .O(N__9934),
            .I(N__9927));
    InMux I__2324 (
            .O(N__9933),
            .I(N__9924));
    Odrv4 I__2323 (
            .O(N__9930),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__2322 (
            .O(N__9927),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__2321 (
            .O(N__9924),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__2320 (
            .O(N__9917),
            .I(N__9914));
    LocalMux I__2319 (
            .O(N__9914),
            .I(N__9911));
    Span4Mux_s3_h I__2318 (
            .O(N__9911),
            .I(N__9908));
    Span4Mux_v I__2317 (
            .O(N__9908),
            .I(N__9905));
    Span4Mux_v I__2316 (
            .O(N__9905),
            .I(N__9902));
    Sp12to4 I__2315 (
            .O(N__9902),
            .I(N__9899));
    Odrv12 I__2314 (
            .O(N__9899),
            .I(WEn_c));
    InMux I__2313 (
            .O(N__9896),
            .I(N__9890));
    CascadeMux I__2312 (
            .O(N__9895),
            .I(N__9886));
    InMux I__2311 (
            .O(N__9894),
            .I(N__9883));
    InMux I__2310 (
            .O(N__9893),
            .I(N__9880));
    LocalMux I__2309 (
            .O(N__9890),
            .I(N__9877));
    InMux I__2308 (
            .O(N__9889),
            .I(N__9872));
    InMux I__2307 (
            .O(N__9886),
            .I(N__9872));
    LocalMux I__2306 (
            .O(N__9883),
            .I(N__9869));
    LocalMux I__2305 (
            .O(N__9880),
            .I(N__9866));
    Span4Mux_v I__2304 (
            .O(N__9877),
            .I(N__9861));
    LocalMux I__2303 (
            .O(N__9872),
            .I(N__9861));
    Span4Mux_h I__2302 (
            .O(N__9869),
            .I(N__9855));
    Span4Mux_h I__2301 (
            .O(N__9866),
            .I(N__9855));
    Span4Mux_h I__2300 (
            .O(N__9861),
            .I(N__9852));
    InMux I__2299 (
            .O(N__9860),
            .I(N__9849));
    Odrv4 I__2298 (
            .O(N__9855),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__2297 (
            .O(N__9852),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__2296 (
            .O(N__9849),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    IoInMux I__2295 (
            .O(N__9842),
            .I(N__9839));
    LocalMux I__2294 (
            .O(N__9839),
            .I(N__9836));
    Span4Mux_s1_v I__2293 (
            .O(N__9836),
            .I(N__9833));
    Span4Mux_v I__2292 (
            .O(N__9833),
            .I(N__9830));
    Span4Mux_v I__2291 (
            .O(N__9830),
            .I(N__9827));
    Span4Mux_h I__2290 (
            .O(N__9827),
            .I(N__9824));
    Odrv4 I__2289 (
            .O(N__9824),
            .I(RASn_c));
    InMux I__2288 (
            .O(N__9821),
            .I(N__9818));
    LocalMux I__2287 (
            .O(N__9818),
            .I(N__9797));
    ClkMux I__2286 (
            .O(N__9817),
            .I(N__9713));
    ClkMux I__2285 (
            .O(N__9816),
            .I(N__9713));
    ClkMux I__2284 (
            .O(N__9815),
            .I(N__9713));
    ClkMux I__2283 (
            .O(N__9814),
            .I(N__9713));
    ClkMux I__2282 (
            .O(N__9813),
            .I(N__9713));
    ClkMux I__2281 (
            .O(N__9812),
            .I(N__9713));
    ClkMux I__2280 (
            .O(N__9811),
            .I(N__9713));
    ClkMux I__2279 (
            .O(N__9810),
            .I(N__9713));
    ClkMux I__2278 (
            .O(N__9809),
            .I(N__9713));
    ClkMux I__2277 (
            .O(N__9808),
            .I(N__9713));
    ClkMux I__2276 (
            .O(N__9807),
            .I(N__9713));
    ClkMux I__2275 (
            .O(N__9806),
            .I(N__9713));
    ClkMux I__2274 (
            .O(N__9805),
            .I(N__9713));
    ClkMux I__2273 (
            .O(N__9804),
            .I(N__9713));
    ClkMux I__2272 (
            .O(N__9803),
            .I(N__9713));
    ClkMux I__2271 (
            .O(N__9802),
            .I(N__9713));
    ClkMux I__2270 (
            .O(N__9801),
            .I(N__9713));
    ClkMux I__2269 (
            .O(N__9800),
            .I(N__9713));
    Glb2LocalMux I__2268 (
            .O(N__9797),
            .I(N__9713));
    ClkMux I__2267 (
            .O(N__9796),
            .I(N__9713));
    ClkMux I__2266 (
            .O(N__9795),
            .I(N__9713));
    ClkMux I__2265 (
            .O(N__9794),
            .I(N__9713));
    ClkMux I__2264 (
            .O(N__9793),
            .I(N__9713));
    ClkMux I__2263 (
            .O(N__9792),
            .I(N__9713));
    ClkMux I__2262 (
            .O(N__9791),
            .I(N__9713));
    ClkMux I__2261 (
            .O(N__9790),
            .I(N__9713));
    ClkMux I__2260 (
            .O(N__9789),
            .I(N__9713));
    ClkMux I__2259 (
            .O(N__9788),
            .I(N__9713));
    ClkMux I__2258 (
            .O(N__9787),
            .I(N__9713));
    ClkMux I__2257 (
            .O(N__9786),
            .I(N__9713));
    ClkMux I__2256 (
            .O(N__9785),
            .I(N__9713));
    ClkMux I__2255 (
            .O(N__9784),
            .I(N__9713));
    ClkMux I__2254 (
            .O(N__9783),
            .I(N__9713));
    ClkMux I__2253 (
            .O(N__9782),
            .I(N__9713));
    GlobalMux I__2252 (
            .O(N__9713),
            .I(CLK80_PLL));
    CascadeMux I__2251 (
            .O(N__9710),
            .I(N__9700));
    InMux I__2250 (
            .O(N__9709),
            .I(N__9696));
    CascadeMux I__2249 (
            .O(N__9708),
            .I(N__9691));
    InMux I__2248 (
            .O(N__9707),
            .I(N__9686));
    InMux I__2247 (
            .O(N__9706),
            .I(N__9683));
    InMux I__2246 (
            .O(N__9705),
            .I(N__9678));
    InMux I__2245 (
            .O(N__9704),
            .I(N__9675));
    InMux I__2244 (
            .O(N__9703),
            .I(N__9670));
    InMux I__2243 (
            .O(N__9700),
            .I(N__9665));
    InMux I__2242 (
            .O(N__9699),
            .I(N__9665));
    LocalMux I__2241 (
            .O(N__9696),
            .I(N__9662));
    CascadeMux I__2240 (
            .O(N__9695),
            .I(N__9658));
    InMux I__2239 (
            .O(N__9694),
            .I(N__9653));
    InMux I__2238 (
            .O(N__9691),
            .I(N__9646));
    InMux I__2237 (
            .O(N__9690),
            .I(N__9646));
    InMux I__2236 (
            .O(N__9689),
            .I(N__9646));
    LocalMux I__2235 (
            .O(N__9686),
            .I(N__9639));
    LocalMux I__2234 (
            .O(N__9683),
            .I(N__9639));
    CascadeMux I__2233 (
            .O(N__9682),
            .I(N__9634));
    InMux I__2232 (
            .O(N__9681),
            .I(N__9631));
    LocalMux I__2231 (
            .O(N__9678),
            .I(N__9626));
    LocalMux I__2230 (
            .O(N__9675),
            .I(N__9626));
    InMux I__2229 (
            .O(N__9674),
            .I(N__9621));
    InMux I__2228 (
            .O(N__9673),
            .I(N__9621));
    LocalMux I__2227 (
            .O(N__9670),
            .I(N__9618));
    LocalMux I__2226 (
            .O(N__9665),
            .I(N__9613));
    Span4Mux_v I__2225 (
            .O(N__9662),
            .I(N__9613));
    InMux I__2224 (
            .O(N__9661),
            .I(N__9608));
    InMux I__2223 (
            .O(N__9658),
            .I(N__9608));
    InMux I__2222 (
            .O(N__9657),
            .I(N__9603));
    InMux I__2221 (
            .O(N__9656),
            .I(N__9603));
    LocalMux I__2220 (
            .O(N__9653),
            .I(N__9598));
    LocalMux I__2219 (
            .O(N__9646),
            .I(N__9598));
    InMux I__2218 (
            .O(N__9645),
            .I(N__9595));
    InMux I__2217 (
            .O(N__9644),
            .I(N__9592));
    Span4Mux_v I__2216 (
            .O(N__9639),
            .I(N__9589));
    InMux I__2215 (
            .O(N__9638),
            .I(N__9586));
    InMux I__2214 (
            .O(N__9637),
            .I(N__9581));
    InMux I__2213 (
            .O(N__9634),
            .I(N__9581));
    LocalMux I__2212 (
            .O(N__9631),
            .I(N__9578));
    Span12Mux_v I__2211 (
            .O(N__9626),
            .I(N__9573));
    LocalMux I__2210 (
            .O(N__9621),
            .I(N__9573));
    Span4Mux_v I__2209 (
            .O(N__9618),
            .I(N__9568));
    Span4Mux_h I__2208 (
            .O(N__9613),
            .I(N__9568));
    LocalMux I__2207 (
            .O(N__9608),
            .I(N__9561));
    LocalMux I__2206 (
            .O(N__9603),
            .I(N__9561));
    Span4Mux_v I__2205 (
            .O(N__9598),
            .I(N__9561));
    LocalMux I__2204 (
            .O(N__9595),
            .I(N__9556));
    LocalMux I__2203 (
            .O(N__9592),
            .I(N__9556));
    Odrv4 I__2202 (
            .O(N__9589),
            .I(CPU_CYCLEm));
    LocalMux I__2201 (
            .O(N__9586),
            .I(CPU_CYCLEm));
    LocalMux I__2200 (
            .O(N__9581),
            .I(CPU_CYCLEm));
    Odrv4 I__2199 (
            .O(N__9578),
            .I(CPU_CYCLEm));
    Odrv12 I__2198 (
            .O(N__9573),
            .I(CPU_CYCLEm));
    Odrv4 I__2197 (
            .O(N__9568),
            .I(CPU_CYCLEm));
    Odrv4 I__2196 (
            .O(N__9561),
            .I(CPU_CYCLEm));
    Odrv12 I__2195 (
            .O(N__9556),
            .I(CPU_CYCLEm));
    InMux I__2194 (
            .O(N__9539),
            .I(N__9536));
    LocalMux I__2193 (
            .O(N__9536),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ));
    CascadeMux I__2192 (
            .O(N__9533),
            .I(N__9528));
    InMux I__2191 (
            .O(N__9532),
            .I(N__9516));
    CascadeMux I__2190 (
            .O(N__9531),
            .I(N__9513));
    InMux I__2189 (
            .O(N__9528),
            .I(N__9509));
    CascadeMux I__2188 (
            .O(N__9527),
            .I(N__9506));
    CascadeMux I__2187 (
            .O(N__9526),
            .I(N__9503));
    InMux I__2186 (
            .O(N__9525),
            .I(N__9499));
    CascadeMux I__2185 (
            .O(N__9524),
            .I(N__9495));
    InMux I__2184 (
            .O(N__9523),
            .I(N__9489));
    InMux I__2183 (
            .O(N__9522),
            .I(N__9484));
    InMux I__2182 (
            .O(N__9521),
            .I(N__9484));
    InMux I__2181 (
            .O(N__9520),
            .I(N__9479));
    InMux I__2180 (
            .O(N__9519),
            .I(N__9479));
    LocalMux I__2179 (
            .O(N__9516),
            .I(N__9476));
    InMux I__2178 (
            .O(N__9513),
            .I(N__9471));
    InMux I__2177 (
            .O(N__9512),
            .I(N__9471));
    LocalMux I__2176 (
            .O(N__9509),
            .I(N__9468));
    InMux I__2175 (
            .O(N__9506),
            .I(N__9465));
    InMux I__2174 (
            .O(N__9503),
            .I(N__9461));
    InMux I__2173 (
            .O(N__9502),
            .I(N__9458));
    LocalMux I__2172 (
            .O(N__9499),
            .I(N__9455));
    InMux I__2171 (
            .O(N__9498),
            .I(N__9448));
    InMux I__2170 (
            .O(N__9495),
            .I(N__9448));
    InMux I__2169 (
            .O(N__9494),
            .I(N__9448));
    InMux I__2168 (
            .O(N__9493),
            .I(N__9443));
    InMux I__2167 (
            .O(N__9492),
            .I(N__9443));
    LocalMux I__2166 (
            .O(N__9489),
            .I(N__9437));
    LocalMux I__2165 (
            .O(N__9484),
            .I(N__9437));
    LocalMux I__2164 (
            .O(N__9479),
            .I(N__9432));
    Span4Mux_v I__2163 (
            .O(N__9476),
            .I(N__9432));
    LocalMux I__2162 (
            .O(N__9471),
            .I(N__9427));
    Span4Mux_h I__2161 (
            .O(N__9468),
            .I(N__9427));
    LocalMux I__2160 (
            .O(N__9465),
            .I(N__9424));
    InMux I__2159 (
            .O(N__9464),
            .I(N__9421));
    LocalMux I__2158 (
            .O(N__9461),
            .I(N__9406));
    LocalMux I__2157 (
            .O(N__9458),
            .I(N__9406));
    Span4Mux_h I__2156 (
            .O(N__9455),
            .I(N__9406));
    LocalMux I__2155 (
            .O(N__9448),
            .I(N__9406));
    LocalMux I__2154 (
            .O(N__9443),
            .I(N__9406));
    InMux I__2153 (
            .O(N__9442),
            .I(N__9403));
    Span4Mux_v I__2152 (
            .O(N__9437),
            .I(N__9400));
    Span4Mux_h I__2151 (
            .O(N__9432),
            .I(N__9397));
    Span4Mux_h I__2150 (
            .O(N__9427),
            .I(N__9394));
    Span4Mux_h I__2149 (
            .O(N__9424),
            .I(N__9389));
    LocalMux I__2148 (
            .O(N__9421),
            .I(N__9389));
    InMux I__2147 (
            .O(N__9420),
            .I(N__9382));
    InMux I__2146 (
            .O(N__9419),
            .I(N__9382));
    InMux I__2145 (
            .O(N__9418),
            .I(N__9382));
    InMux I__2144 (
            .O(N__9417),
            .I(N__9379));
    Span4Mux_v I__2143 (
            .O(N__9406),
            .I(N__9374));
    LocalMux I__2142 (
            .O(N__9403),
            .I(N__9374));
    Odrv4 I__2141 (
            .O(N__9400),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2140 (
            .O(N__9397),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2139 (
            .O(N__9394),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2138 (
            .O(N__9389),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2137 (
            .O(N__9382),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2136 (
            .O(N__9379),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2135 (
            .O(N__9374),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    InMux I__2134 (
            .O(N__9359),
            .I(N__9356));
    LocalMux I__2133 (
            .O(N__9356),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    InMux I__2132 (
            .O(N__9353),
            .I(N__9350));
    LocalMux I__2131 (
            .O(N__9350),
            .I(N__9347));
    Span4Mux_h I__2130 (
            .O(N__9347),
            .I(N__9344));
    Odrv4 I__2129 (
            .O(N__9344),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__2128 (
            .O(N__9341),
            .I(N__9338));
    LocalMux I__2127 (
            .O(N__9338),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__2126 (
            .O(N__9335),
            .I(N__9332));
    LocalMux I__2125 (
            .O(N__9332),
            .I(N__9329));
    Span4Mux_h I__2124 (
            .O(N__9329),
            .I(N__9326));
    Odrv4 I__2123 (
            .O(N__9326),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__2122 (
            .O(N__9323),
            .I(N__9316));
    InMux I__2121 (
            .O(N__9322),
            .I(N__9316));
    InMux I__2120 (
            .O(N__9321),
            .I(N__9313));
    LocalMux I__2119 (
            .O(N__9316),
            .I(N__9310));
    LocalMux I__2118 (
            .O(N__9313),
            .I(N__9307));
    Span4Mux_v I__2117 (
            .O(N__9310),
            .I(N__9303));
    Span4Mux_h I__2116 (
            .O(N__9307),
            .I(N__9300));
    InMux I__2115 (
            .O(N__9306),
            .I(N__9297));
    Span4Mux_v I__2114 (
            .O(N__9303),
            .I(N__9294));
    Span4Mux_v I__2113 (
            .O(N__9300),
            .I(N__9291));
    LocalMux I__2112 (
            .O(N__9297),
            .I(N__9288));
    Sp12to4 I__2111 (
            .O(N__9294),
            .I(N__9281));
    Sp12to4 I__2110 (
            .O(N__9291),
            .I(N__9281));
    Span12Mux_v I__2109 (
            .O(N__9288),
            .I(N__9281));
    Span12Mux_h I__2108 (
            .O(N__9281),
            .I(N__9278));
    Odrv12 I__2107 (
            .O(N__9278),
            .I(DRA_c_6));
    InMux I__2106 (
            .O(N__9275),
            .I(N__9271));
    InMux I__2105 (
            .O(N__9274),
            .I(N__9268));
    LocalMux I__2104 (
            .O(N__9271),
            .I(N__9262));
    LocalMux I__2103 (
            .O(N__9268),
            .I(N__9262));
    InMux I__2102 (
            .O(N__9267),
            .I(N__9259));
    Span4Mux_v I__2101 (
            .O(N__9262),
            .I(N__9255));
    LocalMux I__2100 (
            .O(N__9259),
            .I(N__9252));
    InMux I__2099 (
            .O(N__9258),
            .I(N__9249));
    Span4Mux_v I__2098 (
            .O(N__9255),
            .I(N__9246));
    Sp12to4 I__2097 (
            .O(N__9252),
            .I(N__9241));
    LocalMux I__2096 (
            .O(N__9249),
            .I(N__9241));
    Sp12to4 I__2095 (
            .O(N__9246),
            .I(N__9236));
    Span12Mux_v I__2094 (
            .O(N__9241),
            .I(N__9236));
    Span12Mux_h I__2093 (
            .O(N__9236),
            .I(N__9233));
    Odrv12 I__2092 (
            .O(N__9233),
            .I(DRA_c_5));
    InMux I__2091 (
            .O(N__9230),
            .I(N__9227));
    LocalMux I__2090 (
            .O(N__9227),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__2089 (
            .O(N__9224),
            .I(N__9220));
    InMux I__2088 (
            .O(N__9223),
            .I(N__9217));
    LocalMux I__2087 (
            .O(N__9220),
            .I(N__9211));
    LocalMux I__2086 (
            .O(N__9217),
            .I(N__9211));
    InMux I__2085 (
            .O(N__9216),
            .I(N__9208));
    Span4Mux_v I__2084 (
            .O(N__9211),
            .I(N__9204));
    LocalMux I__2083 (
            .O(N__9208),
            .I(N__9201));
    InMux I__2082 (
            .O(N__9207),
            .I(N__9198));
    Sp12to4 I__2081 (
            .O(N__9204),
            .I(N__9193));
    Span12Mux_v I__2080 (
            .O(N__9201),
            .I(N__9193));
    LocalMux I__2079 (
            .O(N__9198),
            .I(N__9190));
    Span12Mux_h I__2078 (
            .O(N__9193),
            .I(N__9187));
    Span12Mux_h I__2077 (
            .O(N__9190),
            .I(N__9184));
    Odrv12 I__2076 (
            .O(N__9187),
            .I(DRA_c_8));
    Odrv12 I__2075 (
            .O(N__9184),
            .I(DRA_c_8));
    InMux I__2074 (
            .O(N__9179),
            .I(N__9176));
    LocalMux I__2073 (
            .O(N__9176),
            .I(N__9173));
    Odrv4 I__2072 (
            .O(N__9173),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__2071 (
            .O(N__9170),
            .I(N__9167));
    LocalMux I__2070 (
            .O(N__9167),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    CascadeMux I__2069 (
            .O(N__9164),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_ ));
    InMux I__2068 (
            .O(N__9161),
            .I(N__9158));
    LocalMux I__2067 (
            .O(N__9158),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ));
    IoInMux I__2066 (
            .O(N__9155),
            .I(N__9152));
    LocalMux I__2065 (
            .O(N__9152),
            .I(N__9149));
    IoSpan4Mux I__2064 (
            .O(N__9149),
            .I(N__9146));
    Span4Mux_s3_v I__2063 (
            .O(N__9146),
            .I(N__9143));
    Span4Mux_v I__2062 (
            .O(N__9143),
            .I(N__9140));
    Odrv4 I__2061 (
            .O(N__9140),
            .I(CMA_c_1));
    CEMux I__2060 (
            .O(N__9137),
            .I(N__9134));
    LocalMux I__2059 (
            .O(N__9134),
            .I(N__9131));
    Span4Mux_h I__2058 (
            .O(N__9131),
            .I(N__9124));
    CEMux I__2057 (
            .O(N__9130),
            .I(N__9121));
    CEMux I__2056 (
            .O(N__9129),
            .I(N__9118));
    CEMux I__2055 (
            .O(N__9128),
            .I(N__9115));
    CEMux I__2054 (
            .O(N__9127),
            .I(N__9112));
    Odrv4 I__2053 (
            .O(N__9124),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    LocalMux I__2052 (
            .O(N__9121),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    LocalMux I__2051 (
            .O(N__9118),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    LocalMux I__2050 (
            .O(N__9115),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    LocalMux I__2049 (
            .O(N__9112),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    InMux I__2048 (
            .O(N__9101),
            .I(N__9098));
    LocalMux I__2047 (
            .O(N__9098),
            .I(N__9095));
    Span4Mux_v I__2046 (
            .O(N__9095),
            .I(N__9092));
    Sp12to4 I__2045 (
            .O(N__9092),
            .I(N__9089));
    Span12Mux_h I__2044 (
            .O(N__9089),
            .I(N__9086));
    Odrv12 I__2043 (
            .O(N__9086),
            .I(A_c_13));
    InMux I__2042 (
            .O(N__9083),
            .I(N__9080));
    LocalMux I__2041 (
            .O(N__9080),
            .I(N__9077));
    Sp12to4 I__2040 (
            .O(N__9077),
            .I(N__9074));
    Span12Mux_v I__2039 (
            .O(N__9074),
            .I(N__9071));
    Span12Mux_h I__2038 (
            .O(N__9071),
            .I(N__9068));
    Odrv12 I__2037 (
            .O(N__9068),
            .I(A_c_6));
    InMux I__2036 (
            .O(N__9065),
            .I(N__9062));
    LocalMux I__2035 (
            .O(N__9062),
            .I(N__9059));
    Span4Mux_h I__2034 (
            .O(N__9059),
            .I(N__9056));
    Odrv4 I__2033 (
            .O(N__9056),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    CascadeMux I__2032 (
            .O(N__9053),
            .I(N__9050));
    InMux I__2031 (
            .O(N__9050),
            .I(N__9047));
    LocalMux I__2030 (
            .O(N__9047),
            .I(N__9044));
    Odrv4 I__2029 (
            .O(N__9044),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__2028 (
            .O(N__9041),
            .I(N__9036));
    InMux I__2027 (
            .O(N__9040),
            .I(N__9033));
    InMux I__2026 (
            .O(N__9039),
            .I(N__9030));
    LocalMux I__2025 (
            .O(N__9036),
            .I(N__9027));
    LocalMux I__2024 (
            .O(N__9033),
            .I(N__9019));
    LocalMux I__2023 (
            .O(N__9030),
            .I(N__9019));
    Span4Mux_h I__2022 (
            .O(N__9027),
            .I(N__9019));
    InMux I__2021 (
            .O(N__9026),
            .I(N__9016));
    Sp12to4 I__2020 (
            .O(N__9019),
            .I(N__9011));
    LocalMux I__2019 (
            .O(N__9016),
            .I(N__9011));
    Span12Mux_v I__2018 (
            .O(N__9011),
            .I(N__9008));
    Span12Mux_h I__2017 (
            .O(N__9008),
            .I(N__9005));
    Odrv12 I__2016 (
            .O(N__9005),
            .I(DRA_c_7));
    InMux I__2015 (
            .O(N__9002),
            .I(N__8999));
    LocalMux I__2014 (
            .O(N__8999),
            .I(N__8996));
    Span4Mux_h I__2013 (
            .O(N__8996),
            .I(N__8993));
    Odrv4 I__2012 (
            .O(N__8993),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2011 (
            .O(N__8990),
            .I(N__8987));
    LocalMux I__2010 (
            .O(N__8987),
            .I(N__8984));
    Span4Mux_v I__2009 (
            .O(N__8984),
            .I(N__8981));
    Span4Mux_h I__2008 (
            .O(N__8981),
            .I(N__8978));
    Odrv4 I__2007 (
            .O(N__8978),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    InMux I__2006 (
            .O(N__8975),
            .I(N__8972));
    LocalMux I__2005 (
            .O(N__8972),
            .I(N__8969));
    Span4Mux_h I__2004 (
            .O(N__8969),
            .I(N__8966));
    Span4Mux_v I__2003 (
            .O(N__8966),
            .I(N__8963));
    Odrv4 I__2002 (
            .O(N__8963),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__2001 (
            .O(N__8960),
            .I(N__8957));
    LocalMux I__2000 (
            .O(N__8957),
            .I(N__8953));
    InMux I__1999 (
            .O(N__8956),
            .I(N__8950));
    Span4Mux_v I__1998 (
            .O(N__8953),
            .I(N__8945));
    LocalMux I__1997 (
            .O(N__8950),
            .I(N__8945));
    Span4Mux_h I__1996 (
            .O(N__8945),
            .I(N__8942));
    Sp12to4 I__1995 (
            .O(N__8942),
            .I(N__8939));
    Span12Mux_h I__1994 (
            .O(N__8939),
            .I(N__8936));
    Span12Mux_v I__1993 (
            .O(N__8936),
            .I(N__8933));
    Odrv12 I__1992 (
            .O(N__8933),
            .I(DRA_c_0));
    InMux I__1991 (
            .O(N__8930),
            .I(N__8927));
    LocalMux I__1990 (
            .O(N__8927),
            .I(N__8924));
    Odrv12 I__1989 (
            .O(N__8924),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    IoInMux I__1988 (
            .O(N__8921),
            .I(N__8918));
    LocalMux I__1987 (
            .O(N__8918),
            .I(N__8915));
    Span4Mux_s3_v I__1986 (
            .O(N__8915),
            .I(N__8912));
    Span4Mux_v I__1985 (
            .O(N__8912),
            .I(N__8909));
    Sp12to4 I__1984 (
            .O(N__8909),
            .I(N__8906));
    Span12Mux_h I__1983 (
            .O(N__8906),
            .I(N__8903));
    Odrv12 I__1982 (
            .O(N__8903),
            .I(CASn_c));
    InMux I__1981 (
            .O(N__8900),
            .I(N__8897));
    LocalMux I__1980 (
            .O(N__8897),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    IoInMux I__1979 (
            .O(N__8894),
            .I(N__8891));
    LocalMux I__1978 (
            .O(N__8891),
            .I(N__8888));
    Span4Mux_s2_v I__1977 (
            .O(N__8888),
            .I(N__8885));
    Span4Mux_v I__1976 (
            .O(N__8885),
            .I(N__8882));
    Span4Mux_h I__1975 (
            .O(N__8882),
            .I(N__8879));
    Odrv4 I__1974 (
            .O(N__8879),
            .I(CMA_c_0));
    InMux I__1973 (
            .O(N__8876),
            .I(N__8872));
    InMux I__1972 (
            .O(N__8875),
            .I(N__8868));
    LocalMux I__1971 (
            .O(N__8872),
            .I(N__8865));
    InMux I__1970 (
            .O(N__8871),
            .I(N__8862));
    LocalMux I__1969 (
            .O(N__8868),
            .I(N__8856));
    Span4Mux_v I__1968 (
            .O(N__8865),
            .I(N__8856));
    LocalMux I__1967 (
            .O(N__8862),
            .I(N__8853));
    CascadeMux I__1966 (
            .O(N__8861),
            .I(N__8850));
    Span4Mux_v I__1965 (
            .O(N__8856),
            .I(N__8847));
    Span12Mux_h I__1964 (
            .O(N__8853),
            .I(N__8844));
    InMux I__1963 (
            .O(N__8850),
            .I(N__8841));
    Odrv4 I__1962 (
            .O(N__8847),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv12 I__1961 (
            .O(N__8844),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1960 (
            .O(N__8841),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__1959 (
            .O(N__8834),
            .I(N__8831));
    LocalMux I__1958 (
            .O(N__8831),
            .I(N__8828));
    Span12Mux_s10_v I__1957 (
            .O(N__8828),
            .I(N__8825));
    Odrv12 I__1956 (
            .O(N__8825),
            .I(CMA_c_10));
    InMux I__1955 (
            .O(N__8822),
            .I(N__8819));
    LocalMux I__1954 (
            .O(N__8819),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ));
    InMux I__1953 (
            .O(N__8816),
            .I(N__8813));
    LocalMux I__1952 (
            .O(N__8813),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ));
    InMux I__1951 (
            .O(N__8810),
            .I(N__8807));
    LocalMux I__1950 (
            .O(N__8807),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ));
    IoInMux I__1949 (
            .O(N__8804),
            .I(N__8801));
    LocalMux I__1948 (
            .O(N__8801),
            .I(N__8798));
    IoSpan4Mux I__1947 (
            .O(N__8798),
            .I(N__8795));
    Span4Mux_s2_h I__1946 (
            .O(N__8795),
            .I(N__8792));
    Sp12to4 I__1945 (
            .O(N__8792),
            .I(N__8789));
    Span12Mux_h I__1944 (
            .O(N__8789),
            .I(N__8786));
    Odrv12 I__1943 (
            .O(N__8786),
            .I(CMA_c_5));
    CascadeMux I__1942 (
            .O(N__8783),
            .I(N__8778));
    CascadeMux I__1941 (
            .O(N__8782),
            .I(N__8775));
    CascadeMux I__1940 (
            .O(N__8781),
            .I(N__8772));
    InMux I__1939 (
            .O(N__8778),
            .I(N__8767));
    InMux I__1938 (
            .O(N__8775),
            .I(N__8763));
    InMux I__1937 (
            .O(N__8772),
            .I(N__8760));
    InMux I__1936 (
            .O(N__8771),
            .I(N__8752));
    InMux I__1935 (
            .O(N__8770),
            .I(N__8752));
    LocalMux I__1934 (
            .O(N__8767),
            .I(N__8749));
    InMux I__1933 (
            .O(N__8766),
            .I(N__8746));
    LocalMux I__1932 (
            .O(N__8763),
            .I(N__8743));
    LocalMux I__1931 (
            .O(N__8760),
            .I(N__8740));
    InMux I__1930 (
            .O(N__8759),
            .I(N__8733));
    InMux I__1929 (
            .O(N__8758),
            .I(N__8733));
    InMux I__1928 (
            .O(N__8757),
            .I(N__8733));
    LocalMux I__1927 (
            .O(N__8752),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__1926 (
            .O(N__8749),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__1925 (
            .O(N__8746),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__1924 (
            .O(N__8743),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__1923 (
            .O(N__8740),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__1922 (
            .O(N__8733),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    InMux I__1921 (
            .O(N__8720),
            .I(N__8712));
    InMux I__1920 (
            .O(N__8719),
            .I(N__8707));
    InMux I__1919 (
            .O(N__8718),
            .I(N__8707));
    InMux I__1918 (
            .O(N__8717),
            .I(N__8704));
    InMux I__1917 (
            .O(N__8716),
            .I(N__8699));
    InMux I__1916 (
            .O(N__8715),
            .I(N__8699));
    LocalMux I__1915 (
            .O(N__8712),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9 ));
    LocalMux I__1914 (
            .O(N__8707),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9 ));
    LocalMux I__1913 (
            .O(N__8704),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9 ));
    LocalMux I__1912 (
            .O(N__8699),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9 ));
    IoInMux I__1911 (
            .O(N__8690),
            .I(N__8687));
    LocalMux I__1910 (
            .O(N__8687),
            .I(N__8684));
    Span4Mux_s3_h I__1909 (
            .O(N__8684),
            .I(N__8681));
    Sp12to4 I__1908 (
            .O(N__8681),
            .I(N__8678));
    Span12Mux_s9_v I__1907 (
            .O(N__8678),
            .I(N__8675));
    Span12Mux_h I__1906 (
            .O(N__8675),
            .I(N__8672));
    Odrv12 I__1905 (
            .O(N__8672),
            .I(CMA_c_4));
    InMux I__1904 (
            .O(N__8669),
            .I(N__8666));
    LocalMux I__1903 (
            .O(N__8666),
            .I(N__8663));
    Span4Mux_v I__1902 (
            .O(N__8663),
            .I(N__8660));
    Span4Mux_v I__1901 (
            .O(N__8660),
            .I(N__8657));
    Sp12to4 I__1900 (
            .O(N__8657),
            .I(N__8654));
    Span12Mux_h I__1899 (
            .O(N__8654),
            .I(N__8651));
    Odrv12 I__1898 (
            .O(N__8651),
            .I(A_c_19));
    IoInMux I__1897 (
            .O(N__8648),
            .I(N__8645));
    LocalMux I__1896 (
            .O(N__8645),
            .I(N__8642));
    IoSpan4Mux I__1895 (
            .O(N__8642),
            .I(N__8639));
    Span4Mux_s2_h I__1894 (
            .O(N__8639),
            .I(N__8636));
    Sp12to4 I__1893 (
            .O(N__8636),
            .I(N__8633));
    Span12Mux_h I__1892 (
            .O(N__8633),
            .I(N__8630));
    Odrv12 I__1891 (
            .O(N__8630),
            .I(CMA_c_9));
    CascadeMux I__1890 (
            .O(N__8627),
            .I(N__8624));
    InMux I__1889 (
            .O(N__8624),
            .I(N__8621));
    LocalMux I__1888 (
            .O(N__8621),
            .I(N__8618));
    Span4Mux_h I__1887 (
            .O(N__8618),
            .I(N__8615));
    Sp12to4 I__1886 (
            .O(N__8615),
            .I(N__8612));
    Span12Mux_v I__1885 (
            .O(N__8612),
            .I(N__8609));
    Span12Mux_h I__1884 (
            .O(N__8609),
            .I(N__8606));
    Odrv12 I__1883 (
            .O(N__8606),
            .I(A_c_17));
    CascadeMux I__1882 (
            .O(N__8603),
            .I(N__8598));
    CascadeMux I__1881 (
            .O(N__8602),
            .I(N__8595));
    InMux I__1880 (
            .O(N__8601),
            .I(N__8590));
    InMux I__1879 (
            .O(N__8598),
            .I(N__8590));
    InMux I__1878 (
            .O(N__8595),
            .I(N__8587));
    LocalMux I__1877 (
            .O(N__8590),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    LocalMux I__1876 (
            .O(N__8587),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    IoInMux I__1875 (
            .O(N__8582),
            .I(N__8579));
    LocalMux I__1874 (
            .O(N__8579),
            .I(N__8576));
    Span4Mux_s3_h I__1873 (
            .O(N__8576),
            .I(N__8573));
    Sp12to4 I__1872 (
            .O(N__8573),
            .I(N__8570));
    Span12Mux_v I__1871 (
            .O(N__8570),
            .I(N__8567));
    Span12Mux_h I__1870 (
            .O(N__8567),
            .I(N__8564));
    Odrv12 I__1869 (
            .O(N__8564),
            .I(CMA_c_8));
    InMux I__1868 (
            .O(N__8561),
            .I(N__8558));
    LocalMux I__1867 (
            .O(N__8558),
            .I(N__8555));
    Span4Mux_v I__1866 (
            .O(N__8555),
            .I(N__8552));
    Sp12to4 I__1865 (
            .O(N__8552),
            .I(N__8549));
    Span12Mux_h I__1864 (
            .O(N__8549),
            .I(N__8546));
    Span12Mux_v I__1863 (
            .O(N__8546),
            .I(N__8543));
    Odrv12 I__1862 (
            .O(N__8543),
            .I(A_c_3));
    InMux I__1861 (
            .O(N__8540),
            .I(N__8537));
    LocalMux I__1860 (
            .O(N__8537),
            .I(N__8534));
    Span12Mux_h I__1859 (
            .O(N__8534),
            .I(N__8531));
    Odrv12 I__1858 (
            .O(N__8531),
            .I(A_c_10));
    CascadeMux I__1857 (
            .O(N__8528),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ));
    InMux I__1856 (
            .O(N__8525),
            .I(N__8519));
    InMux I__1855 (
            .O(N__8524),
            .I(N__8519));
    LocalMux I__1854 (
            .O(N__8519),
            .I(N__8516));
    Odrv4 I__1853 (
            .O(N__8516),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__1852 (
            .O(N__8513),
            .I(N__8510));
    LocalMux I__1851 (
            .O(N__8510),
            .I(N__8507));
    Span4Mux_h I__1850 (
            .O(N__8507),
            .I(N__8504));
    Odrv4 I__1849 (
            .O(N__8504),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__1848 (
            .O(N__8501),
            .I(N__8498));
    LocalMux I__1847 (
            .O(N__8498),
            .I(N__8495));
    Odrv4 I__1846 (
            .O(N__8495),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__1845 (
            .O(N__8492),
            .I(N__8489));
    LocalMux I__1844 (
            .O(N__8489),
            .I(N__8486));
    Odrv4 I__1843 (
            .O(N__8486),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    CascadeMux I__1842 (
            .O(N__8483),
            .I(N__8478));
    CascadeMux I__1841 (
            .O(N__8482),
            .I(N__8475));
    InMux I__1840 (
            .O(N__8481),
            .I(N__8467));
    InMux I__1839 (
            .O(N__8478),
            .I(N__8467));
    InMux I__1838 (
            .O(N__8475),
            .I(N__8467));
    InMux I__1837 (
            .O(N__8474),
            .I(N__8464));
    LocalMux I__1836 (
            .O(N__8467),
            .I(N__8461));
    LocalMux I__1835 (
            .O(N__8464),
            .I(N__8458));
    Span4Mux_v I__1834 (
            .O(N__8461),
            .I(N__8455));
    Span4Mux_v I__1833 (
            .O(N__8458),
            .I(N__8450));
    Span4Mux_h I__1832 (
            .O(N__8455),
            .I(N__8450));
    Span4Mux_v I__1831 (
            .O(N__8450),
            .I(N__8447));
    Span4Mux_v I__1830 (
            .O(N__8447),
            .I(N__8444));
    Odrv4 I__1829 (
            .O(N__8444),
            .I(CLK40_PLL_i));
    IoInMux I__1828 (
            .O(N__8441),
            .I(N__8437));
    IoInMux I__1827 (
            .O(N__8440),
            .I(N__8434));
    LocalMux I__1826 (
            .O(N__8437),
            .I(N__8431));
    LocalMux I__1825 (
            .O(N__8434),
            .I(N__8428));
    Span4Mux_s0_v I__1824 (
            .O(N__8431),
            .I(N__8425));
    Span4Mux_s0_v I__1823 (
            .O(N__8428),
            .I(N__8422));
    Span4Mux_v I__1822 (
            .O(N__8425),
            .I(N__8419));
    Span4Mux_v I__1821 (
            .O(N__8422),
            .I(N__8416));
    Sp12to4 I__1820 (
            .O(N__8419),
            .I(N__8410));
    Sp12to4 I__1819 (
            .O(N__8416),
            .I(N__8410));
    IoInMux I__1818 (
            .O(N__8415),
            .I(N__8407));
    Span12Mux_h I__1817 (
            .O(N__8410),
            .I(N__8404));
    LocalMux I__1816 (
            .O(N__8407),
            .I(N__8401));
    Span12Mux_v I__1815 (
            .O(N__8404),
            .I(N__8396));
    Span12Mux_s5_h I__1814 (
            .O(N__8401),
            .I(N__8396));
    Odrv12 I__1813 (
            .O(N__8396),
            .I(CLK40_PLL_i_i));
    InMux I__1812 (
            .O(N__8393),
            .I(N__8383));
    InMux I__1811 (
            .O(N__8392),
            .I(N__8376));
    InMux I__1810 (
            .O(N__8391),
            .I(N__8376));
    InMux I__1809 (
            .O(N__8390),
            .I(N__8376));
    InMux I__1808 (
            .O(N__8389),
            .I(N__8365));
    InMux I__1807 (
            .O(N__8388),
            .I(N__8365));
    InMux I__1806 (
            .O(N__8387),
            .I(N__8365));
    InMux I__1805 (
            .O(N__8386),
            .I(N__8356));
    LocalMux I__1804 (
            .O(N__8383),
            .I(N__8353));
    LocalMux I__1803 (
            .O(N__8376),
            .I(N__8350));
    InMux I__1802 (
            .O(N__8375),
            .I(N__8345));
    InMux I__1801 (
            .O(N__8374),
            .I(N__8345));
    InMux I__1800 (
            .O(N__8373),
            .I(N__8342));
    InMux I__1799 (
            .O(N__8372),
            .I(N__8339));
    LocalMux I__1798 (
            .O(N__8365),
            .I(N__8336));
    InMux I__1797 (
            .O(N__8364),
            .I(N__8329));
    InMux I__1796 (
            .O(N__8363),
            .I(N__8329));
    InMux I__1795 (
            .O(N__8362),
            .I(N__8329));
    InMux I__1794 (
            .O(N__8361),
            .I(N__8326));
    InMux I__1793 (
            .O(N__8360),
            .I(N__8321));
    InMux I__1792 (
            .O(N__8359),
            .I(N__8321));
    LocalMux I__1791 (
            .O(N__8356),
            .I(N__8318));
    Span4Mux_v I__1790 (
            .O(N__8353),
            .I(N__8315));
    Span4Mux_v I__1789 (
            .O(N__8350),
            .I(N__8308));
    LocalMux I__1788 (
            .O(N__8345),
            .I(N__8308));
    LocalMux I__1787 (
            .O(N__8342),
            .I(N__8308));
    LocalMux I__1786 (
            .O(N__8339),
            .I(N__8305));
    Span4Mux_h I__1785 (
            .O(N__8336),
            .I(N__8296));
    LocalMux I__1784 (
            .O(N__8329),
            .I(N__8296));
    LocalMux I__1783 (
            .O(N__8326),
            .I(N__8296));
    LocalMux I__1782 (
            .O(N__8321),
            .I(N__8296));
    Sp12to4 I__1781 (
            .O(N__8318),
            .I(N__8292));
    Span4Mux_v I__1780 (
            .O(N__8315),
            .I(N__8287));
    Span4Mux_v I__1779 (
            .O(N__8308),
            .I(N__8287));
    Span4Mux_v I__1778 (
            .O(N__8305),
            .I(N__8282));
    Span4Mux_v I__1777 (
            .O(N__8296),
            .I(N__8282));
    InMux I__1776 (
            .O(N__8295),
            .I(N__8279));
    Span12Mux_v I__1775 (
            .O(N__8292),
            .I(N__8270));
    Sp12to4 I__1774 (
            .O(N__8287),
            .I(N__8270));
    Sp12to4 I__1773 (
            .O(N__8282),
            .I(N__8270));
    LocalMux I__1772 (
            .O(N__8279),
            .I(N__8270));
    Span12Mux_h I__1771 (
            .O(N__8270),
            .I(N__8267));
    Odrv12 I__1770 (
            .O(N__8267),
            .I(RESETn_c));
    IoInMux I__1769 (
            .O(N__8264),
            .I(N__8261));
    LocalMux I__1768 (
            .O(N__8261),
            .I(N__8258));
    Span12Mux_s1_v I__1767 (
            .O(N__8258),
            .I(N__8255));
    Odrv12 I__1766 (
            .O(N__8255),
            .I(RESETn_c_i));
    InMux I__1765 (
            .O(N__8252),
            .I(N__8245));
    InMux I__1764 (
            .O(N__8251),
            .I(N__8245));
    InMux I__1763 (
            .O(N__8250),
            .I(N__8242));
    LocalMux I__1762 (
            .O(N__8245),
            .I(N__8236));
    LocalMux I__1761 (
            .O(N__8242),
            .I(N__8236));
    CascadeMux I__1760 (
            .O(N__8241),
            .I(N__8233));
    Span4Mux_v I__1759 (
            .O(N__8236),
            .I(N__8229));
    InMux I__1758 (
            .O(N__8233),
            .I(N__8226));
    InMux I__1757 (
            .O(N__8232),
            .I(N__8223));
    Span4Mux_v I__1756 (
            .O(N__8229),
            .I(N__8216));
    LocalMux I__1755 (
            .O(N__8226),
            .I(N__8216));
    LocalMux I__1754 (
            .O(N__8223),
            .I(N__8216));
    Span4Mux_v I__1753 (
            .O(N__8216),
            .I(N__8212));
    InMux I__1752 (
            .O(N__8215),
            .I(N__8209));
    Span4Mux_v I__1751 (
            .O(N__8212),
            .I(N__8206));
    LocalMux I__1750 (
            .O(N__8209),
            .I(N__8203));
    Sp12to4 I__1749 (
            .O(N__8206),
            .I(N__8198));
    Span12Mux_v I__1748 (
            .O(N__8203),
            .I(N__8198));
    Span12Mux_h I__1747 (
            .O(N__8198),
            .I(N__8195));
    Odrv12 I__1746 (
            .O(N__8195),
            .I(CASLn_c));
    InMux I__1745 (
            .O(N__8192),
            .I(N__8184));
    InMux I__1744 (
            .O(N__8191),
            .I(N__8184));
    InMux I__1743 (
            .O(N__8190),
            .I(N__8181));
    InMux I__1742 (
            .O(N__8189),
            .I(N__8178));
    LocalMux I__1741 (
            .O(N__8184),
            .I(N__8173));
    LocalMux I__1740 (
            .O(N__8181),
            .I(N__8173));
    LocalMux I__1739 (
            .O(N__8178),
            .I(N__8168));
    Span4Mux_v I__1738 (
            .O(N__8173),
            .I(N__8165));
    InMux I__1737 (
            .O(N__8172),
            .I(N__8160));
    InMux I__1736 (
            .O(N__8171),
            .I(N__8160));
    Span4Mux_v I__1735 (
            .O(N__8168),
            .I(N__8157));
    Sp12to4 I__1734 (
            .O(N__8165),
            .I(N__8154));
    LocalMux I__1733 (
            .O(N__8160),
            .I(N__8151));
    Span4Mux_v I__1732 (
            .O(N__8157),
            .I(N__8148));
    Span12Mux_h I__1731 (
            .O(N__8154),
            .I(N__8145));
    Span12Mux_v I__1730 (
            .O(N__8151),
            .I(N__8142));
    Sp12to4 I__1729 (
            .O(N__8148),
            .I(N__8139));
    Span12Mux_v I__1728 (
            .O(N__8145),
            .I(N__8134));
    Span12Mux_h I__1727 (
            .O(N__8142),
            .I(N__8134));
    Span12Mux_h I__1726 (
            .O(N__8139),
            .I(N__8131));
    Odrv12 I__1725 (
            .O(N__8134),
            .I(CASUn_c));
    Odrv12 I__1724 (
            .O(N__8131),
            .I(CASUn_c));
    InMux I__1723 (
            .O(N__8126),
            .I(N__8121));
    InMux I__1722 (
            .O(N__8125),
            .I(N__8118));
    InMux I__1721 (
            .O(N__8124),
            .I(N__8115));
    LocalMux I__1720 (
            .O(N__8121),
            .I(N__8112));
    LocalMux I__1719 (
            .O(N__8118),
            .I(N__8109));
    LocalMux I__1718 (
            .O(N__8115),
            .I(N__8106));
    Span4Mux_h I__1717 (
            .O(N__8112),
            .I(N__8103));
    Span12Mux_h I__1716 (
            .O(N__8109),
            .I(N__8100));
    Span4Mux_v I__1715 (
            .O(N__8106),
            .I(N__8097));
    Span4Mux_v I__1714 (
            .O(N__8103),
            .I(N__8094));
    Span12Mux_v I__1713 (
            .O(N__8100),
            .I(N__8091));
    Span4Mux_h I__1712 (
            .O(N__8097),
            .I(N__8088));
    Span4Mux_v I__1711 (
            .O(N__8094),
            .I(N__8085));
    Odrv12 I__1710 (
            .O(N__8091),
            .I(REG_CYCLEm));
    Odrv4 I__1709 (
            .O(N__8088),
            .I(REG_CYCLEm));
    Odrv4 I__1708 (
            .O(N__8085),
            .I(REG_CYCLEm));
    IoInMux I__1707 (
            .O(N__8078),
            .I(N__8075));
    LocalMux I__1706 (
            .O(N__8075),
            .I(N__8072));
    Span4Mux_s1_v I__1705 (
            .O(N__8072),
            .I(N__8069));
    Span4Mux_h I__1704 (
            .O(N__8069),
            .I(N__8066));
    Sp12to4 I__1703 (
            .O(N__8066),
            .I(N__8063));
    Span12Mux_h I__1702 (
            .O(N__8063),
            .I(N__8060));
    Odrv12 I__1701 (
            .O(N__8060),
            .I(DRDENn_c));
    IoInMux I__1700 (
            .O(N__8057),
            .I(N__8054));
    LocalMux I__1699 (
            .O(N__8054),
            .I(N__8051));
    Span4Mux_s3_v I__1698 (
            .O(N__8051),
            .I(N__8048));
    Span4Mux_v I__1697 (
            .O(N__8048),
            .I(N__8045));
    Span4Mux_h I__1696 (
            .O(N__8045),
            .I(N__8042));
    Odrv4 I__1695 (
            .O(N__8042),
            .I(CRCSn_c));
    InMux I__1694 (
            .O(N__8039),
            .I(N__8036));
    LocalMux I__1693 (
            .O(N__8036),
            .I(N__8033));
    Span4Mux_v I__1692 (
            .O(N__8033),
            .I(N__8030));
    Span4Mux_h I__1691 (
            .O(N__8030),
            .I(N__8027));
    Odrv4 I__1690 (
            .O(N__8027),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    IoInMux I__1689 (
            .O(N__8024),
            .I(N__8021));
    LocalMux I__1688 (
            .O(N__8021),
            .I(N__8018));
    IoSpan4Mux I__1687 (
            .O(N__8018),
            .I(N__8015));
    Span4Mux_s1_h I__1686 (
            .O(N__8015),
            .I(N__8012));
    Sp12to4 I__1685 (
            .O(N__8012),
            .I(N__8009));
    Span12Mux_h I__1684 (
            .O(N__8009),
            .I(N__8006));
    Odrv12 I__1683 (
            .O(N__8006),
            .I(CMA_c_3));
    InMux I__1682 (
            .O(N__8003),
            .I(N__8000));
    LocalMux I__1681 (
            .O(N__8000),
            .I(N__7997));
    Span4Mux_v I__1680 (
            .O(N__7997),
            .I(N__7994));
    Span4Mux_v I__1679 (
            .O(N__7994),
            .I(N__7991));
    Sp12to4 I__1678 (
            .O(N__7991),
            .I(N__7988));
    Span12Mux_h I__1677 (
            .O(N__7988),
            .I(N__7985));
    Odrv12 I__1676 (
            .O(N__7985),
            .I(A_c_7));
    CascadeMux I__1675 (
            .O(N__7982),
            .I(\U712_CHIP_RAM.N_463_cascade_ ));
    InMux I__1674 (
            .O(N__7979),
            .I(N__7976));
    LocalMux I__1673 (
            .O(N__7976),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i ));
    InMux I__1672 (
            .O(N__7973),
            .I(N__7958));
    InMux I__1671 (
            .O(N__7972),
            .I(N__7958));
    InMux I__1670 (
            .O(N__7971),
            .I(N__7958));
    InMux I__1669 (
            .O(N__7970),
            .I(N__7955));
    InMux I__1668 (
            .O(N__7969),
            .I(N__7952));
    CascadeMux I__1667 (
            .O(N__7968),
            .I(N__7946));
    CascadeMux I__1666 (
            .O(N__7967),
            .I(N__7942));
    InMux I__1665 (
            .O(N__7966),
            .I(N__7937));
    InMux I__1664 (
            .O(N__7965),
            .I(N__7937));
    LocalMux I__1663 (
            .O(N__7958),
            .I(N__7934));
    LocalMux I__1662 (
            .O(N__7955),
            .I(N__7929));
    LocalMux I__1661 (
            .O(N__7952),
            .I(N__7929));
    InMux I__1660 (
            .O(N__7951),
            .I(N__7924));
    InMux I__1659 (
            .O(N__7950),
            .I(N__7924));
    InMux I__1658 (
            .O(N__7949),
            .I(N__7918));
    InMux I__1657 (
            .O(N__7946),
            .I(N__7915));
    InMux I__1656 (
            .O(N__7945),
            .I(N__7910));
    InMux I__1655 (
            .O(N__7942),
            .I(N__7910));
    LocalMux I__1654 (
            .O(N__7937),
            .I(N__7907));
    Span4Mux_h I__1653 (
            .O(N__7934),
            .I(N__7904));
    Span4Mux_v I__1652 (
            .O(N__7929),
            .I(N__7899));
    LocalMux I__1651 (
            .O(N__7924),
            .I(N__7899));
    InMux I__1650 (
            .O(N__7923),
            .I(N__7896));
    InMux I__1649 (
            .O(N__7922),
            .I(N__7893));
    InMux I__1648 (
            .O(N__7921),
            .I(N__7890));
    LocalMux I__1647 (
            .O(N__7918),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1646 (
            .O(N__7915),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1645 (
            .O(N__7910),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1644 (
            .O(N__7907),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1643 (
            .O(N__7904),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1642 (
            .O(N__7899),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1641 (
            .O(N__7896),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1640 (
            .O(N__7893),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1639 (
            .O(N__7890),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__1638 (
            .O(N__7871),
            .I(N__7864));
    InMux I__1637 (
            .O(N__7870),
            .I(N__7861));
    InMux I__1636 (
            .O(N__7869),
            .I(N__7858));
    InMux I__1635 (
            .O(N__7868),
            .I(N__7855));
    CascadeMux I__1634 (
            .O(N__7867),
            .I(N__7852));
    LocalMux I__1633 (
            .O(N__7864),
            .I(N__7841));
    LocalMux I__1632 (
            .O(N__7861),
            .I(N__7841));
    LocalMux I__1631 (
            .O(N__7858),
            .I(N__7836));
    LocalMux I__1630 (
            .O(N__7855),
            .I(N__7836));
    InMux I__1629 (
            .O(N__7852),
            .I(N__7833));
    InMux I__1628 (
            .O(N__7851),
            .I(N__7829));
    InMux I__1627 (
            .O(N__7850),
            .I(N__7826));
    InMux I__1626 (
            .O(N__7849),
            .I(N__7823));
    CascadeMux I__1625 (
            .O(N__7848),
            .I(N__7820));
    CascadeMux I__1624 (
            .O(N__7847),
            .I(N__7816));
    InMux I__1623 (
            .O(N__7846),
            .I(N__7805));
    Span4Mux_v I__1622 (
            .O(N__7841),
            .I(N__7802));
    Span4Mux_v I__1621 (
            .O(N__7836),
            .I(N__7797));
    LocalMux I__1620 (
            .O(N__7833),
            .I(N__7797));
    InMux I__1619 (
            .O(N__7832),
            .I(N__7794));
    LocalMux I__1618 (
            .O(N__7829),
            .I(N__7787));
    LocalMux I__1617 (
            .O(N__7826),
            .I(N__7787));
    LocalMux I__1616 (
            .O(N__7823),
            .I(N__7787));
    InMux I__1615 (
            .O(N__7820),
            .I(N__7778));
    InMux I__1614 (
            .O(N__7819),
            .I(N__7778));
    InMux I__1613 (
            .O(N__7816),
            .I(N__7778));
    InMux I__1612 (
            .O(N__7815),
            .I(N__7778));
    InMux I__1611 (
            .O(N__7814),
            .I(N__7775));
    InMux I__1610 (
            .O(N__7813),
            .I(N__7762));
    InMux I__1609 (
            .O(N__7812),
            .I(N__7762));
    InMux I__1608 (
            .O(N__7811),
            .I(N__7762));
    InMux I__1607 (
            .O(N__7810),
            .I(N__7762));
    InMux I__1606 (
            .O(N__7809),
            .I(N__7762));
    InMux I__1605 (
            .O(N__7808),
            .I(N__7762));
    LocalMux I__1604 (
            .O(N__7805),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1603 (
            .O(N__7802),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1602 (
            .O(N__7797),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1601 (
            .O(N__7794),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1600 (
            .O(N__7787),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1599 (
            .O(N__7778),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1598 (
            .O(N__7775),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1597 (
            .O(N__7762),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__1596 (
            .O(N__7745),
            .I(N__7742));
    LocalMux I__1595 (
            .O(N__7742),
            .I(N__7737));
    InMux I__1594 (
            .O(N__7741),
            .I(N__7734));
    InMux I__1593 (
            .O(N__7740),
            .I(N__7731));
    Span4Mux_v I__1592 (
            .O(N__7737),
            .I(N__7726));
    LocalMux I__1591 (
            .O(N__7734),
            .I(N__7726));
    LocalMux I__1590 (
            .O(N__7731),
            .I(N__7723));
    Span4Mux_h I__1589 (
            .O(N__7726),
            .I(N__7720));
    Odrv12 I__1588 (
            .O(N__7723),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRTZ0Z_2 ));
    Odrv4 I__1587 (
            .O(N__7720),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRTZ0Z_2 ));
    InMux I__1586 (
            .O(N__7715),
            .I(N__7712));
    LocalMux I__1585 (
            .O(N__7712),
            .I(N__7709));
    Odrv4 I__1584 (
            .O(N__7709),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__1583 (
            .O(N__7706),
            .I(N__7703));
    LocalMux I__1582 (
            .O(N__7703),
            .I(N__7700));
    Odrv12 I__1581 (
            .O(N__7700),
            .I(\U712_CHIP_RAM.un3_DMA_CYCLE_START ));
    InMux I__1580 (
            .O(N__7697),
            .I(N__7691));
    InMux I__1579 (
            .O(N__7696),
            .I(N__7691));
    LocalMux I__1578 (
            .O(N__7691),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__1577 (
            .O(N__7688),
            .I(N__7685));
    LocalMux I__1576 (
            .O(N__7685),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__1575 (
            .O(N__7682),
            .I(N__7679));
    LocalMux I__1574 (
            .O(N__7679),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ));
    IoInMux I__1573 (
            .O(N__7676),
            .I(N__7673));
    LocalMux I__1572 (
            .O(N__7673),
            .I(N__7670));
    Span4Mux_s1_v I__1571 (
            .O(N__7670),
            .I(N__7667));
    Span4Mux_v I__1570 (
            .O(N__7667),
            .I(N__7664));
    Span4Mux_v I__1569 (
            .O(N__7664),
            .I(N__7661));
    Odrv4 I__1568 (
            .O(N__7661),
            .I(CMA_c_2));
    InMux I__1567 (
            .O(N__7658),
            .I(N__7655));
    LocalMux I__1566 (
            .O(N__7655),
            .I(N__7652));
    Span4Mux_h I__1565 (
            .O(N__7652),
            .I(N__7649));
    Span4Mux_v I__1564 (
            .O(N__7649),
            .I(N__7646));
    Odrv4 I__1563 (
            .O(N__7646),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ));
    CascadeMux I__1562 (
            .O(N__7643),
            .I(\U712_CHIP_RAM.CMA_5_0_8_cascade_ ));
    InMux I__1561 (
            .O(N__7640),
            .I(N__7634));
    InMux I__1560 (
            .O(N__7639),
            .I(N__7634));
    LocalMux I__1559 (
            .O(N__7634),
            .I(N__7631));
    Span4Mux_v I__1558 (
            .O(N__7631),
            .I(N__7628));
    Span4Mux_v I__1557 (
            .O(N__7628),
            .I(N__7625));
    Sp12to4 I__1556 (
            .O(N__7625),
            .I(N__7622));
    Span12Mux_h I__1555 (
            .O(N__7622),
            .I(N__7619));
    Odrv12 I__1554 (
            .O(N__7619),
            .I(A_c_14));
    CascadeMux I__1553 (
            .O(N__7616),
            .I(N__7613));
    InMux I__1552 (
            .O(N__7613),
            .I(N__7606));
    InMux I__1551 (
            .O(N__7612),
            .I(N__7596));
    InMux I__1550 (
            .O(N__7611),
            .I(N__7596));
    InMux I__1549 (
            .O(N__7610),
            .I(N__7596));
    InMux I__1548 (
            .O(N__7609),
            .I(N__7596));
    LocalMux I__1547 (
            .O(N__7606),
            .I(N__7593));
    InMux I__1546 (
            .O(N__7605),
            .I(N__7590));
    LocalMux I__1545 (
            .O(N__7596),
            .I(N__7585));
    Span4Mux_v I__1544 (
            .O(N__7593),
            .I(N__7580));
    LocalMux I__1543 (
            .O(N__7590),
            .I(N__7580));
    InMux I__1542 (
            .O(N__7589),
            .I(N__7575));
    InMux I__1541 (
            .O(N__7588),
            .I(N__7575));
    Odrv12 I__1540 (
            .O(N__7585),
            .I(DMA_CYCLEm));
    Odrv4 I__1539 (
            .O(N__7580),
            .I(DMA_CYCLEm));
    LocalMux I__1538 (
            .O(N__7575),
            .I(DMA_CYCLEm));
    InMux I__1537 (
            .O(N__7568),
            .I(N__7563));
    CascadeMux I__1536 (
            .O(N__7567),
            .I(N__7559));
    CascadeMux I__1535 (
            .O(N__7566),
            .I(N__7556));
    LocalMux I__1534 (
            .O(N__7563),
            .I(N__7553));
    InMux I__1533 (
            .O(N__7562),
            .I(N__7550));
    InMux I__1532 (
            .O(N__7559),
            .I(N__7547));
    InMux I__1531 (
            .O(N__7556),
            .I(N__7542));
    Span4Mux_v I__1530 (
            .O(N__7553),
            .I(N__7537));
    LocalMux I__1529 (
            .O(N__7550),
            .I(N__7537));
    LocalMux I__1528 (
            .O(N__7547),
            .I(N__7534));
    InMux I__1527 (
            .O(N__7546),
            .I(N__7531));
    InMux I__1526 (
            .O(N__7545),
            .I(N__7528));
    LocalMux I__1525 (
            .O(N__7542),
            .I(N__7525));
    Span4Mux_v I__1524 (
            .O(N__7537),
            .I(N__7522));
    Span4Mux_h I__1523 (
            .O(N__7534),
            .I(N__7518));
    LocalMux I__1522 (
            .O(N__7531),
            .I(N__7513));
    LocalMux I__1521 (
            .O(N__7528),
            .I(N__7513));
    Span4Mux_h I__1520 (
            .O(N__7525),
            .I(N__7507));
    Span4Mux_h I__1519 (
            .O(N__7522),
            .I(N__7504));
    InMux I__1518 (
            .O(N__7521),
            .I(N__7501));
    Span4Mux_h I__1517 (
            .O(N__7518),
            .I(N__7496));
    Span4Mux_h I__1516 (
            .O(N__7513),
            .I(N__7496));
    InMux I__1515 (
            .O(N__7512),
            .I(N__7491));
    InMux I__1514 (
            .O(N__7511),
            .I(N__7491));
    InMux I__1513 (
            .O(N__7510),
            .I(N__7488));
    Odrv4 I__1512 (
            .O(N__7507),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1511 (
            .O(N__7504),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1510 (
            .O(N__7501),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1509 (
            .O(N__7496),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1508 (
            .O(N__7491),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1507 (
            .O(N__7488),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    InMux I__1506 (
            .O(N__7475),
            .I(N__7472));
    LocalMux I__1505 (
            .O(N__7472),
            .I(N__7469));
    Span4Mux_v I__1504 (
            .O(N__7469),
            .I(N__7465));
    InMux I__1503 (
            .O(N__7468),
            .I(N__7462));
    Odrv4 I__1502 (
            .O(N__7465),
            .I(\U712_CHIP_RAM.N_201_i_i_a2_3_1 ));
    LocalMux I__1501 (
            .O(N__7462),
            .I(\U712_CHIP_RAM.N_201_i_i_a2_3_1 ));
    SRMux I__1500 (
            .O(N__7457),
            .I(N__7454));
    LocalMux I__1499 (
            .O(N__7454),
            .I(N__7451));
    Span4Mux_h I__1498 (
            .O(N__7451),
            .I(N__7448));
    Odrv4 I__1497 (
            .O(N__7448),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    CascadeMux I__1496 (
            .O(N__7445),
            .I(N__7440));
    InMux I__1495 (
            .O(N__7444),
            .I(N__7429));
    CascadeMux I__1494 (
            .O(N__7443),
            .I(N__7423));
    InMux I__1493 (
            .O(N__7440),
            .I(N__7420));
    InMux I__1492 (
            .O(N__7439),
            .I(N__7417));
    InMux I__1491 (
            .O(N__7438),
            .I(N__7410));
    InMux I__1490 (
            .O(N__7437),
            .I(N__7403));
    InMux I__1489 (
            .O(N__7436),
            .I(N__7403));
    InMux I__1488 (
            .O(N__7435),
            .I(N__7403));
    InMux I__1487 (
            .O(N__7434),
            .I(N__7396));
    InMux I__1486 (
            .O(N__7433),
            .I(N__7396));
    InMux I__1485 (
            .O(N__7432),
            .I(N__7396));
    LocalMux I__1484 (
            .O(N__7429),
            .I(N__7392));
    InMux I__1483 (
            .O(N__7428),
            .I(N__7387));
    InMux I__1482 (
            .O(N__7427),
            .I(N__7387));
    InMux I__1481 (
            .O(N__7426),
            .I(N__7382));
    InMux I__1480 (
            .O(N__7423),
            .I(N__7375));
    LocalMux I__1479 (
            .O(N__7420),
            .I(N__7372));
    LocalMux I__1478 (
            .O(N__7417),
            .I(N__7369));
    InMux I__1477 (
            .O(N__7416),
            .I(N__7360));
    InMux I__1476 (
            .O(N__7415),
            .I(N__7360));
    InMux I__1475 (
            .O(N__7414),
            .I(N__7360));
    InMux I__1474 (
            .O(N__7413),
            .I(N__7360));
    LocalMux I__1473 (
            .O(N__7410),
            .I(N__7353));
    LocalMux I__1472 (
            .O(N__7403),
            .I(N__7353));
    LocalMux I__1471 (
            .O(N__7396),
            .I(N__7353));
    InMux I__1470 (
            .O(N__7395),
            .I(N__7350));
    Span4Mux_v I__1469 (
            .O(N__7392),
            .I(N__7345));
    LocalMux I__1468 (
            .O(N__7387),
            .I(N__7345));
    InMux I__1467 (
            .O(N__7386),
            .I(N__7340));
    InMux I__1466 (
            .O(N__7385),
            .I(N__7340));
    LocalMux I__1465 (
            .O(N__7382),
            .I(N__7337));
    InMux I__1464 (
            .O(N__7381),
            .I(N__7334));
    InMux I__1463 (
            .O(N__7380),
            .I(N__7327));
    InMux I__1462 (
            .O(N__7379),
            .I(N__7327));
    InMux I__1461 (
            .O(N__7378),
            .I(N__7327));
    LocalMux I__1460 (
            .O(N__7375),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv12 I__1459 (
            .O(N__7372),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1458 (
            .O(N__7369),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1457 (
            .O(N__7360),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1456 (
            .O(N__7353),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1455 (
            .O(N__7350),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1454 (
            .O(N__7345),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1453 (
            .O(N__7340),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1452 (
            .O(N__7337),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1451 (
            .O(N__7334),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1450 (
            .O(N__7327),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__1449 (
            .O(N__7304),
            .I(N__7298));
    InMux I__1448 (
            .O(N__7303),
            .I(N__7298));
    LocalMux I__1447 (
            .O(N__7298),
            .I(N__7295));
    Span4Mux_v I__1446 (
            .O(N__7295),
            .I(N__7291));
    InMux I__1445 (
            .O(N__7294),
            .I(N__7288));
    Span4Mux_v I__1444 (
            .O(N__7291),
            .I(N__7279));
    LocalMux I__1443 (
            .O(N__7288),
            .I(N__7279));
    InMux I__1442 (
            .O(N__7287),
            .I(N__7276));
    InMux I__1441 (
            .O(N__7286),
            .I(N__7273));
    InMux I__1440 (
            .O(N__7285),
            .I(N__7270));
    InMux I__1439 (
            .O(N__7284),
            .I(N__7265));
    Span4Mux_v I__1438 (
            .O(N__7279),
            .I(N__7256));
    LocalMux I__1437 (
            .O(N__7276),
            .I(N__7256));
    LocalMux I__1436 (
            .O(N__7273),
            .I(N__7256));
    LocalMux I__1435 (
            .O(N__7270),
            .I(N__7256));
    InMux I__1434 (
            .O(N__7269),
            .I(N__7251));
    InMux I__1433 (
            .O(N__7268),
            .I(N__7251));
    LocalMux I__1432 (
            .O(N__7265),
            .I(N__7248));
    Span4Mux_v I__1431 (
            .O(N__7256),
            .I(N__7242));
    LocalMux I__1430 (
            .O(N__7251),
            .I(N__7239));
    Span4Mux_v I__1429 (
            .O(N__7248),
            .I(N__7236));
    InMux I__1428 (
            .O(N__7247),
            .I(N__7229));
    InMux I__1427 (
            .O(N__7246),
            .I(N__7229));
    InMux I__1426 (
            .O(N__7245),
            .I(N__7229));
    Odrv4 I__1425 (
            .O(N__7242),
            .I(WRITE_CYCLEm));
    Odrv4 I__1424 (
            .O(N__7239),
            .I(WRITE_CYCLEm));
    Odrv4 I__1423 (
            .O(N__7236),
            .I(WRITE_CYCLEm));
    LocalMux I__1422 (
            .O(N__7229),
            .I(WRITE_CYCLEm));
    InMux I__1421 (
            .O(N__7220),
            .I(N__7214));
    InMux I__1420 (
            .O(N__7219),
            .I(N__7211));
    InMux I__1419 (
            .O(N__7218),
            .I(N__7206));
    InMux I__1418 (
            .O(N__7217),
            .I(N__7203));
    LocalMux I__1417 (
            .O(N__7214),
            .I(N__7199));
    LocalMux I__1416 (
            .O(N__7211),
            .I(N__7196));
    InMux I__1415 (
            .O(N__7210),
            .I(N__7188));
    InMux I__1414 (
            .O(N__7209),
            .I(N__7188));
    LocalMux I__1413 (
            .O(N__7206),
            .I(N__7183));
    LocalMux I__1412 (
            .O(N__7203),
            .I(N__7183));
    InMux I__1411 (
            .O(N__7202),
            .I(N__7180));
    Span4Mux_h I__1410 (
            .O(N__7199),
            .I(N__7175));
    Span4Mux_h I__1409 (
            .O(N__7196),
            .I(N__7175));
    InMux I__1408 (
            .O(N__7195),
            .I(N__7168));
    InMux I__1407 (
            .O(N__7194),
            .I(N__7168));
    InMux I__1406 (
            .O(N__7193),
            .I(N__7168));
    LocalMux I__1405 (
            .O(N__7188),
            .I(N__7161));
    Span4Mux_v I__1404 (
            .O(N__7183),
            .I(N__7161));
    LocalMux I__1403 (
            .O(N__7180),
            .I(N__7161));
    Odrv4 I__1402 (
            .O(N__7175),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1401 (
            .O(N__7168),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1400 (
            .O(N__7161),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    CascadeMux I__1399 (
            .O(N__7154),
            .I(\U712_CHIP_RAM.N_306_cascade_ ));
    InMux I__1398 (
            .O(N__7151),
            .I(N__7147));
    CascadeMux I__1397 (
            .O(N__7150),
            .I(N__7139));
    LocalMux I__1396 (
            .O(N__7147),
            .I(N__7135));
    InMux I__1395 (
            .O(N__7146),
            .I(N__7132));
    InMux I__1394 (
            .O(N__7145),
            .I(N__7127));
    InMux I__1393 (
            .O(N__7144),
            .I(N__7127));
    InMux I__1392 (
            .O(N__7143),
            .I(N__7122));
    CascadeMux I__1391 (
            .O(N__7142),
            .I(N__7118));
    InMux I__1390 (
            .O(N__7139),
            .I(N__7115));
    CascadeMux I__1389 (
            .O(N__7138),
            .I(N__7109));
    Span4Mux_h I__1388 (
            .O(N__7135),
            .I(N__7102));
    LocalMux I__1387 (
            .O(N__7132),
            .I(N__7102));
    LocalMux I__1386 (
            .O(N__7127),
            .I(N__7102));
    InMux I__1385 (
            .O(N__7126),
            .I(N__7099));
    InMux I__1384 (
            .O(N__7125),
            .I(N__7094));
    LocalMux I__1383 (
            .O(N__7122),
            .I(N__7091));
    InMux I__1382 (
            .O(N__7121),
            .I(N__7086));
    InMux I__1381 (
            .O(N__7118),
            .I(N__7086));
    LocalMux I__1380 (
            .O(N__7115),
            .I(N__7083));
    InMux I__1379 (
            .O(N__7114),
            .I(N__7080));
    CascadeMux I__1378 (
            .O(N__7113),
            .I(N__7076));
    CascadeMux I__1377 (
            .O(N__7112),
            .I(N__7073));
    InMux I__1376 (
            .O(N__7109),
            .I(N__7066));
    Span4Mux_v I__1375 (
            .O(N__7102),
            .I(N__7063));
    LocalMux I__1374 (
            .O(N__7099),
            .I(N__7060));
    InMux I__1373 (
            .O(N__7098),
            .I(N__7055));
    InMux I__1372 (
            .O(N__7097),
            .I(N__7055));
    LocalMux I__1371 (
            .O(N__7094),
            .I(N__7044));
    Span4Mux_v I__1370 (
            .O(N__7091),
            .I(N__7044));
    LocalMux I__1369 (
            .O(N__7086),
            .I(N__7044));
    Span4Mux_v I__1368 (
            .O(N__7083),
            .I(N__7044));
    LocalMux I__1367 (
            .O(N__7080),
            .I(N__7044));
    InMux I__1366 (
            .O(N__7079),
            .I(N__7037));
    InMux I__1365 (
            .O(N__7076),
            .I(N__7037));
    InMux I__1364 (
            .O(N__7073),
            .I(N__7037));
    InMux I__1363 (
            .O(N__7072),
            .I(N__7034));
    InMux I__1362 (
            .O(N__7071),
            .I(N__7031));
    InMux I__1361 (
            .O(N__7070),
            .I(N__7026));
    InMux I__1360 (
            .O(N__7069),
            .I(N__7026));
    LocalMux I__1359 (
            .O(N__7066),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1358 (
            .O(N__7063),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv12 I__1357 (
            .O(N__7060),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1356 (
            .O(N__7055),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1355 (
            .O(N__7044),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1354 (
            .O(N__7037),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1353 (
            .O(N__7034),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1352 (
            .O(N__7031),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1351 (
            .O(N__7026),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__1350 (
            .O(N__7007),
            .I(N__7004));
    LocalMux I__1349 (
            .O(N__7004),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_i_0 ));
    InMux I__1348 (
            .O(N__7001),
            .I(N__6997));
    InMux I__1347 (
            .O(N__7000),
            .I(N__6994));
    LocalMux I__1346 (
            .O(N__6997),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    LocalMux I__1345 (
            .O(N__6994),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    InMux I__1344 (
            .O(N__6989),
            .I(N__6985));
    InMux I__1343 (
            .O(N__6988),
            .I(N__6982));
    LocalMux I__1342 (
            .O(N__6985),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__1341 (
            .O(N__6982),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    CascadeMux I__1340 (
            .O(N__6977),
            .I(N__6973));
    InMux I__1339 (
            .O(N__6976),
            .I(N__6970));
    InMux I__1338 (
            .O(N__6973),
            .I(N__6967));
    LocalMux I__1337 (
            .O(N__6970),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    LocalMux I__1336 (
            .O(N__6967),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    InMux I__1335 (
            .O(N__6962),
            .I(N__6958));
    InMux I__1334 (
            .O(N__6961),
            .I(N__6955));
    LocalMux I__1333 (
            .O(N__6958),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    LocalMux I__1332 (
            .O(N__6955),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__1331 (
            .O(N__6950),
            .I(N__6946));
    InMux I__1330 (
            .O(N__6949),
            .I(N__6943));
    LocalMux I__1329 (
            .O(N__6946),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__1328 (
            .O(N__6943),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__1327 (
            .O(N__6938),
            .I(N__6934));
    InMux I__1326 (
            .O(N__6937),
            .I(N__6931));
    LocalMux I__1325 (
            .O(N__6934),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__1324 (
            .O(N__6931),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__1323 (
            .O(N__6926),
            .I(N__6922));
    InMux I__1322 (
            .O(N__6925),
            .I(N__6919));
    LocalMux I__1321 (
            .O(N__6922),
            .I(N__6916));
    LocalMux I__1320 (
            .O(N__6919),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    Odrv4 I__1319 (
            .O(N__6916),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__1318 (
            .O(N__6911),
            .I(N__6908));
    LocalMux I__1317 (
            .O(N__6908),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ));
    CascadeMux I__1316 (
            .O(N__6905),
            .I(N__6902));
    InMux I__1315 (
            .O(N__6902),
            .I(N__6898));
    InMux I__1314 (
            .O(N__6901),
            .I(N__6895));
    LocalMux I__1313 (
            .O(N__6898),
            .I(N__6892));
    LocalMux I__1312 (
            .O(N__6895),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    Odrv12 I__1311 (
            .O(N__6892),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__1310 (
            .O(N__6887),
            .I(N__6884));
    LocalMux I__1309 (
            .O(N__6884),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ));
    InMux I__1308 (
            .O(N__6881),
            .I(N__6877));
    InMux I__1307 (
            .O(N__6880),
            .I(N__6874));
    LocalMux I__1306 (
            .O(N__6877),
            .I(N__6871));
    LocalMux I__1305 (
            .O(N__6874),
            .I(N__6866));
    Span4Mux_h I__1304 (
            .O(N__6871),
            .I(N__6863));
    InMux I__1303 (
            .O(N__6870),
            .I(N__6860));
    InMux I__1302 (
            .O(N__6869),
            .I(N__6857));
    Odrv4 I__1301 (
            .O(N__6866),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    Odrv4 I__1300 (
            .O(N__6863),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__1299 (
            .O(N__6860),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__1298 (
            .O(N__6857),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    InMux I__1297 (
            .O(N__6848),
            .I(N__6835));
    InMux I__1296 (
            .O(N__6847),
            .I(N__6835));
    InMux I__1295 (
            .O(N__6846),
            .I(N__6835));
    InMux I__1294 (
            .O(N__6845),
            .I(N__6828));
    InMux I__1293 (
            .O(N__6844),
            .I(N__6828));
    InMux I__1292 (
            .O(N__6843),
            .I(N__6828));
    InMux I__1291 (
            .O(N__6842),
            .I(N__6825));
    LocalMux I__1290 (
            .O(N__6835),
            .I(N__6820));
    LocalMux I__1289 (
            .O(N__6828),
            .I(N__6820));
    LocalMux I__1288 (
            .O(N__6825),
            .I(\U712_CHIP_RAM.N_62 ));
    Odrv4 I__1287 (
            .O(N__6820),
            .I(\U712_CHIP_RAM.N_62 ));
    InMux I__1286 (
            .O(N__6815),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    CascadeMux I__1285 (
            .O(N__6812),
            .I(N__6808));
    InMux I__1284 (
            .O(N__6811),
            .I(N__6805));
    InMux I__1283 (
            .O(N__6808),
            .I(N__6802));
    LocalMux I__1282 (
            .O(N__6805),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__1281 (
            .O(N__6802),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    CEMux I__1280 (
            .O(N__6797),
            .I(N__6793));
    CEMux I__1279 (
            .O(N__6796),
            .I(N__6790));
    LocalMux I__1278 (
            .O(N__6793),
            .I(N__6787));
    LocalMux I__1277 (
            .O(N__6790),
            .I(N__6784));
    Odrv4 I__1276 (
            .O(N__6787),
            .I(\U712_CHIP_RAM.N_434_i ));
    Odrv4 I__1275 (
            .O(N__6784),
            .I(\U712_CHIP_RAM.N_434_i ));
    InMux I__1274 (
            .O(N__6779),
            .I(bfn_11_7_0_));
    InMux I__1273 (
            .O(N__6776),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__1272 (
            .O(N__6773),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__1271 (
            .O(N__6770),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__1270 (
            .O(N__6767),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__1269 (
            .O(N__6764),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__1268 (
            .O(N__6761),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__1267 (
            .O(N__6758),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    CascadeMux I__1266 (
            .O(N__6755),
            .I(N__6751));
    CascadeMux I__1265 (
            .O(N__6754),
            .I(N__6748));
    InMux I__1264 (
            .O(N__6751),
            .I(N__6744));
    InMux I__1263 (
            .O(N__6748),
            .I(N__6741));
    InMux I__1262 (
            .O(N__6747),
            .I(N__6738));
    LocalMux I__1261 (
            .O(N__6744),
            .I(N__6735));
    LocalMux I__1260 (
            .O(N__6741),
            .I(N__6726));
    LocalMux I__1259 (
            .O(N__6738),
            .I(N__6723));
    Glb2LocalMux I__1258 (
            .O(N__6735),
            .I(N__6704));
    ClkMux I__1257 (
            .O(N__6734),
            .I(N__6704));
    ClkMux I__1256 (
            .O(N__6733),
            .I(N__6704));
    ClkMux I__1255 (
            .O(N__6732),
            .I(N__6704));
    ClkMux I__1254 (
            .O(N__6731),
            .I(N__6704));
    ClkMux I__1253 (
            .O(N__6730),
            .I(N__6704));
    ClkMux I__1252 (
            .O(N__6729),
            .I(N__6704));
    Glb2LocalMux I__1251 (
            .O(N__6726),
            .I(N__6704));
    Glb2LocalMux I__1250 (
            .O(N__6723),
            .I(N__6704));
    GlobalMux I__1249 (
            .O(N__6704),
            .I(N__6701));
    gio2CtrlBuf I__1248 (
            .O(N__6701),
            .I(C1_c_g));
    CascadeMux I__1247 (
            .O(N__6698),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ));
    CascadeMux I__1246 (
            .O(N__6695),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_ ));
    IoInMux I__1245 (
            .O(N__6692),
            .I(N__6689));
    LocalMux I__1244 (
            .O(N__6689),
            .I(N__6686));
    IoSpan4Mux I__1243 (
            .O(N__6686),
            .I(N__6683));
    Span4Mux_s3_h I__1242 (
            .O(N__6683),
            .I(N__6680));
    Sp12to4 I__1241 (
            .O(N__6680),
            .I(N__6677));
    Span12Mux_h I__1240 (
            .O(N__6677),
            .I(N__6674));
    Odrv12 I__1239 (
            .O(N__6674),
            .I(CMA_c_6));
    InMux I__1238 (
            .O(N__6671),
            .I(N__6668));
    LocalMux I__1237 (
            .O(N__6668),
            .I(N__6665));
    Span4Mux_h I__1236 (
            .O(N__6665),
            .I(N__6662));
    Odrv4 I__1235 (
            .O(N__6662),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_1 ));
    InMux I__1234 (
            .O(N__6659),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__1233 (
            .O(N__6656),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    InMux I__1232 (
            .O(N__6653),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__1231 (
            .O(N__6650),
            .I(N__6646));
    InMux I__1230 (
            .O(N__6649),
            .I(N__6643));
    LocalMux I__1229 (
            .O(N__6646),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1228 (
            .O(N__6643),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__1227 (
            .O(N__6638),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__1226 (
            .O(N__6635),
            .I(N__6631));
    InMux I__1225 (
            .O(N__6634),
            .I(N__6628));
    LocalMux I__1224 (
            .O(N__6631),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__1223 (
            .O(N__6628),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    InMux I__1222 (
            .O(N__6623),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__1221 (
            .O(N__6620),
            .I(N__6616));
    InMux I__1220 (
            .O(N__6619),
            .I(N__6613));
    LocalMux I__1219 (
            .O(N__6616),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__1218 (
            .O(N__6613),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__1217 (
            .O(N__6608),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__1216 (
            .O(N__6605),
            .I(N__6602));
    LocalMux I__1215 (
            .O(N__6602),
            .I(N__6599));
    Odrv12 I__1214 (
            .O(N__6599),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2Z0Z_0 ));
    InMux I__1213 (
            .O(N__6596),
            .I(N__6593));
    LocalMux I__1212 (
            .O(N__6593),
            .I(\U712_BYTE_ENABLE.N_431 ));
    CascadeMux I__1211 (
            .O(N__6590),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2Z0Z_0_cascade_ ));
    IoInMux I__1210 (
            .O(N__6587),
            .I(N__6584));
    LocalMux I__1209 (
            .O(N__6584),
            .I(N__6581));
    Span12Mux_s3_v I__1208 (
            .O(N__6581),
            .I(N__6578));
    Span12Mux_v I__1207 (
            .O(N__6578),
            .I(N__6575));
    Odrv12 I__1206 (
            .O(N__6575),
            .I(N_45_i));
    InMux I__1205 (
            .O(N__6572),
            .I(N__6566));
    InMux I__1204 (
            .O(N__6571),
            .I(N__6566));
    LocalMux I__1203 (
            .O(N__6566),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2Z0Z_0 ));
    InMux I__1202 (
            .O(N__6563),
            .I(N__6559));
    InMux I__1201 (
            .O(N__6562),
            .I(N__6556));
    LocalMux I__1200 (
            .O(N__6559),
            .I(N__6551));
    LocalMux I__1199 (
            .O(N__6556),
            .I(N__6548));
    InMux I__1198 (
            .O(N__6555),
            .I(N__6545));
    InMux I__1197 (
            .O(N__6554),
            .I(N__6542));
    Span4Mux_v I__1196 (
            .O(N__6551),
            .I(N__6539));
    Span4Mux_v I__1195 (
            .O(N__6548),
            .I(N__6536));
    LocalMux I__1194 (
            .O(N__6545),
            .I(N__6533));
    LocalMux I__1193 (
            .O(N__6542),
            .I(N__6530));
    Sp12to4 I__1192 (
            .O(N__6539),
            .I(N__6525));
    Sp12to4 I__1191 (
            .O(N__6536),
            .I(N__6525));
    Span4Mux_v I__1190 (
            .O(N__6533),
            .I(N__6522));
    Span12Mux_h I__1189 (
            .O(N__6530),
            .I(N__6519));
    Span12Mux_h I__1188 (
            .O(N__6525),
            .I(N__6516));
    Sp12to4 I__1187 (
            .O(N__6522),
            .I(N__6513));
    Span12Mux_v I__1186 (
            .O(N__6519),
            .I(N__6510));
    Span12Mux_v I__1185 (
            .O(N__6516),
            .I(N__6505));
    Span12Mux_h I__1184 (
            .O(N__6513),
            .I(N__6505));
    Odrv12 I__1183 (
            .O(N__6510),
            .I(RnW_c));
    Odrv12 I__1182 (
            .O(N__6505),
            .I(RnW_c));
    IoInMux I__1181 (
            .O(N__6500),
            .I(N__6497));
    LocalMux I__1180 (
            .O(N__6497),
            .I(N__6494));
    IoSpan4Mux I__1179 (
            .O(N__6494),
            .I(N__6491));
    Span4Mux_s1_h I__1178 (
            .O(N__6491),
            .I(N__6488));
    Span4Mux_v I__1177 (
            .O(N__6488),
            .I(N__6485));
    Sp12to4 I__1176 (
            .O(N__6485),
            .I(N__6482));
    Span12Mux_s10_h I__1175 (
            .O(N__6482),
            .I(N__6479));
    Odrv12 I__1174 (
            .O(N__6479),
            .I(N_344));
    IoInMux I__1173 (
            .O(N__6476),
            .I(N__6473));
    LocalMux I__1172 (
            .O(N__6473),
            .I(N__6470));
    Span12Mux_s8_v I__1171 (
            .O(N__6470),
            .I(N__6467));
    Odrv12 I__1170 (
            .O(N__6467),
            .I(DMA_LATCH_EN_c));
    InMux I__1169 (
            .O(N__6464),
            .I(N__6461));
    LocalMux I__1168 (
            .O(N__6461),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ));
    InMux I__1167 (
            .O(N__6458),
            .I(N__6455));
    LocalMux I__1166 (
            .O(N__6455),
            .I(N__6452));
    Odrv4 I__1165 (
            .O(N__6452),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    CascadeMux I__1164 (
            .O(N__6449),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_ ));
    IoInMux I__1163 (
            .O(N__6446),
            .I(N__6443));
    LocalMux I__1162 (
            .O(N__6443),
            .I(N__6440));
    Span4Mux_s1_h I__1161 (
            .O(N__6440),
            .I(N__6437));
    Sp12to4 I__1160 (
            .O(N__6437),
            .I(N__6434));
    Span12Mux_s10_v I__1159 (
            .O(N__6434),
            .I(N__6431));
    Span12Mux_h I__1158 (
            .O(N__6431),
            .I(N__6428));
    Odrv12 I__1157 (
            .O(N__6428),
            .I(CMA_c_7));
    InMux I__1156 (
            .O(N__6425),
            .I(N__6422));
    LocalMux I__1155 (
            .O(N__6422),
            .I(N__6419));
    Span4Mux_v I__1154 (
            .O(N__6419),
            .I(N__6416));
    Span4Mux_v I__1153 (
            .O(N__6416),
            .I(N__6413));
    Sp12to4 I__1152 (
            .O(N__6413),
            .I(N__6410));
    Span12Mux_h I__1151 (
            .O(N__6410),
            .I(N__6407));
    Odrv12 I__1150 (
            .O(N__6407),
            .I(A_c_8));
    InMux I__1149 (
            .O(N__6404),
            .I(N__6401));
    LocalMux I__1148 (
            .O(N__6401),
            .I(N__6398));
    Sp12to4 I__1147 (
            .O(N__6398),
            .I(N__6395));
    Span12Mux_v I__1146 (
            .O(N__6395),
            .I(N__6392));
    Span12Mux_h I__1145 (
            .O(N__6392),
            .I(N__6389));
    Odrv12 I__1144 (
            .O(N__6389),
            .I(A_c_15));
    CascadeMux I__1143 (
            .O(N__6386),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNO_6Z0Z_1_cascade_ ));
    InMux I__1142 (
            .O(N__6383),
            .I(N__6380));
    LocalMux I__1141 (
            .O(N__6380),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1 ));
    InMux I__1140 (
            .O(N__6377),
            .I(N__6371));
    CascadeMux I__1139 (
            .O(N__6376),
            .I(N__6368));
    InMux I__1138 (
            .O(N__6375),
            .I(N__6365));
    InMux I__1137 (
            .O(N__6374),
            .I(N__6361));
    LocalMux I__1136 (
            .O(N__6371),
            .I(N__6358));
    InMux I__1135 (
            .O(N__6368),
            .I(N__6351));
    LocalMux I__1134 (
            .O(N__6365),
            .I(N__6348));
    InMux I__1133 (
            .O(N__6364),
            .I(N__6345));
    LocalMux I__1132 (
            .O(N__6361),
            .I(N__6340));
    Span4Mux_h I__1131 (
            .O(N__6358),
            .I(N__6340));
    InMux I__1130 (
            .O(N__6357),
            .I(N__6337));
    InMux I__1129 (
            .O(N__6356),
            .I(N__6330));
    InMux I__1128 (
            .O(N__6355),
            .I(N__6330));
    InMux I__1127 (
            .O(N__6354),
            .I(N__6330));
    LocalMux I__1126 (
            .O(N__6351),
            .I(\U712_CHIP_RAM.N_287 ));
    Odrv4 I__1125 (
            .O(N__6348),
            .I(\U712_CHIP_RAM.N_287 ));
    LocalMux I__1124 (
            .O(N__6345),
            .I(\U712_CHIP_RAM.N_287 ));
    Odrv4 I__1123 (
            .O(N__6340),
            .I(\U712_CHIP_RAM.N_287 ));
    LocalMux I__1122 (
            .O(N__6337),
            .I(\U712_CHIP_RAM.N_287 ));
    LocalMux I__1121 (
            .O(N__6330),
            .I(\U712_CHIP_RAM.N_287 ));
    InMux I__1120 (
            .O(N__6317),
            .I(N__6314));
    LocalMux I__1119 (
            .O(N__6314),
            .I(N__6311));
    Span4Mux_v I__1118 (
            .O(N__6311),
            .I(N__6308));
    Odrv4 I__1117 (
            .O(N__6308),
            .I(\U712_CHIP_RAM.N_388 ));
    InMux I__1116 (
            .O(N__6305),
            .I(N__6302));
    LocalMux I__1115 (
            .O(N__6302),
            .I(\U712_CHIP_RAM.N_370 ));
    InMux I__1114 (
            .O(N__6299),
            .I(N__6296));
    LocalMux I__1113 (
            .O(N__6296),
            .I(\U712_BYTE_ENABLE.un1_CUUBEn_i_0_aZ0Z2 ));
    IoInMux I__1112 (
            .O(N__6293),
            .I(N__6290));
    LocalMux I__1111 (
            .O(N__6290),
            .I(N__6287));
    IoSpan4Mux I__1110 (
            .O(N__6287),
            .I(N__6284));
    Span4Mux_s1_h I__1109 (
            .O(N__6284),
            .I(N__6281));
    Span4Mux_v I__1108 (
            .O(N__6281),
            .I(N__6278));
    Sp12to4 I__1107 (
            .O(N__6278),
            .I(N__6275));
    Span12Mux_s10_h I__1106 (
            .O(N__6275),
            .I(N__6272));
    Odrv12 I__1105 (
            .O(N__6272),
            .I(N_38_i));
    CascadeMux I__1104 (
            .O(N__6269),
            .I(\U712_BYTE_ENABLE.N_426_cascade_ ));
    IoInMux I__1103 (
            .O(N__6266),
            .I(N__6263));
    LocalMux I__1102 (
            .O(N__6263),
            .I(N__6260));
    IoSpan4Mux I__1101 (
            .O(N__6260),
            .I(N__6257));
    Span4Mux_s1_h I__1100 (
            .O(N__6257),
            .I(N__6254));
    Sp12to4 I__1099 (
            .O(N__6254),
            .I(N__6251));
    Span12Mux_h I__1098 (
            .O(N__6251),
            .I(N__6248));
    Span12Mux_v I__1097 (
            .O(N__6248),
            .I(N__6245));
    Odrv12 I__1096 (
            .O(N__6245),
            .I(N_47_i));
    InMux I__1095 (
            .O(N__6242),
            .I(N__6239));
    LocalMux I__1094 (
            .O(N__6239),
            .I(N__6236));
    Odrv4 I__1093 (
            .O(N__6236),
            .I(\U712_BYTE_ENABLE.un1_CLMBEn_i_0_aZ0Z2 ));
    IoInMux I__1092 (
            .O(N__6233),
            .I(N__6230));
    LocalMux I__1091 (
            .O(N__6230),
            .I(N__6225));
    CascadeMux I__1090 (
            .O(N__6229),
            .I(N__6220));
    CascadeMux I__1089 (
            .O(N__6228),
            .I(N__6217));
    IoSpan4Mux I__1088 (
            .O(N__6225),
            .I(N__6214));
    InMux I__1087 (
            .O(N__6224),
            .I(N__6205));
    InMux I__1086 (
            .O(N__6223),
            .I(N__6205));
    InMux I__1085 (
            .O(N__6220),
            .I(N__6205));
    InMux I__1084 (
            .O(N__6217),
            .I(N__6205));
    Span4Mux_s3_v I__1083 (
            .O(N__6214),
            .I(N__6202));
    LocalMux I__1082 (
            .O(N__6205),
            .I(N__6199));
    Span4Mux_v I__1081 (
            .O(N__6202),
            .I(N__6195));
    Span4Mux_v I__1080 (
            .O(N__6199),
            .I(N__6192));
    InMux I__1079 (
            .O(N__6198),
            .I(N__6189));
    Odrv4 I__1078 (
            .O(N__6195),
            .I(DBENn_c));
    Odrv4 I__1077 (
            .O(N__6192),
            .I(DBENn_c));
    LocalMux I__1076 (
            .O(N__6189),
            .I(DBENn_c));
    IoInMux I__1075 (
            .O(N__6182),
            .I(N__6179));
    LocalMux I__1074 (
            .O(N__6179),
            .I(N__6176));
    Span4Mux_s2_h I__1073 (
            .O(N__6176),
            .I(N__6173));
    Span4Mux_h I__1072 (
            .O(N__6173),
            .I(N__6170));
    Sp12to4 I__1071 (
            .O(N__6170),
            .I(N__6167));
    Span12Mux_v I__1070 (
            .O(N__6167),
            .I(N__6164));
    Odrv12 I__1069 (
            .O(N__6164),
            .I(N_46_i));
    CascadeMux I__1068 (
            .O(N__6161),
            .I(\U712_CHIP_RAM.N_287_cascade_ ));
    InMux I__1067 (
            .O(N__6158),
            .I(N__6155));
    LocalMux I__1066 (
            .O(N__6155),
            .I(\U712_CHIP_RAM.N_436 ));
    CascadeMux I__1065 (
            .O(N__6152),
            .I(N__6148));
    InMux I__1064 (
            .O(N__6151),
            .I(N__6141));
    InMux I__1063 (
            .O(N__6148),
            .I(N__6141));
    InMux I__1062 (
            .O(N__6147),
            .I(N__6136));
    InMux I__1061 (
            .O(N__6146),
            .I(N__6136));
    LocalMux I__1060 (
            .O(N__6141),
            .I(N__6133));
    LocalMux I__1059 (
            .O(N__6136),
            .I(N__6130));
    Span4Mux_h I__1058 (
            .O(N__6133),
            .I(N__6127));
    Odrv4 I__1057 (
            .O(N__6130),
            .I(\U712_CHIP_RAM.N_283 ));
    Odrv4 I__1056 (
            .O(N__6127),
            .I(\U712_CHIP_RAM.N_283 ));
    CascadeMux I__1055 (
            .O(N__6122),
            .I(N__6119));
    InMux I__1054 (
            .O(N__6119),
            .I(N__6116));
    LocalMux I__1053 (
            .O(N__6116),
            .I(N__6113));
    Odrv12 I__1052 (
            .O(N__6113),
            .I(\U712_CHIP_RAM.N_347 ));
    InMux I__1051 (
            .O(N__6110),
            .I(N__6107));
    LocalMux I__1050 (
            .O(N__6107),
            .I(N__6104));
    Odrv4 I__1049 (
            .O(N__6104),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_i_0_2 ));
    CascadeMux I__1048 (
            .O(N__6101),
            .I(N__6098));
    InMux I__1047 (
            .O(N__6098),
            .I(N__6095));
    LocalMux I__1046 (
            .O(N__6095),
            .I(N__6092));
    Odrv4 I__1045 (
            .O(N__6092),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_129_i_0_0 ));
    CascadeMux I__1044 (
            .O(N__6089),
            .I(N__6084));
    InMux I__1043 (
            .O(N__6088),
            .I(N__6078));
    InMux I__1042 (
            .O(N__6087),
            .I(N__6075));
    InMux I__1041 (
            .O(N__6084),
            .I(N__6070));
    InMux I__1040 (
            .O(N__6083),
            .I(N__6059));
    InMux I__1039 (
            .O(N__6082),
            .I(N__6059));
    InMux I__1038 (
            .O(N__6081),
            .I(N__6059));
    LocalMux I__1037 (
            .O(N__6078),
            .I(N__6056));
    LocalMux I__1036 (
            .O(N__6075),
            .I(N__6053));
    InMux I__1035 (
            .O(N__6074),
            .I(N__6050));
    InMux I__1034 (
            .O(N__6073),
            .I(N__6047));
    LocalMux I__1033 (
            .O(N__6070),
            .I(N__6044));
    InMux I__1032 (
            .O(N__6069),
            .I(N__6039));
    InMux I__1031 (
            .O(N__6068),
            .I(N__6039));
    InMux I__1030 (
            .O(N__6067),
            .I(N__6034));
    InMux I__1029 (
            .O(N__6066),
            .I(N__6034));
    LocalMux I__1028 (
            .O(N__6059),
            .I(\U712_CHIP_RAM.N_286 ));
    Odrv4 I__1027 (
            .O(N__6056),
            .I(\U712_CHIP_RAM.N_286 ));
    Odrv4 I__1026 (
            .O(N__6053),
            .I(\U712_CHIP_RAM.N_286 ));
    LocalMux I__1025 (
            .O(N__6050),
            .I(\U712_CHIP_RAM.N_286 ));
    LocalMux I__1024 (
            .O(N__6047),
            .I(\U712_CHIP_RAM.N_286 ));
    Odrv12 I__1023 (
            .O(N__6044),
            .I(\U712_CHIP_RAM.N_286 ));
    LocalMux I__1022 (
            .O(N__6039),
            .I(\U712_CHIP_RAM.N_286 ));
    LocalMux I__1021 (
            .O(N__6034),
            .I(\U712_CHIP_RAM.N_286 ));
    CEMux I__1020 (
            .O(N__6017),
            .I(N__6014));
    LocalMux I__1019 (
            .O(N__6014),
            .I(N__6011));
    Odrv4 I__1018 (
            .O(N__6011),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ));
    CascadeMux I__1017 (
            .O(N__6008),
            .I(N__6005));
    InMux I__1016 (
            .O(N__6005),
            .I(N__6000));
    InMux I__1015 (
            .O(N__6004),
            .I(N__5997));
    InMux I__1014 (
            .O(N__6003),
            .I(N__5994));
    LocalMux I__1013 (
            .O(N__6000),
            .I(N__5988));
    LocalMux I__1012 (
            .O(N__5997),
            .I(N__5983));
    LocalMux I__1011 (
            .O(N__5994),
            .I(N__5983));
    InMux I__1010 (
            .O(N__5993),
            .I(N__5980));
    InMux I__1009 (
            .O(N__5992),
            .I(N__5977));
    InMux I__1008 (
            .O(N__5991),
            .I(N__5974));
    Span4Mux_h I__1007 (
            .O(N__5988),
            .I(N__5971));
    Span4Mux_h I__1006 (
            .O(N__5983),
            .I(N__5966));
    LocalMux I__1005 (
            .O(N__5980),
            .I(N__5966));
    LocalMux I__1004 (
            .O(N__5977),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1003 (
            .O(N__5974),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__1002 (
            .O(N__5971),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__1001 (
            .O(N__5966),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    CascadeMux I__1000 (
            .O(N__5957),
            .I(N__5954));
    InMux I__999 (
            .O(N__5954),
            .I(N__5950));
    InMux I__998 (
            .O(N__5953),
            .I(N__5945));
    LocalMux I__997 (
            .O(N__5950),
            .I(N__5942));
    InMux I__996 (
            .O(N__5949),
            .I(N__5939));
    InMux I__995 (
            .O(N__5948),
            .I(N__5936));
    LocalMux I__994 (
            .O(N__5945),
            .I(N__5929));
    Span4Mux_h I__993 (
            .O(N__5942),
            .I(N__5929));
    LocalMux I__992 (
            .O(N__5939),
            .I(N__5929));
    LocalMux I__991 (
            .O(N__5936),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__990 (
            .O(N__5929),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    CascadeMux I__989 (
            .O(N__5924),
            .I(N__5921));
    InMux I__988 (
            .O(N__5921),
            .I(N__5916));
    InMux I__987 (
            .O(N__5920),
            .I(N__5911));
    InMux I__986 (
            .O(N__5919),
            .I(N__5908));
    LocalMux I__985 (
            .O(N__5916),
            .I(N__5905));
    InMux I__984 (
            .O(N__5915),
            .I(N__5902));
    InMux I__983 (
            .O(N__5914),
            .I(N__5899));
    LocalMux I__982 (
            .O(N__5911),
            .I(N__5892));
    LocalMux I__981 (
            .O(N__5908),
            .I(N__5892));
    Span4Mux_h I__980 (
            .O(N__5905),
            .I(N__5892));
    LocalMux I__979 (
            .O(N__5902),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__978 (
            .O(N__5899),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    Odrv4 I__977 (
            .O(N__5892),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    InMux I__976 (
            .O(N__5885),
            .I(N__5880));
    InMux I__975 (
            .O(N__5884),
            .I(N__5877));
    InMux I__974 (
            .O(N__5883),
            .I(N__5874));
    LocalMux I__973 (
            .O(N__5880),
            .I(N__5866));
    LocalMux I__972 (
            .O(N__5877),
            .I(N__5863));
    LocalMux I__971 (
            .O(N__5874),
            .I(N__5860));
    InMux I__970 (
            .O(N__5873),
            .I(N__5857));
    InMux I__969 (
            .O(N__5872),
            .I(N__5854));
    InMux I__968 (
            .O(N__5871),
            .I(N__5851));
    InMux I__967 (
            .O(N__5870),
            .I(N__5846));
    InMux I__966 (
            .O(N__5869),
            .I(N__5846));
    Span4Mux_h I__965 (
            .O(N__5866),
            .I(N__5843));
    Span4Mux_h I__964 (
            .O(N__5863),
            .I(N__5836));
    Span4Mux_h I__963 (
            .O(N__5860),
            .I(N__5836));
    LocalMux I__962 (
            .O(N__5857),
            .I(N__5836));
    LocalMux I__961 (
            .O(N__5854),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__960 (
            .O(N__5851),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__959 (
            .O(N__5846),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    Odrv4 I__958 (
            .O(N__5843),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    Odrv4 I__957 (
            .O(N__5836),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    CascadeMux I__956 (
            .O(N__5825),
            .I(\U712_REG_SM.C1_SYNC_RNIAS4F1_0Z0Z_1_cascade_ ));
    InMux I__955 (
            .O(N__5822),
            .I(N__5819));
    LocalMux I__954 (
            .O(N__5819),
            .I(N__5816));
    Span4Mux_v I__953 (
            .O(N__5816),
            .I(N__5812));
    InMux I__952 (
            .O(N__5815),
            .I(N__5809));
    Sp12to4 I__951 (
            .O(N__5812),
            .I(N__5804));
    LocalMux I__950 (
            .O(N__5809),
            .I(N__5804));
    Odrv12 I__949 (
            .O(N__5804),
            .I(\U712_REG_SM.ASn_0_sqmuxa_1 ));
    InMux I__948 (
            .O(N__5801),
            .I(N__5798));
    LocalMux I__947 (
            .O(N__5798),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a2_0_1 ));
    CascadeMux I__946 (
            .O(N__5795),
            .I(N__5787));
    InMux I__945 (
            .O(N__5794),
            .I(N__5782));
    InMux I__944 (
            .O(N__5793),
            .I(N__5782));
    InMux I__943 (
            .O(N__5792),
            .I(N__5777));
    InMux I__942 (
            .O(N__5791),
            .I(N__5777));
    InMux I__941 (
            .O(N__5790),
            .I(N__5774));
    InMux I__940 (
            .O(N__5787),
            .I(N__5771));
    LocalMux I__939 (
            .O(N__5782),
            .I(N__5766));
    LocalMux I__938 (
            .O(N__5777),
            .I(N__5766));
    LocalMux I__937 (
            .O(N__5774),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__936 (
            .O(N__5771),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    Odrv12 I__935 (
            .O(N__5766),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    CascadeMux I__934 (
            .O(N__5759),
            .I(N__5756));
    InMux I__933 (
            .O(N__5756),
            .I(N__5752));
    CascadeMux I__932 (
            .O(N__5755),
            .I(N__5749));
    LocalMux I__931 (
            .O(N__5752),
            .I(N__5744));
    InMux I__930 (
            .O(N__5749),
            .I(N__5741));
    InMux I__929 (
            .O(N__5748),
            .I(N__5738));
    InMux I__928 (
            .O(N__5747),
            .I(N__5735));
    Span4Mux_h I__927 (
            .O(N__5744),
            .I(N__5732));
    LocalMux I__926 (
            .O(N__5741),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__925 (
            .O(N__5738),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__924 (
            .O(N__5735),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    Odrv4 I__923 (
            .O(N__5732),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    CascadeMux I__922 (
            .O(N__5723),
            .I(N__5719));
    InMux I__921 (
            .O(N__5722),
            .I(N__5716));
    InMux I__920 (
            .O(N__5719),
            .I(N__5713));
    LocalMux I__919 (
            .O(N__5716),
            .I(N__5707));
    LocalMux I__918 (
            .O(N__5713),
            .I(N__5707));
    InMux I__917 (
            .O(N__5712),
            .I(N__5704));
    Odrv12 I__916 (
            .O(N__5707),
            .I(\U712_REG_SM.C1_SYNC_RNIAS4F1_0Z0Z_1 ));
    LocalMux I__915 (
            .O(N__5704),
            .I(\U712_REG_SM.C1_SYNC_RNIAS4F1_0Z0Z_1 ));
    CascadeMux I__914 (
            .O(N__5699),
            .I(N__5696));
    InMux I__913 (
            .O(N__5696),
            .I(N__5693));
    LocalMux I__912 (
            .O(N__5693),
            .I(N__5690));
    Odrv4 I__911 (
            .O(N__5690),
            .I(\U712_REG_SM.N_104 ));
    CascadeMux I__910 (
            .O(N__5687),
            .I(\U712_CHIP_RAM.N_414_cascade_ ));
    InMux I__909 (
            .O(N__5684),
            .I(N__5681));
    LocalMux I__908 (
            .O(N__5681),
            .I(N__5678));
    Span4Mux_h I__907 (
            .O(N__5678),
            .I(N__5675));
    Odrv4 I__906 (
            .O(N__5675),
            .I(\U712_CHIP_RAM.N_86 ));
    InMux I__905 (
            .O(N__5672),
            .I(N__5666));
    InMux I__904 (
            .O(N__5671),
            .I(N__5663));
    InMux I__903 (
            .O(N__5670),
            .I(N__5660));
    CascadeMux I__902 (
            .O(N__5669),
            .I(N__5657));
    LocalMux I__901 (
            .O(N__5666),
            .I(N__5654));
    LocalMux I__900 (
            .O(N__5663),
            .I(N__5651));
    LocalMux I__899 (
            .O(N__5660),
            .I(N__5648));
    InMux I__898 (
            .O(N__5657),
            .I(N__5644));
    Span4Mux_v I__897 (
            .O(N__5654),
            .I(N__5641));
    Span4Mux_v I__896 (
            .O(N__5651),
            .I(N__5636));
    Span4Mux_h I__895 (
            .O(N__5648),
            .I(N__5636));
    InMux I__894 (
            .O(N__5647),
            .I(N__5633));
    LocalMux I__893 (
            .O(N__5644),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__892 (
            .O(N__5641),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__891 (
            .O(N__5636),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__890 (
            .O(N__5633),
            .I(DBR_SYNCZ0Z_1));
    CascadeMux I__889 (
            .O(N__5624),
            .I(N__5621));
    InMux I__888 (
            .O(N__5621),
            .I(N__5614));
    InMux I__887 (
            .O(N__5620),
            .I(N__5611));
    InMux I__886 (
            .O(N__5619),
            .I(N__5608));
    InMux I__885 (
            .O(N__5618),
            .I(N__5605));
    InMux I__884 (
            .O(N__5617),
            .I(N__5602));
    LocalMux I__883 (
            .O(N__5614),
            .I(N__5599));
    LocalMux I__882 (
            .O(N__5611),
            .I(N__5596));
    LocalMux I__881 (
            .O(N__5608),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__880 (
            .O(N__5605),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__879 (
            .O(N__5602),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    Odrv4 I__878 (
            .O(N__5599),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    Odrv12 I__877 (
            .O(N__5596),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    InMux I__876 (
            .O(N__5585),
            .I(N__5579));
    InMux I__875 (
            .O(N__5584),
            .I(N__5579));
    LocalMux I__874 (
            .O(N__5579),
            .I(N__5576));
    Odrv4 I__873 (
            .O(N__5576),
            .I(\U712_CHIP_RAM.N_373 ));
    InMux I__872 (
            .O(N__5573),
            .I(N__5569));
    InMux I__871 (
            .O(N__5572),
            .I(N__5564));
    LocalMux I__870 (
            .O(N__5569),
            .I(N__5560));
    InMux I__869 (
            .O(N__5568),
            .I(N__5555));
    InMux I__868 (
            .O(N__5567),
            .I(N__5555));
    LocalMux I__867 (
            .O(N__5564),
            .I(N__5552));
    InMux I__866 (
            .O(N__5563),
            .I(N__5549));
    Span4Mux_v I__865 (
            .O(N__5560),
            .I(N__5544));
    LocalMux I__864 (
            .O(N__5555),
            .I(N__5544));
    Odrv4 I__863 (
            .O(N__5552),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    LocalMux I__862 (
            .O(N__5549),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    Odrv4 I__861 (
            .O(N__5544),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    CascadeMux I__860 (
            .O(N__5537),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15_cascade_ ));
    InMux I__859 (
            .O(N__5534),
            .I(N__5531));
    LocalMux I__858 (
            .O(N__5531),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_1 ));
    CascadeMux I__857 (
            .O(N__5528),
            .I(\U712_CHIP_RAM.N_286_cascade_ ));
    InMux I__856 (
            .O(N__5525),
            .I(N__5522));
    LocalMux I__855 (
            .O(N__5522),
            .I(N__5517));
    InMux I__854 (
            .O(N__5521),
            .I(N__5512));
    InMux I__853 (
            .O(N__5520),
            .I(N__5512));
    Odrv4 I__852 (
            .O(N__5517),
            .I(\U712_CHIP_RAM.N_486 ));
    LocalMux I__851 (
            .O(N__5512),
            .I(\U712_CHIP_RAM.N_486 ));
    InMux I__850 (
            .O(N__5507),
            .I(N__5504));
    LocalMux I__849 (
            .O(N__5504),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a2_1 ));
    CascadeMux I__848 (
            .O(N__5501),
            .I(\U712_CHIP_RAM.N_371_1_cascade_ ));
    InMux I__847 (
            .O(N__5498),
            .I(N__5495));
    LocalMux I__846 (
            .O(N__5495),
            .I(N__5492));
    Span4Mux_v I__845 (
            .O(N__5492),
            .I(N__5489));
    Span4Mux_h I__844 (
            .O(N__5489),
            .I(N__5486));
    Odrv4 I__843 (
            .O(N__5486),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_a2_0 ));
    CascadeMux I__842 (
            .O(N__5483),
            .I(N__5480));
    InMux I__841 (
            .O(N__5480),
            .I(N__5477));
    LocalMux I__840 (
            .O(N__5477),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_0_0_0 ));
    InMux I__839 (
            .O(N__5474),
            .I(N__5471));
    LocalMux I__838 (
            .O(N__5471),
            .I(\U712_CHIP_RAM.N_371_1 ));
    InMux I__837 (
            .O(N__5468),
            .I(N__5465));
    LocalMux I__836 (
            .O(N__5465),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    CascadeMux I__835 (
            .O(N__5462),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_ ));
    CascadeMux I__834 (
            .O(N__5459),
            .I(N__5456));
    InMux I__833 (
            .O(N__5456),
            .I(N__5449));
    InMux I__832 (
            .O(N__5455),
            .I(N__5449));
    InMux I__831 (
            .O(N__5454),
            .I(N__5439));
    LocalMux I__830 (
            .O(N__5449),
            .I(N__5436));
    InMux I__829 (
            .O(N__5448),
            .I(N__5433));
    InMux I__828 (
            .O(N__5447),
            .I(N__5430));
    InMux I__827 (
            .O(N__5446),
            .I(N__5427));
    InMux I__826 (
            .O(N__5445),
            .I(N__5424));
    InMux I__825 (
            .O(N__5444),
            .I(N__5417));
    InMux I__824 (
            .O(N__5443),
            .I(N__5417));
    InMux I__823 (
            .O(N__5442),
            .I(N__5417));
    LocalMux I__822 (
            .O(N__5439),
            .I(N__5414));
    Span4Mux_h I__821 (
            .O(N__5436),
            .I(N__5411));
    LocalMux I__820 (
            .O(N__5433),
            .I(\U712_CHIP_RAM.N_288 ));
    LocalMux I__819 (
            .O(N__5430),
            .I(\U712_CHIP_RAM.N_288 ));
    LocalMux I__818 (
            .O(N__5427),
            .I(\U712_CHIP_RAM.N_288 ));
    LocalMux I__817 (
            .O(N__5424),
            .I(\U712_CHIP_RAM.N_288 ));
    LocalMux I__816 (
            .O(N__5417),
            .I(\U712_CHIP_RAM.N_288 ));
    Odrv4 I__815 (
            .O(N__5414),
            .I(\U712_CHIP_RAM.N_288 ));
    Odrv4 I__814 (
            .O(N__5411),
            .I(\U712_CHIP_RAM.N_288 ));
    CEMux I__813 (
            .O(N__5396),
            .I(N__5393));
    LocalMux I__812 (
            .O(N__5393),
            .I(N__5390));
    Span4Mux_v I__811 (
            .O(N__5390),
            .I(N__5387));
    Odrv4 I__810 (
            .O(N__5387),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0 ));
    InMux I__809 (
            .O(N__5384),
            .I(N__5381));
    LocalMux I__808 (
            .O(N__5381),
            .I(\U712_CHIP_RAM.N_329 ));
    InMux I__807 (
            .O(N__5378),
            .I(N__5375));
    LocalMux I__806 (
            .O(N__5375),
            .I(\U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ));
    CascadeMux I__805 (
            .O(N__5372),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_i_0_cascade_ ));
    InMux I__804 (
            .O(N__5369),
            .I(N__5366));
    LocalMux I__803 (
            .O(N__5366),
            .I(N__5362));
    InMux I__802 (
            .O(N__5365),
            .I(N__5359));
    Odrv4 I__801 (
            .O(N__5362),
            .I(\U712_CHIP_RAM.N_11_2 ));
    LocalMux I__800 (
            .O(N__5359),
            .I(\U712_CHIP_RAM.N_11_2 ));
    InMux I__799 (
            .O(N__5354),
            .I(N__5350));
    InMux I__798 (
            .O(N__5353),
            .I(N__5347));
    LocalMux I__797 (
            .O(N__5350),
            .I(N__5344));
    LocalMux I__796 (
            .O(N__5347),
            .I(REG_TACK));
    Odrv4 I__795 (
            .O(N__5344),
            .I(REG_TACK));
    InMux I__794 (
            .O(N__5339),
            .I(N__5333));
    InMux I__793 (
            .O(N__5338),
            .I(N__5333));
    LocalMux I__792 (
            .O(N__5333),
            .I(CPU_TACKm));
    CascadeMux I__791 (
            .O(N__5330),
            .I(N__5327));
    InMux I__790 (
            .O(N__5327),
            .I(N__5322));
    InMux I__789 (
            .O(N__5326),
            .I(N__5319));
    InMux I__788 (
            .O(N__5325),
            .I(N__5316));
    LocalMux I__787 (
            .O(N__5322),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    LocalMux I__786 (
            .O(N__5319),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    LocalMux I__785 (
            .O(N__5316),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    CascadeMux I__784 (
            .O(N__5309),
            .I(N__5306));
    InMux I__783 (
            .O(N__5306),
            .I(N__5302));
    InMux I__782 (
            .O(N__5305),
            .I(N__5299));
    LocalMux I__781 (
            .O(N__5302),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    LocalMux I__780 (
            .O(N__5299),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    CascadeMux I__779 (
            .O(N__5294),
            .I(\U712_CYCLE_TERM.TACK_EN6_0_cascade_ ));
    InMux I__778 (
            .O(N__5291),
            .I(N__5286));
    InMux I__777 (
            .O(N__5290),
            .I(N__5283));
    InMux I__776 (
            .O(N__5289),
            .I(N__5280));
    LocalMux I__775 (
            .O(N__5286),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__774 (
            .O(N__5283),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__773 (
            .O(N__5280),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    InMux I__772 (
            .O(N__5273),
            .I(N__5270));
    LocalMux I__771 (
            .O(N__5270),
            .I(\U712_CYCLE_TERM.N_316_i_0_en ));
    CEMux I__770 (
            .O(N__5267),
            .I(N__5264));
    LocalMux I__769 (
            .O(N__5264),
            .I(\U712_CYCLE_TERM.N_316_i_0_en_0 ));
    InMux I__768 (
            .O(N__5261),
            .I(N__5258));
    LocalMux I__767 (
            .O(N__5258),
            .I(N__5254));
    InMux I__766 (
            .O(N__5257),
            .I(N__5251));
    Odrv4 I__765 (
            .O(N__5254),
            .I(\U712_BYTE_ENABLE.N_282_i ));
    LocalMux I__764 (
            .O(N__5251),
            .I(\U712_BYTE_ENABLE.N_282_i ));
    InMux I__763 (
            .O(N__5246),
            .I(N__5243));
    LocalMux I__762 (
            .O(N__5243),
            .I(N__5240));
    Span12Mux_v I__761 (
            .O(N__5240),
            .I(N__5237));
    Span12Mux_h I__760 (
            .O(N__5237),
            .I(N__5234));
    Odrv12 I__759 (
            .O(N__5234),
            .I(A_c_4));
    InMux I__758 (
            .O(N__5231),
            .I(N__5228));
    LocalMux I__757 (
            .O(N__5228),
            .I(N__5225));
    Span4Mux_v I__756 (
            .O(N__5225),
            .I(N__5222));
    Sp12to4 I__755 (
            .O(N__5222),
            .I(N__5219));
    Span12Mux_h I__754 (
            .O(N__5219),
            .I(N__5216));
    Odrv12 I__753 (
            .O(N__5216),
            .I(A_c_11));
    InMux I__752 (
            .O(N__5213),
            .I(N__5210));
    LocalMux I__751 (
            .O(N__5210),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ));
    CascadeMux I__750 (
            .O(N__5207),
            .I(\U712_CHIP_RAM.N_15_cascade_ ));
    InMux I__749 (
            .O(N__5204),
            .I(N__5201));
    LocalMux I__748 (
            .O(N__5201),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_0_0 ));
    InMux I__747 (
            .O(N__5198),
            .I(N__5195));
    LocalMux I__746 (
            .O(N__5195),
            .I(N__5192));
    Span4Mux_v I__745 (
            .O(N__5192),
            .I(N__5189));
    Span4Mux_v I__744 (
            .O(N__5189),
            .I(N__5186));
    Sp12to4 I__743 (
            .O(N__5186),
            .I(N__5183));
    Odrv12 I__742 (
            .O(N__5183),
            .I(A_c_5));
    InMux I__741 (
            .O(N__5180),
            .I(N__5177));
    LocalMux I__740 (
            .O(N__5177),
            .I(N__5174));
    Span4Mux_v I__739 (
            .O(N__5174),
            .I(N__5171));
    Span4Mux_h I__738 (
            .O(N__5171),
            .I(N__5168));
    Sp12to4 I__737 (
            .O(N__5168),
            .I(N__5165));
    Odrv12 I__736 (
            .O(N__5165),
            .I(A_c_12));
    CascadeMux I__735 (
            .O(N__5162),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ));
    InMux I__734 (
            .O(N__5159),
            .I(N__5156));
    LocalMux I__733 (
            .O(N__5156),
            .I(N__5153));
    Odrv4 I__732 (
            .O(N__5153),
            .I(\U712_CHIP_RAM.N_448 ));
    CascadeMux I__731 (
            .O(N__5150),
            .I(\U712_CHIP_RAM.N_345_cascade_ ));
    InMux I__730 (
            .O(N__5147),
            .I(N__5144));
    LocalMux I__729 (
            .O(N__5144),
            .I(N__5141));
    Span12Mux_h I__728 (
            .O(N__5141),
            .I(N__5138));
    Span12Mux_v I__727 (
            .O(N__5138),
            .I(N__5135));
    Odrv12 I__726 (
            .O(N__5135),
            .I(A_c_2));
    InMux I__725 (
            .O(N__5132),
            .I(N__5129));
    LocalMux I__724 (
            .O(N__5129),
            .I(N__5126));
    Span4Mux_v I__723 (
            .O(N__5126),
            .I(N__5123));
    Sp12to4 I__722 (
            .O(N__5123),
            .I(N__5120));
    Odrv12 I__721 (
            .O(N__5120),
            .I(A_c_9));
    CascadeMux I__720 (
            .O(N__5117),
            .I(\U712_CHIP_RAM.N_288_cascade_ ));
    CascadeMux I__719 (
            .O(N__5114),
            .I(\U712_CHIP_RAM.N_372_cascade_ ));
    InMux I__718 (
            .O(N__5111),
            .I(N__5108));
    LocalMux I__717 (
            .O(N__5108),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0 ));
    CascadeMux I__716 (
            .O(N__5105),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_ ));
    CascadeMux I__715 (
            .O(N__5102),
            .I(N__5099));
    InMux I__714 (
            .O(N__5099),
            .I(N__5096));
    LocalMux I__713 (
            .O(N__5096),
            .I(N__5087));
    InMux I__712 (
            .O(N__5095),
            .I(N__5084));
    InMux I__711 (
            .O(N__5094),
            .I(N__5081));
    InMux I__710 (
            .O(N__5093),
            .I(N__5076));
    InMux I__709 (
            .O(N__5092),
            .I(N__5076));
    InMux I__708 (
            .O(N__5091),
            .I(N__5071));
    InMux I__707 (
            .O(N__5090),
            .I(N__5071));
    Odrv4 I__706 (
            .O(N__5087),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3 ));
    LocalMux I__705 (
            .O(N__5084),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3 ));
    LocalMux I__704 (
            .O(N__5081),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3 ));
    LocalMux I__703 (
            .O(N__5076),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3 ));
    LocalMux I__702 (
            .O(N__5071),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3 ));
    CascadeMux I__701 (
            .O(N__5060),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1_1_cascade_ ));
    CascadeMux I__700 (
            .O(N__5057),
            .I(\U712_CHIP_RAM.N_366_cascade_ ));
    CascadeMux I__699 (
            .O(N__5054),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_0_cascade_ ));
    IoInMux I__698 (
            .O(N__5051),
            .I(N__5048));
    LocalMux I__697 (
            .O(N__5048),
            .I(N__5045));
    Span4Mux_s0_v I__696 (
            .O(N__5045),
            .I(N__5042));
    Sp12to4 I__695 (
            .O(N__5042),
            .I(N__5038));
    InMux I__694 (
            .O(N__5041),
            .I(N__5035));
    Span12Mux_h I__693 (
            .O(N__5038),
            .I(N__5032));
    LocalMux I__692 (
            .O(N__5035),
            .I(N__5029));
    Odrv12 I__691 (
            .O(N__5032),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__690 (
            .O(N__5029),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__689 (
            .O(N__5024),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_cascade_ ));
    CascadeMux I__688 (
            .O(N__5021),
            .I(N__5017));
    InMux I__687 (
            .O(N__5020),
            .I(N__5012));
    InMux I__686 (
            .O(N__5017),
            .I(N__5012));
    LocalMux I__685 (
            .O(N__5012),
            .I(N__5009));
    Odrv4 I__684 (
            .O(N__5009),
            .I(\U712_CHIP_RAM.N_304 ));
    CascadeMux I__683 (
            .O(N__5006),
            .I(\U712_CHIP_RAM.N_62_cascade_ ));
    CascadeMux I__682 (
            .O(N__5003),
            .I(N__4999));
    InMux I__681 (
            .O(N__5002),
            .I(N__4995));
    InMux I__680 (
            .O(N__4999),
            .I(N__4992));
    InMux I__679 (
            .O(N__4998),
            .I(N__4989));
    LocalMux I__678 (
            .O(N__4995),
            .I(\U712_CHIP_RAM.N_452 ));
    LocalMux I__677 (
            .O(N__4992),
            .I(\U712_CHIP_RAM.N_452 ));
    LocalMux I__676 (
            .O(N__4989),
            .I(\U712_CHIP_RAM.N_452 ));
    CascadeMux I__675 (
            .O(N__4982),
            .I(\U712_CHIP_RAM.N_452_cascade_ ));
    InMux I__674 (
            .O(N__4979),
            .I(N__4974));
    InMux I__673 (
            .O(N__4978),
            .I(N__4971));
    InMux I__672 (
            .O(N__4977),
            .I(N__4968));
    LocalMux I__671 (
            .O(N__4974),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    LocalMux I__670 (
            .O(N__4971),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    LocalMux I__669 (
            .O(N__4968),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    CascadeMux I__668 (
            .O(N__4961),
            .I(\U712_CHIP_RAM.N_11_cascade_ ));
    IoInMux I__667 (
            .O(N__4958),
            .I(N__4955));
    LocalMux I__666 (
            .O(N__4955),
            .I(N__4952));
    Span4Mux_s0_h I__665 (
            .O(N__4952),
            .I(N__4949));
    Sp12to4 I__664 (
            .O(N__4949),
            .I(N__4946));
    Span12Mux_v I__663 (
            .O(N__4946),
            .I(N__4943));
    Span12Mux_h I__662 (
            .O(N__4943),
            .I(N__4939));
    InMux I__661 (
            .O(N__4942),
            .I(N__4936));
    Odrv12 I__660 (
            .O(N__4939),
            .I(CLK_EN_c));
    LocalMux I__659 (
            .O(N__4936),
            .I(CLK_EN_c));
    InMux I__658 (
            .O(N__4931),
            .I(N__4927));
    InMux I__657 (
            .O(N__4930),
            .I(N__4924));
    LocalMux I__656 (
            .O(N__4927),
            .I(DBR_SYNCZ0Z_0));
    LocalMux I__655 (
            .O(N__4924),
            .I(DBR_SYNCZ0Z_0));
    InMux I__654 (
            .O(N__4919),
            .I(N__4907));
    InMux I__653 (
            .O(N__4918),
            .I(N__4907));
    InMux I__652 (
            .O(N__4917),
            .I(N__4907));
    InMux I__651 (
            .O(N__4916),
            .I(N__4907));
    LocalMux I__650 (
            .O(N__4907),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    InMux I__649 (
            .O(N__4904),
            .I(N__4897));
    InMux I__648 (
            .O(N__4903),
            .I(N__4897));
    InMux I__647 (
            .O(N__4902),
            .I(N__4894));
    LocalMux I__646 (
            .O(N__4897),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__645 (
            .O(N__4894),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    IoInMux I__644 (
            .O(N__4889),
            .I(N__4886));
    LocalMux I__643 (
            .O(N__4886),
            .I(N__4883));
    Span4Mux_s0_h I__642 (
            .O(N__4883),
            .I(N__4880));
    Sp12to4 I__641 (
            .O(N__4880),
            .I(N__4877));
    Span12Mux_v I__640 (
            .O(N__4877),
            .I(N__4873));
    InMux I__639 (
            .O(N__4876),
            .I(N__4870));
    Odrv12 I__638 (
            .O(N__4873),
            .I(TACK_OUTn));
    LocalMux I__637 (
            .O(N__4870),
            .I(TACK_OUTn));
    InMux I__636 (
            .O(N__4865),
            .I(N__4862));
    LocalMux I__635 (
            .O(N__4862),
            .I(N__4859));
    Span4Mux_h I__634 (
            .O(N__4859),
            .I(N__4856));
    Span4Mux_v I__633 (
            .O(N__4856),
            .I(N__4853));
    Odrv4 I__632 (
            .O(N__4853),
            .I(TACK_EN_i_ess));
    InMux I__631 (
            .O(N__4850),
            .I(N__4847));
    LocalMux I__630 (
            .O(N__4847),
            .I(N__4844));
    Sp12to4 I__629 (
            .O(N__4844),
            .I(N__4841));
    Span12Mux_v I__628 (
            .O(N__4841),
            .I(N__4838));
    Span12Mux_h I__627 (
            .O(N__4838),
            .I(N__4835));
    Odrv12 I__626 (
            .O(N__4835),
            .I(A_c_18));
    InMux I__625 (
            .O(N__4832),
            .I(N__4829));
    LocalMux I__624 (
            .O(N__4829),
            .I(N__4826));
    Sp12to4 I__623 (
            .O(N__4826),
            .I(N__4823));
    Span12Mux_v I__622 (
            .O(N__4823),
            .I(N__4820));
    Span12Mux_h I__621 (
            .O(N__4820),
            .I(N__4817));
    Odrv12 I__620 (
            .O(N__4817),
            .I(A_c_16));
    InMux I__619 (
            .O(N__4814),
            .I(N__4810));
    InMux I__618 (
            .O(N__4813),
            .I(N__4807));
    LocalMux I__617 (
            .O(N__4810),
            .I(\U712_CHIP_RAM.N_489 ));
    LocalMux I__616 (
            .O(N__4807),
            .I(\U712_CHIP_RAM.N_489 ));
    InMux I__615 (
            .O(N__4802),
            .I(N__4799));
    LocalMux I__614 (
            .O(N__4799),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0 ));
    InMux I__613 (
            .O(N__4796),
            .I(N__4793));
    LocalMux I__612 (
            .O(N__4793),
            .I(N__4789));
    InMux I__611 (
            .O(N__4792),
            .I(N__4786));
    Span4Mux_h I__610 (
            .O(N__4789),
            .I(N__4781));
    LocalMux I__609 (
            .O(N__4786),
            .I(N__4781));
    Span4Mux_v I__608 (
            .O(N__4781),
            .I(N__4778));
    Sp12to4 I__607 (
            .O(N__4778),
            .I(N__4775));
    Span12Mux_h I__606 (
            .O(N__4775),
            .I(N__4772));
    Span12Mux_v I__605 (
            .O(N__4772),
            .I(N__4769));
    Odrv12 I__604 (
            .O(N__4769),
            .I(TSn_c));
    CascadeMux I__603 (
            .O(N__4766),
            .I(N__4763));
    InMux I__602 (
            .O(N__4763),
            .I(N__4760));
    LocalMux I__601 (
            .O(N__4760),
            .I(N__4757));
    Span12Mux_h I__600 (
            .O(N__4757),
            .I(N__4754));
    Span12Mux_v I__599 (
            .O(N__4754),
            .I(N__4751));
    Odrv12 I__598 (
            .O(N__4751),
            .I(RAMSPACEn_c));
    InMux I__597 (
            .O(N__4748),
            .I(N__4744));
    InMux I__596 (
            .O(N__4747),
            .I(N__4741));
    LocalMux I__595 (
            .O(N__4744),
            .I(N__4738));
    LocalMux I__594 (
            .O(N__4741),
            .I(N__4735));
    Span4Mux_v I__593 (
            .O(N__4738),
            .I(N__4732));
    Span4Mux_v I__592 (
            .O(N__4735),
            .I(N__4729));
    Sp12to4 I__591 (
            .O(N__4732),
            .I(N__4726));
    Span4Mux_h I__590 (
            .O(N__4729),
            .I(N__4723));
    Span12Mux_h I__589 (
            .O(N__4726),
            .I(N__4718));
    Sp12to4 I__588 (
            .O(N__4723),
            .I(N__4718));
    Span12Mux_v I__587 (
            .O(N__4718),
            .I(N__4715));
    Odrv12 I__586 (
            .O(N__4715),
            .I(AWEn_c));
    IoInMux I__585 (
            .O(N__4712),
            .I(N__4709));
    LocalMux I__584 (
            .O(N__4709),
            .I(N__4706));
    Span4Mux_s2_v I__583 (
            .O(N__4706),
            .I(N__4703));
    Span4Mux_v I__582 (
            .O(N__4703),
            .I(N__4700));
    Span4Mux_v I__581 (
            .O(N__4700),
            .I(N__4696));
    InMux I__580 (
            .O(N__4699),
            .I(N__4693));
    Odrv4 I__579 (
            .O(N__4696),
            .I(DBDIR_c));
    LocalMux I__578 (
            .O(N__4693),
            .I(DBDIR_c));
    InMux I__577 (
            .O(N__4688),
            .I(N__4684));
    InMux I__576 (
            .O(N__4687),
            .I(N__4681));
    LocalMux I__575 (
            .O(N__4684),
            .I(\U712_REG_SM.STATE_COUNT_RNI4BRHZ0Z_3 ));
    LocalMux I__574 (
            .O(N__4681),
            .I(\U712_REG_SM.STATE_COUNT_RNI4BRHZ0Z_3 ));
    InMux I__573 (
            .O(N__4676),
            .I(N__4673));
    LocalMux I__572 (
            .O(N__4673),
            .I(\U712_REG_SM.N_400 ));
    InMux I__571 (
            .O(N__4670),
            .I(N__4667));
    LocalMux I__570 (
            .O(N__4667),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_12_0 ));
    IoInMux I__569 (
            .O(N__4664),
            .I(N__4661));
    LocalMux I__568 (
            .O(N__4661),
            .I(N__4658));
    IoSpan4Mux I__567 (
            .O(N__4658),
            .I(N__4655));
    Sp12to4 I__566 (
            .O(N__4655),
            .I(N__4652));
    Span12Mux_s6_v I__565 (
            .O(N__4652),
            .I(N__4649));
    Span12Mux_v I__564 (
            .O(N__4649),
            .I(N__4645));
    InMux I__563 (
            .O(N__4648),
            .I(N__4642));
    Odrv12 I__562 (
            .O(N__4645),
            .I(LATCH_CLK_c));
    LocalMux I__561 (
            .O(N__4642),
            .I(LATCH_CLK_c));
    InMux I__560 (
            .O(N__4637),
            .I(N__4633));
    InMux I__559 (
            .O(N__4636),
            .I(N__4630));
    LocalMux I__558 (
            .O(N__4633),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    LocalMux I__557 (
            .O(N__4630),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    InMux I__556 (
            .O(N__4625),
            .I(N__4622));
    LocalMux I__555 (
            .O(N__4622),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ));
    CascadeMux I__554 (
            .O(N__4619),
            .I(\U712_CHIP_RAM.N_361_cascade_ ));
    CascadeMux I__553 (
            .O(N__4616),
            .I(N__4613));
    InMux I__552 (
            .O(N__4613),
            .I(N__4610));
    LocalMux I__551 (
            .O(N__4610),
            .I(N__4607));
    Span4Mux_v I__550 (
            .O(N__4607),
            .I(N__4604));
    Sp12to4 I__549 (
            .O(N__4604),
            .I(N__4601));
    Span12Mux_h I__548 (
            .O(N__4601),
            .I(N__4598));
    Span12Mux_v I__547 (
            .O(N__4598),
            .I(N__4595));
    Odrv12 I__546 (
            .O(N__4595),
            .I(A_c_20));
    InMux I__545 (
            .O(N__4592),
            .I(N__4588));
    InMux I__544 (
            .O(N__4591),
            .I(N__4585));
    LocalMux I__543 (
            .O(N__4588),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    LocalMux I__542 (
            .O(N__4585),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    CascadeMux I__541 (
            .O(N__4580),
            .I(\U712_CHIP_RAM.N_416_cascade_ ));
    CascadeMux I__540 (
            .O(N__4577),
            .I(\U712_CHIP_RAM.BANK0_RNOZ0Z_0_cascade_ ));
    InMux I__539 (
            .O(N__4574),
            .I(N__4571));
    LocalMux I__538 (
            .O(N__4571),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_i_i_0 ));
    IoInMux I__537 (
            .O(N__4568),
            .I(N__4565));
    LocalMux I__536 (
            .O(N__4565),
            .I(N__4562));
    Span4Mux_s3_v I__535 (
            .O(N__4562),
            .I(N__4559));
    Span4Mux_v I__534 (
            .O(N__4559),
            .I(N__4556));
    Span4Mux_v I__533 (
            .O(N__4556),
            .I(N__4553));
    Span4Mux_h I__532 (
            .O(N__4553),
            .I(N__4549));
    InMux I__531 (
            .O(N__4552),
            .I(N__4546));
    Odrv4 I__530 (
            .O(N__4549),
            .I(BANK0_c));
    LocalMux I__529 (
            .O(N__4546),
            .I(BANK0_c));
    CascadeMux I__528 (
            .O(N__4541),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3_cascade_ ));
    CascadeMux I__527 (
            .O(N__4538),
            .I(\U712_CHIP_RAM.N_410_cascade_ ));
    IoInMux I__526 (
            .O(N__4535),
            .I(N__4532));
    LocalMux I__525 (
            .O(N__4532),
            .I(N__4529));
    IoSpan4Mux I__524 (
            .O(N__4529),
            .I(N__4526));
    Span4Mux_s3_h I__523 (
            .O(N__4526),
            .I(N__4522));
    InMux I__522 (
            .O(N__4525),
            .I(N__4519));
    Span4Mux_h I__521 (
            .O(N__4522),
            .I(N__4516));
    LocalMux I__520 (
            .O(N__4519),
            .I(N__4513));
    Sp12to4 I__519 (
            .O(N__4516),
            .I(N__4510));
    Span4Mux_v I__518 (
            .O(N__4513),
            .I(N__4507));
    Span12Mux_h I__517 (
            .O(N__4510),
            .I(N__4502));
    Sp12to4 I__516 (
            .O(N__4507),
            .I(N__4502));
    Span12Mux_h I__515 (
            .O(N__4502),
            .I(N__4499));
    Span12Mux_v I__514 (
            .O(N__4499),
            .I(N__4496));
    Odrv12 I__513 (
            .O(N__4496),
            .I(C3_c));
    CEMux I__512 (
            .O(N__4493),
            .I(N__4490));
    LocalMux I__511 (
            .O(N__4490),
            .I(N__4487));
    Odrv12 I__510 (
            .O(N__4487),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0 ));
    InMux I__509 (
            .O(N__4484),
            .I(N__4481));
    LocalMux I__508 (
            .O(N__4481),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0 ));
    InMux I__507 (
            .O(N__4478),
            .I(N__4475));
    LocalMux I__506 (
            .O(N__4475),
            .I(\U712_CHIP_RAM.N_409 ));
    InMux I__505 (
            .O(N__4472),
            .I(N__4468));
    InMux I__504 (
            .O(N__4471),
            .I(N__4465));
    LocalMux I__503 (
            .O(N__4468),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0_1 ));
    LocalMux I__502 (
            .O(N__4465),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0_1 ));
    CascadeMux I__501 (
            .O(N__4460),
            .I(\U712_CHIP_RAM.N_489_cascade_ ));
    CascadeMux I__500 (
            .O(N__4457),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_0_cascade_ ));
    CascadeMux I__499 (
            .O(N__4454),
            .I(\U712_REG_SM.N_346_cascade_ ));
    InMux I__498 (
            .O(N__4451),
            .I(N__4447));
    InMux I__497 (
            .O(N__4450),
            .I(N__4443));
    LocalMux I__496 (
            .O(N__4447),
            .I(N__4437));
    InMux I__495 (
            .O(N__4446),
            .I(N__4434));
    LocalMux I__494 (
            .O(N__4443),
            .I(N__4431));
    InMux I__493 (
            .O(N__4442),
            .I(N__4424));
    InMux I__492 (
            .O(N__4441),
            .I(N__4424));
    InMux I__491 (
            .O(N__4440),
            .I(N__4424));
    Odrv4 I__490 (
            .O(N__4437),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__489 (
            .O(N__4434),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    Odrv4 I__488 (
            .O(N__4431),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__487 (
            .O(N__4424),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    InMux I__486 (
            .O(N__4415),
            .I(N__4409));
    InMux I__485 (
            .O(N__4414),
            .I(N__4400));
    InMux I__484 (
            .O(N__4413),
            .I(N__4400));
    InMux I__483 (
            .O(N__4412),
            .I(N__4400));
    LocalMux I__482 (
            .O(N__4409),
            .I(N__4397));
    InMux I__481 (
            .O(N__4408),
            .I(N__4394));
    InMux I__480 (
            .O(N__4407),
            .I(N__4391));
    LocalMux I__479 (
            .O(N__4400),
            .I(N__4388));
    Span4Mux_h I__478 (
            .O(N__4397),
            .I(N__4385));
    LocalMux I__477 (
            .O(N__4394),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__476 (
            .O(N__4391),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    Odrv4 I__475 (
            .O(N__4388),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    Odrv4 I__474 (
            .O(N__4385),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    CascadeMux I__473 (
            .O(N__4376),
            .I(\U712_REG_SM.STATE_COUNT_srsts_i_i_0_o2_0_1_3_cascade_ ));
    InMux I__472 (
            .O(N__4373),
            .I(N__4370));
    LocalMux I__471 (
            .O(N__4370),
            .I(N__4366));
    InMux I__470 (
            .O(N__4369),
            .I(N__4363));
    Odrv4 I__469 (
            .O(N__4366),
            .I(\U712_REG_SM.N_342 ));
    LocalMux I__468 (
            .O(N__4363),
            .I(\U712_REG_SM.N_342 ));
    InMux I__467 (
            .O(N__4358),
            .I(N__4355));
    LocalMux I__466 (
            .O(N__4355),
            .I(\U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0_0 ));
    CascadeMux I__465 (
            .O(N__4352),
            .I(N__4349));
    InMux I__464 (
            .O(N__4349),
            .I(N__4346));
    LocalMux I__463 (
            .O(N__4346),
            .I(\U712_REG_SM.N_106 ));
    InMux I__462 (
            .O(N__4343),
            .I(N__4340));
    LocalMux I__461 (
            .O(N__4340),
            .I(\U712_REG_SM.N_379 ));
    InMux I__460 (
            .O(N__4337),
            .I(N__4333));
    InMux I__459 (
            .O(N__4336),
            .I(N__4330));
    LocalMux I__458 (
            .O(N__4333),
            .I(N__4326));
    LocalMux I__457 (
            .O(N__4330),
            .I(N__4323));
    InMux I__456 (
            .O(N__4329),
            .I(N__4320));
    Span4Mux_v I__455 (
            .O(N__4326),
            .I(N__4317));
    Span4Mux_v I__454 (
            .O(N__4323),
            .I(N__4312));
    LocalMux I__453 (
            .O(N__4320),
            .I(N__4312));
    Span4Mux_v I__452 (
            .O(N__4317),
            .I(N__4309));
    Span4Mux_v I__451 (
            .O(N__4312),
            .I(N__4306));
    Sp12to4 I__450 (
            .O(N__4309),
            .I(N__4301));
    Sp12to4 I__449 (
            .O(N__4306),
            .I(N__4301));
    Span12Mux_h I__448 (
            .O(N__4301),
            .I(N__4298));
    Odrv12 I__447 (
            .O(N__4298),
            .I(DBRn_c));
    IoInMux I__446 (
            .O(N__4295),
            .I(N__4292));
    LocalMux I__445 (
            .O(N__4292),
            .I(N__4289));
    Span4Mux_s2_v I__444 (
            .O(N__4289),
            .I(N__4285));
    InMux I__443 (
            .O(N__4288),
            .I(N__4282));
    Sp12to4 I__442 (
            .O(N__4285),
            .I(N__4279));
    LocalMux I__441 (
            .O(N__4282),
            .I(N__4275));
    Span12Mux_s9_h I__440 (
            .O(N__4279),
            .I(N__4272));
    CascadeMux I__439 (
            .O(N__4278),
            .I(N__4269));
    Span4Mux_v I__438 (
            .O(N__4275),
            .I(N__4266));
    Span12Mux_v I__437 (
            .O(N__4272),
            .I(N__4263));
    InMux I__436 (
            .O(N__4269),
            .I(N__4260));
    Span4Mux_v I__435 (
            .O(N__4266),
            .I(N__4257));
    Odrv12 I__434 (
            .O(N__4263),
            .I(REGENn_c));
    LocalMux I__433 (
            .O(N__4260),
            .I(REGENn_c));
    Odrv4 I__432 (
            .O(N__4257),
            .I(REGENn_c));
    IoInMux I__431 (
            .O(N__4250),
            .I(N__4247));
    LocalMux I__430 (
            .O(N__4247),
            .I(N__4244));
    Odrv12 I__429 (
            .O(N__4244),
            .I(VBENn_c));
    InMux I__428 (
            .O(N__4241),
            .I(N__4235));
    InMux I__427 (
            .O(N__4240),
            .I(N__4235));
    LocalMux I__426 (
            .O(N__4235),
            .I(\U712_REG_SM.N_319 ));
    IoInMux I__425 (
            .O(N__4232),
            .I(N__4229));
    LocalMux I__424 (
            .O(N__4229),
            .I(N__4226));
    Span4Mux_s1_v I__423 (
            .O(N__4226),
            .I(N__4223));
    Span4Mux_v I__422 (
            .O(N__4223),
            .I(N__4220));
    Sp12to4 I__421 (
            .O(N__4220),
            .I(N__4217));
    Span12Mux_h I__420 (
            .O(N__4217),
            .I(N__4214));
    Span12Mux_v I__419 (
            .O(N__4214),
            .I(N__4210));
    InMux I__418 (
            .O(N__4213),
            .I(N__4207));
    Odrv12 I__417 (
            .O(N__4210),
            .I(ASn_c));
    LocalMux I__416 (
            .O(N__4207),
            .I(ASn_c));
    CascadeMux I__415 (
            .O(N__4202),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_cascade_ ));
    InMux I__414 (
            .O(N__4199),
            .I(N__4196));
    LocalMux I__413 (
            .O(N__4196),
            .I(N__4193));
    Span4Mux_v I__412 (
            .O(N__4193),
            .I(N__4190));
    Odrv4 I__411 (
            .O(N__4190),
            .I(DBRn_c_i));
    CascadeMux I__410 (
            .O(N__4187),
            .I(N__4181));
    InMux I__409 (
            .O(N__4186),
            .I(N__4177));
    InMux I__408 (
            .O(N__4185),
            .I(N__4174));
    InMux I__407 (
            .O(N__4184),
            .I(N__4171));
    InMux I__406 (
            .O(N__4181),
            .I(N__4166));
    InMux I__405 (
            .O(N__4180),
            .I(N__4166));
    LocalMux I__404 (
            .O(N__4177),
            .I(\U712_REG_SM.C1_SYNC_RNIAS4F1Z0Z_1 ));
    LocalMux I__403 (
            .O(N__4174),
            .I(\U712_REG_SM.C1_SYNC_RNIAS4F1Z0Z_1 ));
    LocalMux I__402 (
            .O(N__4171),
            .I(\U712_REG_SM.C1_SYNC_RNIAS4F1Z0Z_1 ));
    LocalMux I__401 (
            .O(N__4166),
            .I(\U712_REG_SM.C1_SYNC_RNIAS4F1Z0Z_1 ));
    InMux I__400 (
            .O(N__4157),
            .I(N__4154));
    LocalMux I__399 (
            .O(N__4154),
            .I(N__4151));
    Odrv4 I__398 (
            .O(N__4151),
            .I(\U712_REG_SM.N_348 ));
    CascadeMux I__397 (
            .O(N__4148),
            .I(DBRn_c_i_cascade_));
    IoInMux I__396 (
            .O(N__4145),
            .I(N__4142));
    LocalMux I__395 (
            .O(N__4142),
            .I(N__4139));
    IoSpan4Mux I__394 (
            .O(N__4139),
            .I(N__4136));
    Span4Mux_s3_h I__393 (
            .O(N__4136),
            .I(N__4133));
    Span4Mux_h I__392 (
            .O(N__4133),
            .I(N__4130));
    Odrv4 I__391 (
            .O(N__4130),
            .I(DBRn_c_i_0));
    InMux I__390 (
            .O(N__4127),
            .I(N__4124));
    LocalMux I__389 (
            .O(N__4124),
            .I(N__4120));
    IoInMux I__388 (
            .O(N__4123),
            .I(N__4117));
    Span4Mux_v I__387 (
            .O(N__4120),
            .I(N__4114));
    LocalMux I__386 (
            .O(N__4117),
            .I(N__4111));
    Sp12to4 I__385 (
            .O(N__4114),
            .I(N__4108));
    IoSpan4Mux I__384 (
            .O(N__4111),
            .I(N__4105));
    Span12Mux_h I__383 (
            .O(N__4108),
            .I(N__4102));
    IoSpan4Mux I__382 (
            .O(N__4105),
            .I(N__4099));
    Span12Mux_v I__381 (
            .O(N__4102),
            .I(N__4096));
    IoSpan4Mux I__380 (
            .O(N__4099),
            .I(N__4093));
    Odrv12 I__379 (
            .O(N__4096),
            .I(C1_c));
    Odrv4 I__378 (
            .O(N__4093),
            .I(C1_c));
    InMux I__377 (
            .O(N__4088),
            .I(N__4082));
    InMux I__376 (
            .O(N__4087),
            .I(N__4082));
    LocalMux I__375 (
            .O(N__4082),
            .I(\U712_REG_SM.REG_CYCLE_START_RNITO6SZ0Z1 ));
    InMux I__374 (
            .O(N__4079),
            .I(N__4075));
    InMux I__373 (
            .O(N__4078),
            .I(N__4072));
    LocalMux I__372 (
            .O(N__4075),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    LocalMux I__371 (
            .O(N__4072),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    IoInMux I__370 (
            .O(N__4067),
            .I(N__4064));
    LocalMux I__369 (
            .O(N__4064),
            .I(N__4061));
    Span12Mux_s5_h I__368 (
            .O(N__4061),
            .I(N__4058));
    Odrv12 I__367 (
            .O(N__4058),
            .I(N_1062_i));
    IoInMux I__366 (
            .O(N__4055),
            .I(N__4052));
    LocalMux I__365 (
            .O(N__4052),
            .I(N__4049));
    Span4Mux_s3_v I__364 (
            .O(N__4049),
            .I(N__4046));
    Span4Mux_h I__363 (
            .O(N__4046),
            .I(N__4043));
    Odrv4 I__362 (
            .O(N__4043),
            .I(CLK80_PLL_i_i));
    CascadeMux I__361 (
            .O(N__4040),
            .I(N__4037));
    InMux I__360 (
            .O(N__4037),
            .I(N__4034));
    LocalMux I__359 (
            .O(N__4034),
            .I(N__4031));
    Span4Mux_h I__358 (
            .O(N__4031),
            .I(N__4028));
    Span4Mux_v I__357 (
            .O(N__4028),
            .I(N__4025));
    Span4Mux_v I__356 (
            .O(N__4025),
            .I(N__4022));
    Odrv4 I__355 (
            .O(N__4022),
            .I(REGSPACEn_c));
    InMux I__354 (
            .O(N__4019),
            .I(N__4014));
    InMux I__353 (
            .O(N__4018),
            .I(N__4009));
    InMux I__352 (
            .O(N__4017),
            .I(N__4009));
    LocalMux I__351 (
            .O(N__4014),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__350 (
            .O(N__4009),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    IoInMux I__349 (
            .O(N__4004),
            .I(N__4001));
    LocalMux I__348 (
            .O(N__4001),
            .I(N__3998));
    IoSpan4Mux I__347 (
            .O(N__3998),
            .I(N__3995));
    Span4Mux_s2_v I__346 (
            .O(N__3995),
            .I(N__3992));
    Sp12to4 I__345 (
            .O(N__3992),
            .I(N__3989));
    Span12Mux_v I__344 (
            .O(N__3989),
            .I(N__3986));
    Odrv12 I__343 (
            .O(N__3986),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .I(N__6732));
    INV \INVU712_CHIP_RAM.DMA_A1_nesrC  (
            .O(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .I(N__6729));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .I(N__6730));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .I(N__6731));
    INV \INVU712_CHIP_RAM.DMA_A20C  (
            .O(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .I(N__6734));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_7_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__8264),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__4123),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__4145),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__4535),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam TACKn_obuft_RNO_LC_2_15_6.C_ON=1'b0;
    defparam TACKn_obuft_RNO_LC_2_15_6.SEQ_MODE=4'b0000;
    defparam TACKn_obuft_RNO_LC_2_15_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 TACKn_obuft_RNO_LC_2_15_6 (
            .in0(N__4865),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_1062_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_3_1_0.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_3_1_0.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_3_1_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLKRAM_obuf_RNO_LC_3_1_0 (
            .in0(N__9821),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_5_6_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_5_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_5_6_6 .LUT_INIT=16'b0000010111001101;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_5_6_6  (
            .in0(N__4792),
            .in1(N__4019),
            .in2(N__4040),
            .in3(N__8126),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9810),
            .ce(),
            .sr(N__10806));
    defparam \U712_REG_SM.REG_CYCLE_START_RNITO6S1_LC_5_7_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNITO6S1_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNITO6S1_LC_5_7_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNITO6S1_LC_5_7_4  (
            .in0(_gnd_net_),
            .in1(N__4017),
            .in2(_gnd_net_),
            .in3(N__4180),
            .lcout(\U712_REG_SM.REG_CYCLE_START_RNITO6SZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_5_7_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_5_7_7 .LUT_INIT=16'b1100010011110111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_5_7_7  (
            .in0(N__4018),
            .in1(N__4078),
            .in2(N__4187),
            .in3(N__4408),
            .lcout(\U712_REG_SM.N_348 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_5_8_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_5_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_5_8_1 .LUT_INIT=16'b0011000000110010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_5_8_1  (
            .in0(N__5748),
            .in1(N__5722),
            .in2(N__5795),
            .in3(N__4186),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9817),
            .ce(),
            .sr(N__10805));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_5_8_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_5_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_5_8_4 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_5_8_4  (
            .in0(N__6004),
            .in1(N__5884),
            .in2(N__6755),
            .in3(N__4157),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9817),
            .ce(),
            .sr(N__10805));
    defparam \U712_REG_SM.STATE_COUNT_RNIBMB91_1_LC_5_9_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIBMB91_1_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIBMB91_1_LC_5_9_7 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIBMB91_1_LC_5_9_7  (
            .in0(N__4407),
            .in1(N__5885),
            .in2(N__6008),
            .in3(N__6747),
            .lcout(\U712_REG_SM.N_319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBRn_ibuf_RNIBAB_LC_5_10_6.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_5_10_6.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_5_10_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_5_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4337),
            .lcout(DBRn_c_i),
            .ltout(DBRn_c_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_10_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4148),
            .in3(N__10824),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_6_7_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_6_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_6_7_7 .LUT_INIT=16'b0111001000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_6_7_7  (
            .in0(N__4451),
            .in1(N__4373),
            .in2(N__5755),
            .in3(N__4185),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9808),
            .ce(),
            .sr(N__10800));
    defparam \U712_REG_SM.C1_SYNC_0_LC_6_8_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_6_8_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_6_8_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_6_8_0  (
            .in0(N__4127),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9811),
            .ce(),
            .sr(N__10793));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_6_8_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_6_8_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_6_8_2 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_6_8_2  (
            .in0(N__5790),
            .in1(N__4688),
            .in2(N__5723),
            .in3(N__4088),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9811),
            .ce(),
            .sr(N__10793));
    defparam \U712_REG_SM.REGENn_LC_6_8_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_LC_6_8_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_LC_6_8_4 .LUT_INIT=16'b1110101011111010;
    LogicCell40 \U712_REG_SM.REGENn_LC_6_8_4  (
            .in0(N__5815),
            .in1(N__4087),
            .in2(N__4278),
            .in3(N__4079),
            .lcout(REGENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9811),
            .ce(),
            .sr(N__10793));
    defparam \U712_REG_SM.C1_SYNC_RNIAS4F1_1_LC_6_8_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNIAS4F1_1_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNIAS4F1_1_LC_6_8_5 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNIAS4F1_1_LC_6_8_5  (
            .in0(N__5883),
            .in1(N__6003),
            .in2(N__5957),
            .in3(N__5914),
            .lcout(\U712_REG_SM.C1_SYNC_RNIAS4F1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_6_9_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_6_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_6_9_2 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_6_9_2  (
            .in0(N__4446),
            .in1(N__4369),
            .in2(_gnd_net_),
            .in3(N__4240),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9814),
            .ce(),
            .sr(N__10786));
    defparam \U712_REG_SM.ASn_LC_6_9_6 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_LC_6_9_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_LC_6_9_6 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \U712_REG_SM.ASn_LC_6_9_6  (
            .in0(N__4213),
            .in1(N__5822),
            .in2(_gnd_net_),
            .in3(N__4241),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9814),
            .ce(),
            .sr(N__10786));
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_7_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_7_6_0 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNO_0_LC_7_6_0  (
            .in0(N__7428),
            .in1(N__6151),
            .in2(N__5459),
            .in3(N__4478),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_LC_7_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_7_6_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_7_6_1 .LUT_INIT=16'b0011101011111010;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_7_6_1  (
            .in0(N__6198),
            .in1(N__5573),
            .in2(N__4202),
            .in3(N__8990),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9803),
            .ce(),
            .sr(N__10801));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_0_LC_7_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_0_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_0_LC_7_6_3 .LUT_INIT=16'b0000000010111010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_0_LC_7_6_3  (
            .in0(N__4472),
            .in1(N__7427),
            .in2(N__6152),
            .in3(N__5455),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_A20_LC_7_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A20_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A20_LC_7_7_0 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_A20_LC_7_7_0  (
            .in0(N__11153),
            .in1(N__4199),
            .in2(N__11075),
            .in3(N__4592),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .ce(),
            .sr(N__10794));
    defparam \U712_REG_SM.STATE_COUNT_RNI4BRH_3_LC_7_7_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI4BRH_3_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI4BRH_3_LC_7_7_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI4BRH_3_LC_7_7_1  (
            .in0(N__4415),
            .in1(N__5747),
            .in2(_gnd_net_),
            .in3(N__4450),
            .lcout(\U712_REG_SM.STATE_COUNT_RNI4BRHZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_7_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_7_8_1 .LUT_INIT=16'b1100110000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_7_8_1  (
            .in0(N__7869),
            .in1(N__7969),
            .in2(N__7150),
            .in3(N__7219),
            .lcout(\U712_CHIP_RAM.N_347 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_7_8_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_7_8_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_7_8_2  (
            .in0(N__4184),
            .in1(N__4413),
            .in2(_gnd_net_),
            .in3(N__4441),
            .lcout(\U712_REG_SM.N_400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_7_8_3 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_7_8_3 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_0_LC_7_8_3  (
            .in0(N__5870),
            .in1(N__6562),
            .in2(_gnd_net_),
            .in3(N__5793),
            .lcout(\U712_REG_SM.N_106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_3_LC_7_8_4 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_3_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_3_LC_7_8_4 .LUT_INIT=16'b0111011111101110;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_3_LC_7_8_4  (
            .in0(N__5991),
            .in1(N__4440),
            .in2(_gnd_net_),
            .in3(N__5869),
            .lcout(),
            .ltout(\U712_REG_SM.N_346_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_7_8_5 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_7_8_5 .LUT_INIT=16'b1111000111110101;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_2_LC_7_8_5  (
            .in0(N__4412),
            .in1(N__5919),
            .in2(N__4454),
            .in3(N__5953),
            .lcout(\U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_7_8_6 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_7_8_6 .LUT_INIT=16'b0001000000010001;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_1_LC_7_8_6  (
            .in0(N__5794),
            .in1(N__4442),
            .in2(N__6754),
            .in3(N__4414),
            .lcout(\U712_REG_SM.N_379 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNIS63V_1_LC_7_9_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNIS63V_1_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNIS63V_1_LC_7_9_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNIS63V_1_LC_7_9_1  (
            .in0(N__5948),
            .in1(N__5915),
            .in2(N__5669),
            .in3(N__4930),
            .lcout(),
            .ltout(\U712_REG_SM.STATE_COUNT_srsts_i_i_0_o2_0_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNI35EO1_1_LC_7_9_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI35EO1_1_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI35EO1_1_LC_7_9_2 .LUT_INIT=16'b1111001111111111;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI35EO1_1_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(N__5871),
            .in2(N__4376),
            .in3(N__5992),
            .lcout(\U712_REG_SM.N_342 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_LC_7_9_7 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_LC_7_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DS_EN_LC_7_9_7 .LUT_INIT=16'b1010101010001011;
    LogicCell40 \U712_REG_SM.DS_EN_LC_7_9_7  (
            .in0(N__10357),
            .in1(N__4358),
            .in2(N__4352),
            .in3(N__4343),
            .lcout(DS_ENm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9812),
            .ce(),
            .sr(N__10779));
    defparam DBR_SYNC_0_LC_7_10_2.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_7_10_2.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_7_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_0_LC_7_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4336),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9815),
            .ce(),
            .sr(N__10775));
    defparam \U712_REG_SM.REG_CYCLE_LC_7_16_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_7_16_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_7_16_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_7_16_7  (
            .in0(N__4329),
            .in1(N__8386),
            .in2(_gnd_net_),
            .in3(N__4288),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10889),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_0_a3_0_a2_LC_8_4_0 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a3_0_a2_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a3_0_a2_LC_8_4_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a3_0_a2_LC_8_4_0  (
            .in0(_gnd_net_),
            .in1(N__8125),
            .in2(_gnd_net_),
            .in3(N__9638),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_8_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_8_5_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_8_5_0  (
            .in0(N__4747),
            .in1(N__6554),
            .in2(_gnd_net_),
            .in3(N__7568),
            .lcout(WRITE_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9794),
            .ce(N__4493),
            .sr(N__10802));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_8_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_8_6_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_8_6_0  (
            .in0(_gnd_net_),
            .in1(N__10826),
            .in2(_gnd_net_),
            .in3(N__4977),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_8_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_8_6_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_8_6_1  (
            .in0(N__10825),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4484),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNISNC52_LC_8_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNISNC52_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNISNC52_LC_8_6_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNISNC52_LC_8_6_2  (
            .in0(N__7381),
            .in1(N__7740),
            .in2(N__7112),
            .in3(N__7245),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_RNO_1_LC_8_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNO_1_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNO_1_LC_8_6_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNO_1_LC_8_6_3  (
            .in0(N__7247),
            .in1(N__6377),
            .in2(_gnd_net_),
            .in3(N__5092),
            .lcout(\U712_CHIP_RAM.N_409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI71B91_LC_8_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI71B91_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI71B91_LC_8_6_4 .LUT_INIT=16'b1010111110101100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI71B91_LC_8_6_4  (
            .in0(N__7605),
            .in1(N__7950),
            .in2(N__7113),
            .in3(N__7246),
            .lcout(\U712_CHIP_RAM.N_304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIR9VE1_LC_8_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIR9VE1_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIR9VE1_LC_8_6_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIR9VE1_LC_8_6_5  (
            .in0(N__5617),
            .in1(N__6881),
            .in2(N__7567),
            .in3(N__5671),
            .lcout(\U712_CHIP_RAM.N_489 ),
            .ltout(\U712_CHIP_RAM.N_489_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_1_LC_8_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_1_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_1_LC_8_6_6 .LUT_INIT=16'b1100000011101010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_RNO_1_LC_8_6_6  (
            .in0(N__4471),
            .in1(N__4998),
            .in2(N__4460),
            .in3(N__5446),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_8_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_8_6_7 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_8_6_7  (
            .in0(N__7951),
            .in1(N__7079),
            .in2(N__4457),
            .in3(N__5093),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_3_LC_8_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_3_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_3_LC_8_7_0 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_3_LC_8_7_0  (
            .in0(N__7970),
            .in1(N__7269),
            .in2(N__7138),
            .in3(N__5095),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_361_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_8_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_8_7_1 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_1_LC_8_7_1  (
            .in0(N__6147),
            .in1(N__7434),
            .in2(N__4619),
            .in3(N__5444),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_i_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_2_LC_8_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_2_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_2_LC_8_7_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_2_LC_8_7_2  (
            .in0(N__11071),
            .in1(N__4813),
            .in2(N__4616),
            .in3(N__5567),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_416_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_8_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_8_7_3 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_0_LC_8_7_3  (
            .in0(N__5568),
            .in1(N__4591),
            .in2(N__4580),
            .in3(N__7562),
            .lcout(),
            .ltout(\U712_CHIP_RAM.BANK0_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_LC_8_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.BANK0_LC_8_7_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \U712_CHIP_RAM.BANK0_LC_8_7_4  (
            .in0(N__4552),
            .in1(N__4978),
            .in2(N__4577),
            .in3(N__4574),
            .lcout(BANK0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9804),
            .ce(),
            .sr(N__10787));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_3_LC_8_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_3_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_3_LC_8_7_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_3_LC_8_7_5  (
            .in0(N__7868),
            .in1(N__7432),
            .in2(_gnd_net_),
            .in3(N__5442),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_3_LC_8_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_3_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_3_LC_8_7_6 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_3_LC_8_7_6  (
            .in0(_gnd_net_),
            .in1(N__7268),
            .in2(N__4541),
            .in3(N__6375),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_410_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_7_7 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_7_7  (
            .in0(N__6146),
            .in1(N__7433),
            .in2(N__4538),
            .in3(N__5443),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_1_LC_8_8_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_8_8_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_8_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5872),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9807),
            .ce(),
            .sr(N__10780));
    defparam \U712_REG_SM.C3_SYNC_0_LC_8_8_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_8_8_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_8_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4525),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9807),
            .ce(),
            .sr(N__10780));
    defparam \U712_REG_SM.REG_TACK_LC_8_8_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_8_8_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_8_8_2  (
            .in0(N__4687),
            .in1(N__4676),
            .in2(N__5699),
            .in3(N__5353),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9807),
            .ce(),
            .sr(N__10780));
    defparam \U712_REG_SM.C1_SYNC_1_LC_8_8_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_8_8_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_8_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5920),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9807),
            .ce(),
            .sr(N__10780));
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_8_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_8_8_7 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_LC_8_8_7  (
            .in0(N__4648),
            .in1(N__5684),
            .in2(_gnd_net_),
            .in3(N__4670),
            .lcout(LATCH_CLK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9807),
            .ce(),
            .sr(N__10780));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_9_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_9_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__4902),
            .in2(_gnd_net_),
            .in3(N__4636),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_8_10_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_8_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4637),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9813),
            .ce(),
            .sr(N__10770));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_8_10_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_8_10_2 .LUT_INIT=16'b1110111000001010;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_8_10_2  (
            .in0(N__5290),
            .in1(N__8481),
            .in2(N__5330),
            .in3(N__4919),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9813),
            .ce(),
            .sr(N__10770));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_8_10_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_8_10_3 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_8_10_3  (
            .in0(N__4917),
            .in1(_gnd_net_),
            .in2(N__8483),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9813),
            .ce(),
            .sr(N__10770));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_8_10_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_8_10_4 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_8_10_4 .LUT_INIT=16'b0000000011111000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_8_10_4  (
            .in0(N__4625),
            .in1(N__5326),
            .in2(N__5309),
            .in3(N__4916),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9813),
            .ce(),
            .sr(N__10770));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_8_10_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_8_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_8_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_8_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4904),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9813),
            .ce(),
            .sr(N__10770));
    defparam DBR_SYNC_1_LC_8_10_6.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_8_10_6.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_8_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_8_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4931),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9813),
            .ce(),
            .sr(N__10770));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_10_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_10_7 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_10_7 .LUT_INIT=16'b1111111111000100;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_8_10_7  (
            .in0(N__4918),
            .in1(N__4876),
            .in2(N__8482),
            .in3(N__4903),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9813),
            .ce(),
            .sr(N__10770));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_11_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_11_3 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_11_3 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_11_3  (
            .in0(N__5325),
            .in1(N__8295),
            .in2(_gnd_net_),
            .in3(N__5291),
            .lcout(TACK_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9816),
            .ce(N__5267),
            .sr(N__10767));
    defparam CONSTANT_ONE_LUT4_LC_9_3_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_9_3_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_9_3_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_9_3_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_5_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_5_2  (
            .in0(N__4850),
            .in1(N__4832),
            .in2(_gnd_net_),
            .in3(N__9464),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_9_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_9_5_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_9_5_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_LC_9_5_4  (
            .in0(N__4814),
            .in1(N__5572),
            .in2(N__9682),
            .in3(N__4802),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9792),
            .ce(),
            .sr(N__10795));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_5_5 .LUT_INIT=16'b0011011100000101;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_5_5  (
            .in0(N__4796),
            .in1(N__9637),
            .in2(N__4766),
            .in3(N__5619),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9792),
            .ce(),
            .sr(N__10795));
    defparam \U712_CHIP_RAM.DBDIR_LC_9_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_9_5_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_9_5_7 .LUT_INIT=16'b0011101010101010;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_9_5_7  (
            .in0(N__4699),
            .in1(N__4748),
            .in2(N__7566),
            .in3(N__5002),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9792),
            .ce(),
            .sr(N__10795));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_6_0 .LUT_INIT=16'b1111101111110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_6_0  (
            .in0(N__5091),
            .in1(N__8392),
            .in2(N__5483),
            .in3(N__5020),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_6_1 .LUT_INIT=16'b0000111101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_6_1  (
            .in0(N__5041),
            .in1(N__7125),
            .in2(N__5024),
            .in3(N__6842),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9795),
            .ce(N__6796),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI49DCG_LC_9_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI49DCG_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI49DCG_LC_9_6_3 .LUT_INIT=16'b1111110111011101;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI49DCG_LC_9_6_3  (
            .in0(N__8390),
            .in1(N__5534),
            .in2(N__5021),
            .in3(N__5090),
            .lcout(\U712_CHIP_RAM.N_62 ),
            .ltout(\U712_CHIP_RAM.N_62_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_6_4 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_6_4  (
            .in0(N__4979),
            .in1(N__6671),
            .in2(N__5006),
            .in3(N__8391),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9795),
            .ce(N__6796),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIGGM16_LC_9_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIGGM16_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIGGM16_LC_9_6_5 .LUT_INIT=16'b1101111101011111;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIGGM16_LC_9_6_5  (
            .in0(N__7475),
            .in1(N__5672),
            .in2(N__5003),
            .in3(N__5618),
            .lcout(\U712_CHIP_RAM.N_434_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_3_LC_9_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_3_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_3_LC_9_6_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_3_LC_9_6_6  (
            .in0(N__7395),
            .in1(N__6357),
            .in2(N__7867),
            .in3(N__5454),
            .lcout(\U712_CHIP_RAM.N_452 ),
            .ltout(\U712_CHIP_RAM.N_452_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIQ6QH5_LC_9_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIQ6QH5_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIQ6QH5_LC_9_6_7 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIQ6QH5_LC_9_6_7  (
            .in0(_gnd_net_),
            .in1(N__7545),
            .in2(N__4982),
            .in3(N__5159),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_7_0 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_7_0  (
            .in0(N__7098),
            .in1(N__5384),
            .in2(N__7443),
            .in3(N__5365),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_7_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_7_1 .LUT_INIT=16'b1010001110101111;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_9_7_1  (
            .in0(N__4942),
            .in1(N__9681),
            .in2(N__4961),
            .in3(N__7973),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9800),
            .ce(),
            .sr(N__10781));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4GV43_2_LC_9_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4GV43_2_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4GV43_2_LC_9_7_2 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4GV43_2_LC_9_7_2  (
            .in0(N__7972),
            .in1(N__7871),
            .in2(_gnd_net_),
            .in3(N__5445),
            .lcout(\U712_CHIP_RAM.N_11_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_7_3 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_7_3  (
            .in0(N__5585),
            .in1(N__8388),
            .in2(N__5102),
            .in3(N__5111),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_9_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_9_7_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(N__7202),
            .in2(_gnd_net_),
            .in3(N__6066),
            .lcout(\U712_CHIP_RAM.N_288 ),
            .ltout(\U712_CHIP_RAM.N_288_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_2_LC_9_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_2_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_2_LC_9_7_5 .LUT_INIT=16'b0000100000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_2_LC_9_7_5  (
            .in0(N__5801),
            .in1(N__7971),
            .in2(N__5117),
            .in3(N__7097),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_372_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIADE59_LC_9_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIADE59_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIADE59_LC_9_7_6 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIADE59_LC_9_7_6  (
            .in0(N__8389),
            .in1(N__5498),
            .in2(N__5114),
            .in3(N__6067),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNILV2DI_LC_9_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNILV2DI_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNILV2DI_LC_9_7_7 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNILV2DI_LC_9_7_7  (
            .in0(N__5584),
            .in1(N__8387),
            .in2(N__5105),
            .in3(N__5094),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_7_1_LC_9_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_7_1_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_7_1_LC_9_8_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_7_1_LC_9_8_0  (
            .in0(N__8375),
            .in1(N__7217),
            .in2(_gnd_net_),
            .in3(N__7146),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_4_1_LC_9_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_4_1_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_4_1_LC_9_8_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_4_1_LC_9_8_1  (
            .in0(N__7436),
            .in1(N__6073),
            .in2(N__5060),
            .in3(N__7741),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_366_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_8_2 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_8_2  (
            .in0(N__8374),
            .in1(N__5204),
            .in2(N__5057),
            .in3(N__6088),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_9_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_9_8_3 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_9_8_3  (
            .in0(N__7437),
            .in1(N__6383),
            .in2(N__5054),
            .in3(N__5447),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_8_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__5213),
            .in2(N__5207),
            .in3(N__9420),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9805),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_5_1_LC_9_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_5_1_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_5_1_LC_9_8_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_5_1_LC_9_8_5  (
            .in0(N__7435),
            .in1(N__7870),
            .in2(_gnd_net_),
            .in3(N__6364),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_8_6  (
            .in0(N__5198),
            .in1(N__5180),
            .in2(_gnd_net_),
            .in3(N__9418),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_9_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_9_8_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_9_8_7  (
            .in0(N__9419),
            .in1(N__9644),
            .in2(N__5162),
            .in3(N__8513),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIEH9V_LC_9_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIEH9V_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIEH9V_LC_9_9_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIEH9V_LC_9_9_1  (
            .in0(N__5647),
            .in1(N__5620),
            .in2(_gnd_net_),
            .in3(N__6880),
            .lcout(\U712_CHIP_RAM.N_448 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_9_2 .LUT_INIT=16'b1100110000100010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_9_2  (
            .in0(N__7286),
            .in1(N__7438),
            .in2(_gnd_net_),
            .in3(N__7126),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_345_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_9_3 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_9_3  (
            .in0(N__9645),
            .in1(N__7745),
            .in2(N__5150),
            .in3(N__6087),
            .lcout(\U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_9_6  (
            .in0(N__5147),
            .in1(N__5132),
            .in2(_gnd_net_),
            .in3(N__9417),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_9_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_9_10_1 .LUT_INIT=16'b1111110011011100;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_9_10_1  (
            .in0(N__7151),
            .in1(N__6317),
            .in2(N__7445),
            .in3(N__7294),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_9_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_9_10_2 .LUT_INIT=16'b1100110011000101;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_9_10_2  (
            .in0(N__5378),
            .in1(N__5339),
            .in2(N__5372),
            .in3(N__5369),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9809),
            .ce(),
            .sr(N__10768));
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_9_10_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_9_10_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN6_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__5354),
            .in2(_gnd_net_),
            .in3(N__5338),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(\U712_CYCLE_TERM.TACK_EN6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_10_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_10_5 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_10_5  (
            .in0(N__8373),
            .in1(N__5305),
            .in2(N__5294),
            .in3(N__5289),
            .lcout(\U712_CYCLE_TERM.N_316_i_0_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_9_11_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_9_11_1 .LUT_INIT=16'b0000001010101010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_9_11_1  (
            .in0(N__9704),
            .in1(N__10328),
            .in2(N__10246),
            .in3(N__5261),
            .lcout(\U712_BYTE_ENABLE.un1_CUUBEn_i_0_aZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_11_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_11_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_11_2  (
            .in0(N__10822),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5273),
            .lcout(\U712_CYCLE_TERM.N_316_i_0_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_9_12_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_9_12_2 .LUT_INIT=16'b0000100010101010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_9_12_2  (
            .in0(N__9705),
            .in1(N__10322),
            .in2(N__10244),
            .in3(N__5257),
            .lcout(\U712_BYTE_ENABLE.un1_CLMBEn_i_0_aZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_x2_LC_9_13_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_x2_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_x2_LC_9_13_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_x2_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(N__10055),
            .in2(_gnd_net_),
            .in3(N__10139),
            .lcout(\U712_BYTE_ENABLE.N_282_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_4_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_4_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_4_3  (
            .in0(N__5246),
            .in1(N__5231),
            .in2(_gnd_net_),
            .in3(N__9525),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_0_2_LC_10_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_0_2_LC_10_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_0_2_LC_10_5_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_0_2_LC_10_5_2  (
            .in0(_gnd_net_),
            .in1(N__7832),
            .in2(_gnd_net_),
            .in3(N__7923),
            .lcout(\U712_CHIP_RAM.N_371_1 ),
            .ltout(\U712_CHIP_RAM.N_371_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_10_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_10_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_10_5_3 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_10_5_3  (
            .in0(N__7378),
            .in1(N__7193),
            .in2(N__5501),
            .in3(N__7072),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_5_4 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_5_4  (
            .in0(N__5468),
            .in1(N__7380),
            .in2(_gnd_net_),
            .in3(N__5525),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI27TJ3_LC_10_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI27TJ3_LC_10_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI27TJ3_LC_10_5_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI27TJ3_LC_10_5_6  (
            .in0(N__7194),
            .in1(N__5474),
            .in2(N__6089),
            .in3(N__7379),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_5_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5462),
            .in3(N__7195),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9789),
            .ce(),
            .sr(N__10788));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_10_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_10_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_10_6_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_10_6_1  (
            .in0(N__7813),
            .in1(N__7416),
            .in2(N__6376),
            .in3(N__5448),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9793),
            .ce(N__5396),
            .sr(N__10782));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI68LV_LC_10_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI68LV_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI68LV_LC_10_6_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI68LV_LC_10_6_2  (
            .in0(N__7588),
            .in1(N__7069),
            .in2(_gnd_net_),
            .in3(N__7808),
            .lcout(\U712_CHIP_RAM.N_436 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_6_3 .LUT_INIT=16'b1110111111111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_6_3  (
            .in0(N__7812),
            .in1(N__7415),
            .in2(N__7968),
            .in3(N__7121),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_i_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_6_4 .LUT_INIT=16'b1110111010101100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_6_4  (
            .in0(N__7414),
            .in1(N__7070),
            .in2(N__7967),
            .in3(N__7811),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_129_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_6_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_6_5  (
            .in0(N__7810),
            .in1(N__7285),
            .in2(_gnd_net_),
            .in3(N__7945),
            .lcout(\U712_CHIP_RAM.N_329 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_2_LC_10_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_2_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_2_LC_10_6_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_2_LC_10_6_6  (
            .in0(N__7413),
            .in1(N__7809),
            .in2(N__7142),
            .in3(N__6074),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_414_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_10_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_10_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_10_6_7 .LUT_INIT=16'b1111101111110011;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_10_6_7  (
            .in0(N__7546),
            .in1(N__7589),
            .in2(N__5687),
            .in3(N__5563),
            .lcout(\U712_CHIP_RAM.N_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIIPOI5_LC_10_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIIPOI5_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIIPOI5_LC_10_7_0 .LUT_INIT=16'b0100110000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIIPOI5_LC_10_7_0  (
            .in0(N__5670),
            .in1(N__7468),
            .in2(N__5624),
            .in3(N__5520),
            .lcout(\U712_CHIP_RAM.N_373 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_3_LC_10_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_3_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_3_LC_10_7_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_3_LC_10_7_1  (
            .in0(N__6356),
            .in1(N__7386),
            .in2(N__7848),
            .in3(N__6068),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER15 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4F6EB_LC_10_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4F6EB_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4F6EB_LC_10_7_2 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4F6EB_LC_10_7_2  (
            .in0(N__6069),
            .in1(N__5507),
            .in2(N__5537),
            .in3(N__5521),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_7_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_7_3  (
            .in0(N__6619),
            .in1(N__6634),
            .in2(N__6812),
            .in3(N__6649),
            .lcout(\U712_CHIP_RAM.N_286 ),
            .ltout(\U712_CHIP_RAM.N_286_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI16TJ3_LC_10_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI16TJ3_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI16TJ3_LC_10_7_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI16TJ3_LC_10_7_4  (
            .in0(N__7209),
            .in1(N__7819),
            .in2(N__5528),
            .in3(N__6355),
            .lcout(\U712_CHIP_RAM.N_486 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_0_LC_10_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_0_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_0_LC_10_7_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_0_LC_10_7_5  (
            .in0(N__6354),
            .in1(N__7385),
            .in2(N__7847),
            .in3(N__7210),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_2_LC_10_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_2_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_2_LC_10_7_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_2_LC_10_7_6  (
            .in0(_gnd_net_),
            .in1(N__7922),
            .in2(_gnd_net_),
            .in3(N__7071),
            .lcout(\U712_CHIP_RAM.N_287 ),
            .ltout(\U712_CHIP_RAM.N_287_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIF74S2_LC_10_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIF74S2_LC_10_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIF74S2_LC_10_7_7 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIF74S2_LC_10_7_7  (
            .in0(N__7815),
            .in1(N__7510),
            .in2(N__6161),
            .in3(N__6158),
            .lcout(\U712_CHIP_RAM.N_283 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_8_0 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_8_0  (
            .in0(N__8362),
            .in1(N__7007),
            .in2(N__6122),
            .in3(N__6082),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9801),
            .ce(N__6017),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_8_1 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_8_1  (
            .in0(N__6081),
            .in1(N__8363),
            .in2(_gnd_net_),
            .in3(N__6110),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9801),
            .ce(N__6017),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_8_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_8_2  (
            .in0(N__8364),
            .in1(N__6305),
            .in2(N__6101),
            .in3(N__6083),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9801),
            .ce(N__6017),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNIAS4F1_0_1_LC_10_8_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNIAS4F1_0_1_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNIAS4F1_0_1_LC_10_8_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNIAS4F1_0_1_LC_10_8_4  (
            .in0(N__5993),
            .in1(N__5949),
            .in2(N__5924),
            .in3(N__5873),
            .lcout(\U712_REG_SM.C1_SYNC_RNIAS4F1_0Z0Z_1 ),
            .ltout(\U712_REG_SM.C1_SYNC_RNIAS4F1_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIOC3L1_4_LC_10_8_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIOC3L1_4_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIOC3L1_4_LC_10_8_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIOC3L1_4_LC_10_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5825),
            .in3(N__5791),
            .lcout(\U712_REG_SM.ASn_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIKPND1_3_LC_10_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIKPND1_3_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIKPND1_3_LC_10_8_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIKPND1_3_LC_10_8_6  (
            .in0(N__7849),
            .in1(N__7426),
            .in2(_gnd_net_),
            .in3(N__8372),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_8_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_8_7 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_10_8_7  (
            .in0(N__6563),
            .in1(N__5792),
            .in2(N__5759),
            .in3(N__5712),
            .lcout(\U712_REG_SM.N_104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_6_1_LC_10_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_6_1_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_6_1_LC_10_9_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_6_1_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(N__7521),
            .in2(_gnd_net_),
            .in3(N__6869),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_RNO_6Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_10_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_10_9_4 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_10_9_4  (
            .in0(N__7965),
            .in1(N__8361),
            .in2(N__6386),
            .in3(N__7144),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_10_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_10_9_5 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_10_9_5  (
            .in0(N__7287),
            .in1(N__7850),
            .in2(_gnd_net_),
            .in3(N__6374),
            .lcout(\U712_CHIP_RAM.N_388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_9_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_9_6  (
            .in0(N__7966),
            .in1(N__7218),
            .in2(_gnd_net_),
            .in3(N__7145),
            .lcout(\U712_CHIP_RAM.N_370 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_38_i_LC_10_10_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_38_i_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_38_i_LC_10_10_0 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \U712_BYTE_ENABLE.N_38_i_LC_10_10_0  (
            .in0(N__8191),
            .in1(N__6299),
            .in2(N__6228),
            .in3(N__7609),
            .lcout(N_38_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_1_LC_10_10_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_1_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_1_LC_10_10_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_1_LC_10_10_1  (
            .in0(N__7612),
            .in1(N__8252),
            .in2(_gnd_net_),
            .in3(N__6224),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_426_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_47_i_LC_10_10_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_47_i_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_47_i_LC_10_10_2 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \U712_BYTE_ENABLE.N_47_i_LC_10_10_2  (
            .in0(N__6605),
            .in1(N__6572),
            .in2(N__6269),
            .in3(N__10327),
            .lcout(N_47_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_10_10_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_10_10_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_10_10_3  (
            .in0(N__7611),
            .in1(N__8251),
            .in2(_gnd_net_),
            .in3(N__6223),
            .lcout(\U712_BYTE_ENABLE.N_431 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_46_i_LC_10_10_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_46_i_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_46_i_LC_10_10_4 .LUT_INIT=16'b0011001000110011;
    LogicCell40 \U712_BYTE_ENABLE.N_46_i_LC_10_10_4  (
            .in0(N__8192),
            .in1(N__6242),
            .in2(N__6229),
            .in3(N__7610),
            .lcout(N_46_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_LC_10_10_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_LC_10_10_5 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_LC_10_10_5  (
            .in0(N__10061),
            .in1(N__10157),
            .in2(_gnd_net_),
            .in3(N__9706),
            .lcout(\U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2Z0Z_0 ),
            .ltout(\U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_45_i_LC_10_10_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_45_i_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_45_i_LC_10_10_6 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \U712_BYTE_ENABLE.N_45_i_LC_10_10_6  (
            .in0(N__6596),
            .in1(N__10326),
            .in2(N__6590),
            .in3(N__6571),
            .lcout(N_45_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_1_LC_10_11_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_1_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_1_LC_10_11_0 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_1_LC_10_11_0  (
            .in0(N__9707),
            .in1(N__10245),
            .in2(_gnd_net_),
            .in3(N__10156),
            .lcout(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DRDDIR_0_m2_i_m2_LC_10_18_0 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_0_m2_i_m2_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_0_m2_i_m2_LC_10_18_0 .LUT_INIT=16'b0010000001111111;
    LogicCell40 \U712_BUFFERS.DRDDIR_0_m2_i_m2_LC_10_18_0  (
            .in0(N__8172),
            .in1(N__6555),
            .in2(N__8241),
            .in3(N__7304),
            .lcout(N_344),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DMA_LATCH_EN_0_a2_0_a2_LC_10_18_2 .C_ON=1'b0;
    defparam \U712_BUFFERS.DMA_LATCH_EN_0_a2_0_a2_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DMA_LATCH_EN_0_a2_0_a2_LC_10_18_2 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \U712_BUFFERS.DMA_LATCH_EN_0_a2_0_a2_LC_10_18_2  (
            .in0(N__8171),
            .in1(N__8232),
            .in2(_gnd_net_),
            .in3(N__7303),
            .lcout(DMA_LATCH_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_5 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_5  (
            .in0(N__9703),
            .in1(N__6464),
            .in2(N__9527),
            .in3(N__9335),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_5_3 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_5_3  (
            .in0(N__6458),
            .in1(N__9522),
            .in2(N__9695),
            .in3(N__8975),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_11_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_11_5_4 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_11_5_4  (
            .in0(N__8770),
            .in1(N__8719),
            .in2(N__6449),
            .in3(N__9002),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9786),
            .ce(N__9127),
            .sr(N__10783));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_11_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_11_5_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_11_5_5  (
            .in0(N__6425),
            .in1(N__6404),
            .in2(_gnd_net_),
            .in3(N__9521),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_5_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_5_6  (
            .in0(N__8501),
            .in1(N__9523),
            .in2(N__6698),
            .in3(N__9661),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_11_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_11_5_7 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_11_5_7  (
            .in0(N__8718),
            .in1(N__7715),
            .in2(N__6695),
            .in3(N__8771),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9786),
            .ce(N__9127),
            .sr(N__10783));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_cry_c_0_LC_11_6_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_cry_c_0_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_cry_c_0_LC_11_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_cry_c_0_LC_11_6_0  (
            .in0(_gnd_net_),
            .in1(N__7114),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_11_6_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_11_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(N__7439),
            .in2(_gnd_net_),
            .in3(N__6659),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_6_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_6_2  (
            .in0(N__6846),
            .in1(N__7949),
            .in2(_gnd_net_),
            .in3(N__6656),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(N__9790),
            .ce(N__6797),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_6_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_6_3  (
            .in0(N__6843),
            .in1(N__7846),
            .in2(_gnd_net_),
            .in3(N__6653),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__9790),
            .ce(N__6797),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_6_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_6_4  (
            .in0(N__6847),
            .in1(N__6650),
            .in2(_gnd_net_),
            .in3(N__6638),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__9790),
            .ce(N__6797),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_11_6_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_11_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_11_6_5  (
            .in0(N__6844),
            .in1(N__6635),
            .in2(_gnd_net_),
            .in3(N__6623),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__9790),
            .ce(N__6797),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_6_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_6_6  (
            .in0(N__6848),
            .in1(N__6620),
            .in2(_gnd_net_),
            .in3(N__6608),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__9790),
            .ce(N__6797),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_6_7  (
            .in0(N__6845),
            .in1(N__6811),
            .in2(_gnd_net_),
            .in3(N__6815),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9790),
            .ce(N__6797),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_7_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_7_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__6962),
            .in2(_gnd_net_),
            .in3(N__6779),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__6733),
            .ce(),
            .sr(N__7457));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_7_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_7_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__7001),
            .in2(_gnd_net_),
            .in3(N__6776),
            .lcout(\U712_CHIP_RAM.REFRESH5lto1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__6733),
            .ce(),
            .sr(N__7457));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_7_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_7_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__6976),
            .in2(_gnd_net_),
            .in3(N__6773),
            .lcout(\U712_CHIP_RAM.REFRESH5lto2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__6733),
            .ce(),
            .sr(N__7457));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_7_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_7_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__6925),
            .in2(_gnd_net_),
            .in3(N__6770),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__6733),
            .ce(),
            .sr(N__7457));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_7_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_7_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__6989),
            .in2(_gnd_net_),
            .in3(N__6767),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__6733),
            .ce(),
            .sr(N__7457));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_7_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_7_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__6938),
            .in2(_gnd_net_),
            .in3(N__6764),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__6733),
            .ce(),
            .sr(N__7457));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_7_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_7_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(N__6950),
            .in2(_gnd_net_),
            .in3(N__6761),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__6733),
            .ce(),
            .sr(N__7457));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_7_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_7_7  (
            .in0(_gnd_net_),
            .in1(N__6901),
            .in2(_gnd_net_),
            .in3(N__6758),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6733),
            .ce(),
            .sr(N__7457));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_8_0 .LUT_INIT=16'b1011111110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_8_0  (
            .in0(N__7706),
            .in1(N__8359),
            .in2(N__7616),
            .in3(N__7512),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9796),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIHSHE1_LC_11_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIHSHE1_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIHSHE1_LC_11_8_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIHSHE1_LC_11_8_2  (
            .in0(N__6870),
            .in1(N__8360),
            .in2(_gnd_net_),
            .in3(N__7511),
            .lcout(\U712_CHIP_RAM.N_201_i_i_a2_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_8_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_8_3  (
            .in0(N__9860),
            .in1(N__9933),
            .in2(N__8861),
            .in3(N__9442),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_11_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_11_8_4 .LUT_INIT=16'b1011101110111011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_11_8_4  (
            .in0(N__7444),
            .in1(N__7284),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_306_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_11_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_11_8_5 .LUT_INIT=16'b1010000011100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_11_8_5  (
            .in0(N__7851),
            .in1(N__7220),
            .in2(N__7154),
            .in3(N__7143),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_8_6 .LUT_INIT=16'b0011011100111111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_8_6  (
            .in0(N__7000),
            .in1(N__6988),
            .in2(N__6977),
            .in3(N__6961),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(N__6949),
            .in2(_gnd_net_),
            .in3(N__6937),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_11_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_11_9_3 .LUT_INIT=16'b1111001111111011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_11_9_3  (
            .in0(N__6926),
            .in1(N__6911),
            .in2(N__6905),
            .in3(N__6887),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9802),
            .ce(),
            .sr(N__10761));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_11_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_11_10_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__8190),
            .in2(_gnd_net_),
            .in3(N__8250),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9806),
            .ce(),
            .sr(N__10758));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_10_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(N__7688),
            .in2(_gnd_net_),
            .in3(N__7696),
            .lcout(\U712_CHIP_RAM.un3_DMA_CYCLE_START ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_11_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_11_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_11_10_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_11_10_5  (
            .in0(N__7697),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9806),
            .ce(),
            .sr(N__10758));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_4_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_4_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_12_4_7  (
            .in0(N__8717),
            .in1(N__9065),
            .in2(N__8781),
            .in3(N__7682),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9783),
            .ce(N__9128),
            .sr(N__10778));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_5_0 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_5_0  (
            .in0(N__7658),
            .in1(N__9498),
            .in2(N__9710),
            .in3(N__9353),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_5_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_5_2  (
            .in0(N__10823),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7979),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_12_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_12_5_3 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_12_5_3  (
            .in0(N__9494),
            .in1(N__9893),
            .in2(_gnd_net_),
            .in3(N__9963),
            .lcout(\U712_CHIP_RAM.CMA_5_0_8 ),
            .ltout(\U712_CHIP_RAM.CMA_5_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_5_4 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_5_4  (
            .in0(N__7639),
            .in1(N__9657),
            .in2(N__7643),
            .in3(N__8524),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_5_6 .LUT_INIT=16'b1011111110001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_5_6  (
            .in0(N__7640),
            .in1(N__9656),
            .in2(N__8602),
            .in3(N__8525),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNI8NM9_LC_12_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNI8NM9_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNI8NM9_LC_12_5_7 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_RNI8NM9_LC_12_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9524),
            .in3(N__9699),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_6_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(N__9889),
            .in2(_gnd_net_),
            .in3(N__9959),
            .lcout(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_6_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_6_1  (
            .in0(N__8003),
            .in1(N__9689),
            .in2(_gnd_net_),
            .in3(N__8492),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_463_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_6_2 .LUT_INIT=16'b0101010111110000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_6_2  (
            .in0(N__9493),
            .in1(_gnd_net_),
            .in2(N__7982),
            .in3(N__8758),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_6_3 .LUT_INIT=16'b0101111101001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_6_3  (
            .in0(N__8757),
            .in1(N__10520),
            .in2(N__9531),
            .in3(N__9690),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_6_4 .LUT_INIT=16'b0011001100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_6_4  (
            .in0(N__10519),
            .in1(N__9512),
            .in2(N__9708),
            .in3(N__8759),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_6_5 .LUT_INIT=16'b0000001100110001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_6_5  (
            .in0(N__9958),
            .in1(N__8871),
            .in2(N__9895),
            .in3(N__9492),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_12_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_12_6_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_12_6_7  (
            .in0(N__7921),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7814),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_12_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_12_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_12_7_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_12_7_0  (
            .in0(N__9323),
            .in1(N__11062),
            .in2(_gnd_net_),
            .in3(N__9040),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10888),
            .ce(N__10857),
            .sr(N__10766));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_7_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_7_5  (
            .in0(N__11061),
            .in1(N__9322),
            .in2(_gnd_net_),
            .in3(N__9275),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10888),
            .ce(N__10857),
            .sr(N__10766));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_12_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_12_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_12_8_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_12_8_0  (
            .in0(N__10466),
            .in1(N__9274),
            .in2(_gnd_net_),
            .in3(N__11059),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .ce(N__10855),
            .sr(N__10760));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_12_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_12_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_12_8_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_12_8_3  (
            .in0(N__11060),
            .in1(N__9224),
            .in2(_gnd_net_),
            .in3(N__9039),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .ce(N__10855),
            .sr(N__10760));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_12_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_12_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_12_9_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_12_9_4  (
            .in0(N__9026),
            .in1(N__11053),
            .in2(_gnd_net_),
            .in3(N__9321),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__10853),
            .sr(N__10757));
    defparam pll_RNI8MQ3_LC_12_10_6.C_ON=1'b0;
    defparam pll_RNI8MQ3_LC_12_10_6.SEQ_MODE=4'b0000;
    defparam pll_RNI8MQ3_LC_12_10_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 pll_RNI8MQ3_LC_12_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8474),
            .lcout(CLK40_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_16_1.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_16_1.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_16_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_16_1 (
            .in0(N__8393),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_12_17_0 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_12_17_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_0_a2_LC_12_17_0  (
            .in0(N__8215),
            .in1(N__8189),
            .in2(_gnd_net_),
            .in3(N__8124),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CRCSn_LC_13_2_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_13_2_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_13_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_13_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8876),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9782),
            .ce(),
            .sr(N__10803));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_4_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_4_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_13_4_7  (
            .in0(N__8720),
            .in1(N__10403),
            .in2(N__8783),
            .in3(N__8039),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9784),
            .ce(N__9130),
            .sr(N__10789));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_5_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_5_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_13_5_0  (
            .in0(N__8715),
            .in1(N__8930),
            .in2(N__8782),
            .in3(N__8900),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9787),
            .ce(N__9129),
            .sr(N__10784));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_13_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_13_5_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_13_5_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_13_5_1  (
            .in0(N__9968),
            .in1(N__9894),
            .in2(N__9526),
            .in3(N__8875),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9787),
            .ce(N__9129),
            .sr(N__10784));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_5_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_13_5_2  (
            .in0(N__8822),
            .in1(N__8816),
            .in2(_gnd_net_),
            .in3(N__8810),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9787),
            .ce(N__9129),
            .sr(N__10784));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_13_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_13_5_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_13_5_3 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_13_5_3  (
            .in0(N__8766),
            .in1(N__8716),
            .in2(N__9053),
            .in3(N__9359),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9787),
            .ce(N__9129),
            .sr(N__10784));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_5_6 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_13_5_6  (
            .in0(N__9673),
            .in1(N__8669),
            .in2(N__8603),
            .in3(N__10901),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9787),
            .ce(N__9129),
            .sr(N__10784));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_5_7 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_13_5_7  (
            .in0(N__9179),
            .in1(N__9674),
            .in2(N__8627),
            .in3(N__8601),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9787),
            .ce(N__9129),
            .sr(N__10784));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_13_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_13_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_13_6_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_13_6_2  (
            .in0(N__8561),
            .in1(N__8540),
            .in2(_gnd_net_),
            .in3(N__9519),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_6_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_6_3  (
            .in0(N__9520),
            .in1(N__9694),
            .in2(N__8528),
            .in3(N__9341),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_13_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_13_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_13_6_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_13_6_4  (
            .in0(_gnd_net_),
            .in1(N__9170),
            .in2(N__9164),
            .in3(N__9161),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9791),
            .ce(N__9137),
            .sr(N__10776));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_13_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_13_7_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_13_7_4  (
            .in0(N__9101),
            .in1(N__9083),
            .in2(_gnd_net_),
            .in3(N__9502),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_0  (
            .in0(N__10613),
            .in1(N__11054),
            .in2(_gnd_net_),
            .in3(N__10505),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10887),
            .ce(N__10858),
            .sr(N__10769));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_8_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_8_4  (
            .in0(N__9267),
            .in1(N__11055),
            .in2(_gnd_net_),
            .in3(N__10465),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10887),
            .ce(N__10858),
            .sr(N__10769));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_8_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_8_7  (
            .in0(N__9223),
            .in1(_gnd_net_),
            .in2(N__11070),
            .in3(N__9041),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10887),
            .ce(N__10858),
            .sr(N__10769));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_9_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_13_9_4  (
            .in0(N__8960),
            .in1(N__11049),
            .in2(_gnd_net_),
            .in3(N__10568),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__10856),
            .sr(N__10762));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_7  (
            .in0(N__11145),
            .in1(_gnd_net_),
            .in2(N__11069),
            .in3(N__9207),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__10856),
            .sr(N__10762));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_10_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_10_3  (
            .in0(N__11016),
            .in1(N__10575),
            .in2(_gnd_net_),
            .in3(N__8956),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10884),
            .ce(N__10854),
            .sr(N__10759));
    defparam \U712_CHIP_RAM.CASn_LC_14_3_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_14_3_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_14_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_14_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9532),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9785),
            .ce(),
            .sr(N__10804));
    defparam \U712_CHIP_RAM.WEn_LC_14_3_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_14_3_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_14_3_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_14_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9967),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9785),
            .ce(),
            .sr(N__10804));
    defparam \U712_CHIP_RAM.RASn_LC_14_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_14_4_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_14_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_14_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9896),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9788),
            .ce(),
            .sr(N__10796));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_6_0 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_6_0  (
            .in0(N__9709),
            .in1(N__9539),
            .in2(N__9533),
            .in3(N__9230),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_7_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_7_1  (
            .in0(N__11000),
            .in1(N__10608),
            .in2(_gnd_net_),
            .in3(N__10577),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__10860),
            .sr(N__10777));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_7_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_7_2  (
            .in0(N__10609),
            .in1(N__11001),
            .in2(_gnd_net_),
            .in3(N__10500),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__10860),
            .sr(N__10777));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_7_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_7_3  (
            .in0(N__10501),
            .in1(N__11002),
            .in2(_gnd_net_),
            .in3(N__10464),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__10860),
            .sr(N__10777));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_7_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_7_5  (
            .in0(N__9306),
            .in1(N__11003),
            .in2(_gnd_net_),
            .in3(N__9258),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__10860),
            .sr(N__10777));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_8_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_8_0  (
            .in0(N__9216),
            .in1(N__11012),
            .in2(_gnd_net_),
            .in3(N__11152),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10885),
            .ce(N__10859),
            .sr(N__10771));
    defparam \U712_BYTE_ENABLE.N_357_i_LC_14_19_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_357_i_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_357_i_LC_14_19_3 .LUT_INIT=16'b0000111011100000;
    LogicCell40 \U712_BYTE_ENABLE.N_357_i_LC_14_19_3  (
            .in0(N__10276),
            .in1(N__10236),
            .in2(N__10155),
            .in3(N__10035),
            .lcout(N_357_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_0_LC_14_20_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_0_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_0_LC_14_20_4 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \U712_BYTE_ENABLE.un1_UDSn_i_0_0_LC_14_20_4  (
            .in0(N__10241),
            .in1(N__10376),
            .in2(_gnd_net_),
            .in3(N__10122),
            .lcout(N_42),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UMBE_i_o2_i_LC_14_20_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UMBE_i_o2_i_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UMBE_i_o2_i_LC_14_20_6 .LUT_INIT=16'b0000110111000000;
    LogicCell40 \U712_BYTE_ENABLE.UMBE_i_o2_i_LC_14_20_6  (
            .in0(N__10240),
            .in1(N__10306),
            .in2(N__10048),
            .in3(N__10121),
            .lcout(N_231),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_7_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_7_1  (
            .in0(N__10996),
            .in1(N__10607),
            .in2(_gnd_net_),
            .in3(N__10576),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10886),
            .ce(N__10861),
            .sr(N__10785));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_7_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_7_3  (
            .in0(N__10499),
            .in1(_gnd_net_),
            .in2(N__11032),
            .in3(N__10454),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10886),
            .ce(N__10861),
            .sr(N__10785));
    defparam \U712_BYTE_ENABLE.N_358_i_LC_15_19_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_358_i_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_358_i_LC_15_19_6 .LUT_INIT=16'b0011000111000100;
    LogicCell40 \U712_BYTE_ENABLE.N_358_i_LC_15_19_6  (
            .in0(N__10291),
            .in1(N__10060),
            .in2(N__10247),
            .in3(N__10147),
            .lcout(N_358_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_15_20_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_15_20_1 .LUT_INIT=16'b0010001011111111;
    LogicCell40 \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_15_20_1  (
            .in0(N__10143),
            .in1(N__10243),
            .in2(_gnd_net_),
            .in3(N__10375),
            .lcout(N_40),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LLBE_0_0_LC_15_20_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LLBE_0_0_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LLBE_0_0_LC_15_20_7 .LUT_INIT=16'b0000010101110000;
    LogicCell40 \U712_BYTE_ENABLE.LLBE_0_0_LC_15_20_7  (
            .in0(N__10307),
            .in1(N__10242),
            .in2(N__10154),
            .in3(N__10059),
            .lcout(LLBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_22_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_22_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_22_8_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_22_8_1  (
            .in0(N__11127),
            .in1(N__11084),
            .in2(_gnd_net_),
            .in3(N__11048),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10883),
            .ce(N__10862),
            .sr(N__10807));
endmodule // U712_TOP
